module systemcomplete (clk, reset, data_in, target, finished, nonce_out);

input clk;
input reset;
output finished;
input [95:0] data_in;
input [7:0] target;
output [31:0] nonce_out;

wire vdd = 1'b1;
wire gnd = 1'b0;

BUFX4 BUFX4_1 ( .A(clk), .Y(clk_hier0_bF_buf8) );
BUFX4 BUFX4_2 ( .A(clk), .Y(clk_hier0_bF_buf7) );
BUFX4 BUFX4_3 ( .A(clk), .Y(clk_hier0_bF_buf6) );
BUFX4 BUFX4_4 ( .A(clk), .Y(clk_hier0_bF_buf5) );
BUFX4 BUFX4_5 ( .A(clk), .Y(clk_hier0_bF_buf4) );
BUFX4 BUFX4_6 ( .A(clk), .Y(clk_hier0_bF_buf3) );
BUFX4 BUFX4_7 ( .A(clk), .Y(clk_hier0_bF_buf2) );
BUFX4 BUFX4_8 ( .A(clk), .Y(clk_hier0_bF_buf1) );
BUFX4 BUFX4_9 ( .A(clk), .Y(clk_hier0_bF_buf0) );
BUFX4 BUFX4_10 ( .A(_4283_), .Y(_4283__hier0_bF_buf5) );
BUFX4 BUFX4_11 ( .A(_4283_), .Y(_4283__hier0_bF_buf4) );
BUFX4 BUFX4_12 ( .A(_4283_), .Y(_4283__hier0_bF_buf3) );
BUFX4 BUFX4_13 ( .A(_4283_), .Y(_4283__hier0_bF_buf2) );
BUFX4 BUFX4_14 ( .A(_4283_), .Y(_4283__hier0_bF_buf1) );
BUFX4 BUFX4_15 ( .A(_4283_), .Y(_4283__hier0_bF_buf0) );
BUFX4 BUFX4_16 ( .A(_588_), .Y(_588__bF_buf4) );
BUFX4 BUFX4_17 ( .A(_588_), .Y(_588__bF_buf3) );
BUFX4 BUFX4_18 ( .A(_588_), .Y(_588__bF_buf2) );
BUFX4 BUFX4_19 ( .A(_588_), .Y(_588__bF_buf1) );
BUFX4 BUFX4_20 ( .A(_588_), .Y(_588__bF_buf0) );
BUFX4 BUFX4_21 ( .A(_4226_), .Y(_4226__bF_buf3) );
BUFX4 BUFX4_22 ( .A(_4226_), .Y(_4226__bF_buf2) );
BUFX4 BUFX4_23 ( .A(_4226_), .Y(_4226__bF_buf1) );
BUFX4 BUFX4_24 ( .A(_4226_), .Y(_4226__bF_buf0) );
BUFX4 BUFX4_25 ( .A(_1122_), .Y(_1122__bF_buf4) );
BUFX4 BUFX4_26 ( .A(_1122_), .Y(_1122__bF_buf3) );
BUFX4 BUFX4_27 ( .A(_1122_), .Y(_1122__bF_buf2) );
BUFX4 BUFX4_28 ( .A(_1122_), .Y(_1122__bF_buf1) );
BUFX4 BUFX4_29 ( .A(_1122_), .Y(_1122__bF_buf0) );
BUFX4 BUFX4_30 ( .A(_832_), .Y(_832__bF_buf4) );
BUFX4 BUFX4_31 ( .A(_832_), .Y(_832__bF_buf3) );
BUFX4 BUFX4_32 ( .A(_832_), .Y(_832__bF_buf2) );
BUFX4 BUFX4_33 ( .A(_832_), .Y(_832__bF_buf1) );
BUFX4 BUFX4_34 ( .A(_832_), .Y(_832__bF_buf0) );
BUFX4 BUFX4_35 ( .A(micro_hash_ucr_pipe50), .Y(micro_hash_ucr_pipe50_bF_buf3) );
BUFX4 BUFX4_36 ( .A(micro_hash_ucr_pipe50), .Y(micro_hash_ucr_pipe50_bF_buf2) );
BUFX4 BUFX4_37 ( .A(micro_hash_ucr_pipe50), .Y(micro_hash_ucr_pipe50_bF_buf1) );
BUFX4 BUFX4_38 ( .A(micro_hash_ucr_pipe50), .Y(micro_hash_ucr_pipe50_bF_buf0) );
BUFX4 BUFX4_39 ( .A(micro_hash_ucr_pipe52), .Y(micro_hash_ucr_pipe52_bF_buf3) );
BUFX4 BUFX4_40 ( .A(micro_hash_ucr_pipe52), .Y(micro_hash_ucr_pipe52_bF_buf2) );
BUFX4 BUFX4_41 ( .A(micro_hash_ucr_pipe52), .Y(micro_hash_ucr_pipe52_bF_buf1) );
BUFX4 BUFX4_42 ( .A(micro_hash_ucr_pipe52), .Y(micro_hash_ucr_pipe52_bF_buf0) );
BUFX4 BUFX4_43 ( .A(micro_hash_ucr_pipe53), .Y(micro_hash_ucr_pipe53_bF_buf3) );
BUFX4 BUFX4_44 ( .A(micro_hash_ucr_pipe53), .Y(micro_hash_ucr_pipe53_bF_buf2) );
BUFX4 BUFX4_45 ( .A(micro_hash_ucr_pipe53), .Y(micro_hash_ucr_pipe53_bF_buf1) );
BUFX4 BUFX4_46 ( .A(micro_hash_ucr_pipe53), .Y(micro_hash_ucr_pipe53_bF_buf0) );
BUFX4 BUFX4_47 ( .A(micro_hash_ucr_pipe54), .Y(micro_hash_ucr_pipe54_bF_buf4) );
BUFX4 BUFX4_48 ( .A(micro_hash_ucr_pipe54), .Y(micro_hash_ucr_pipe54_bF_buf3) );
BUFX4 BUFX4_49 ( .A(micro_hash_ucr_pipe54), .Y(micro_hash_ucr_pipe54_bF_buf2) );
BUFX4 BUFX4_50 ( .A(micro_hash_ucr_pipe54), .Y(micro_hash_ucr_pipe54_bF_buf1) );
BUFX4 BUFX4_51 ( .A(micro_hash_ucr_pipe54), .Y(micro_hash_ucr_pipe54_bF_buf0) );
BUFX4 BUFX4_52 ( .A(micro_hash_ucr_pipe56), .Y(micro_hash_ucr_pipe56_bF_buf3) );
BUFX4 BUFX4_53 ( .A(micro_hash_ucr_pipe56), .Y(micro_hash_ucr_pipe56_bF_buf2) );
BUFX4 BUFX4_54 ( .A(micro_hash_ucr_pipe56), .Y(micro_hash_ucr_pipe56_bF_buf1) );
BUFX4 BUFX4_55 ( .A(micro_hash_ucr_pipe56), .Y(micro_hash_ucr_pipe56_bF_buf0) );
BUFX4 BUFX4_56 ( .A(micro_hash_ucr_pipe57), .Y(micro_hash_ucr_pipe57_bF_buf3) );
BUFX4 BUFX4_57 ( .A(micro_hash_ucr_pipe57), .Y(micro_hash_ucr_pipe57_bF_buf2) );
BUFX4 BUFX4_58 ( .A(micro_hash_ucr_pipe57), .Y(micro_hash_ucr_pipe57_bF_buf1) );
BUFX4 BUFX4_59 ( .A(micro_hash_ucr_pipe57), .Y(micro_hash_ucr_pipe57_bF_buf0) );
BUFX4 BUFX4_60 ( .A(micro_hash_ucr_pipe58), .Y(micro_hash_ucr_pipe58_bF_buf3) );
BUFX4 BUFX4_61 ( .A(micro_hash_ucr_pipe58), .Y(micro_hash_ucr_pipe58_bF_buf2) );
BUFX4 BUFX4_62 ( .A(micro_hash_ucr_pipe58), .Y(micro_hash_ucr_pipe58_bF_buf1) );
BUFX4 BUFX4_63 ( .A(micro_hash_ucr_pipe58), .Y(micro_hash_ucr_pipe58_bF_buf0) );
BUFX4 BUFX4_64 ( .A(micro_hash_ucr_c_3_), .Y(micro_hash_ucr_c_3_bF_buf3_) );
BUFX4 BUFX4_65 ( .A(micro_hash_ucr_c_3_), .Y(micro_hash_ucr_c_3_bF_buf2_) );
BUFX4 BUFX4_66 ( .A(micro_hash_ucr_c_3_), .Y(micro_hash_ucr_c_3_bF_buf1_) );
BUFX4 BUFX4_67 ( .A(micro_hash_ucr_c_3_), .Y(micro_hash_ucr_c_3_bF_buf0_) );
BUFX4 BUFX4_68 ( .A(micro_hash_ucr_b_6_), .Y(micro_hash_ucr_b_6_bF_buf3_) );
BUFX4 BUFX4_69 ( .A(micro_hash_ucr_b_6_), .Y(micro_hash_ucr_b_6_bF_buf2_) );
BUFX4 BUFX4_70 ( .A(micro_hash_ucr_b_6_), .Y(micro_hash_ucr_b_6_bF_buf1_) );
BUFX4 BUFX4_71 ( .A(micro_hash_ucr_b_6_), .Y(micro_hash_ucr_b_6_bF_buf0_) );
BUFX4 BUFX4_72 ( .A(_4199_), .Y(_4199__bF_buf5) );
BUFX4 BUFX4_73 ( .A(_4199_), .Y(_4199__bF_buf4) );
BUFX4 BUFX4_74 ( .A(_4199_), .Y(_4199__bF_buf3) );
BUFX4 BUFX4_75 ( .A(_4199_), .Y(_4199__bF_buf2) );
BUFX4 BUFX4_76 ( .A(_4199_), .Y(_4199__bF_buf1) );
BUFX4 BUFX4_77 ( .A(_4199_), .Y(_4199__bF_buf0) );
BUFX4 BUFX4_78 ( .A(_4220_), .Y(_4220__bF_buf4) );
BUFX4 BUFX4_79 ( .A(_4220_), .Y(_4220__bF_buf3) );
BUFX4 BUFX4_80 ( .A(_4220_), .Y(_4220__bF_buf2) );
BUFX4 BUFX4_81 ( .A(_4220_), .Y(_4220__bF_buf1) );
BUFX4 BUFX4_82 ( .A(_4220_), .Y(_4220__bF_buf0) );
BUFX4 BUFX4_83 ( .A(_4217_), .Y(_4217__bF_buf3) );
BUFX4 BUFX4_84 ( .A(_4217_), .Y(_4217__bF_buf2) );
BUFX4 BUFX4_85 ( .A(_4217_), .Y(_4217__bF_buf1) );
BUFX4 BUFX4_86 ( .A(_4217_), .Y(_4217__bF_buf0) );
BUFX4 BUFX4_87 ( .A(_2932_), .Y(_2932__bF_buf3) );
BUFX4 BUFX4_88 ( .A(_2932_), .Y(_2932__bF_buf2) );
BUFX4 BUFX4_89 ( .A(_2932_), .Y(_2932__bF_buf1) );
BUFX4 BUFX4_90 ( .A(_2932_), .Y(_2932__bF_buf0) );
BUFX4 BUFX4_91 ( .A(micro_hash_ucr_pipe20), .Y(micro_hash_ucr_pipe20_bF_buf3) );
BUFX4 BUFX4_92 ( .A(micro_hash_ucr_pipe20), .Y(micro_hash_ucr_pipe20_bF_buf2) );
BUFX4 BUFX4_93 ( .A(micro_hash_ucr_pipe20), .Y(micro_hash_ucr_pipe20_bF_buf1) );
BUFX4 BUFX4_94 ( .A(micro_hash_ucr_pipe20), .Y(micro_hash_ucr_pipe20_bF_buf0) );
BUFX4 BUFX4_95 ( .A(micro_hash_ucr_pipe22), .Y(micro_hash_ucr_pipe22_bF_buf3) );
BUFX4 BUFX4_96 ( .A(micro_hash_ucr_pipe22), .Y(micro_hash_ucr_pipe22_bF_buf2) );
BUFX4 BUFX4_97 ( .A(micro_hash_ucr_pipe22), .Y(micro_hash_ucr_pipe22_bF_buf1) );
BUFX4 BUFX4_98 ( .A(micro_hash_ucr_pipe22), .Y(micro_hash_ucr_pipe22_bF_buf0) );
BUFX4 BUFX4_99 ( .A(micro_hash_ucr_pipe24), .Y(micro_hash_ucr_pipe24_bF_buf3) );
BUFX4 BUFX4_100 ( .A(micro_hash_ucr_pipe24), .Y(micro_hash_ucr_pipe24_bF_buf2) );
BUFX4 BUFX4_101 ( .A(micro_hash_ucr_pipe24), .Y(micro_hash_ucr_pipe24_bF_buf1) );
BUFX4 BUFX4_102 ( .A(micro_hash_ucr_pipe24), .Y(micro_hash_ucr_pipe24_bF_buf0) );
BUFX4 BUFX4_103 ( .A(micro_hash_ucr_pipe25), .Y(micro_hash_ucr_pipe25_bF_buf3) );
BUFX4 BUFX4_104 ( .A(micro_hash_ucr_pipe25), .Y(micro_hash_ucr_pipe25_bF_buf2) );
BUFX4 BUFX4_105 ( .A(micro_hash_ucr_pipe25), .Y(micro_hash_ucr_pipe25_bF_buf1) );
BUFX4 BUFX4_106 ( .A(micro_hash_ucr_pipe25), .Y(micro_hash_ucr_pipe25_bF_buf0) );
BUFX4 BUFX4_107 ( .A(micro_hash_ucr_pipe26), .Y(micro_hash_ucr_pipe26_bF_buf3) );
BUFX4 BUFX4_108 ( .A(micro_hash_ucr_pipe26), .Y(micro_hash_ucr_pipe26_bF_buf2) );
BUFX4 BUFX4_109 ( .A(micro_hash_ucr_pipe26), .Y(micro_hash_ucr_pipe26_bF_buf1) );
BUFX4 BUFX4_110 ( .A(micro_hash_ucr_pipe26), .Y(micro_hash_ucr_pipe26_bF_buf0) );
BUFX4 BUFX4_111 ( .A(micro_hash_ucr_pipe27), .Y(micro_hash_ucr_pipe27_bF_buf3) );
BUFX4 BUFX4_112 ( .A(micro_hash_ucr_pipe27), .Y(micro_hash_ucr_pipe27_bF_buf2) );
BUFX4 BUFX4_113 ( .A(micro_hash_ucr_pipe27), .Y(micro_hash_ucr_pipe27_bF_buf1) );
BUFX4 BUFX4_114 ( .A(micro_hash_ucr_pipe27), .Y(micro_hash_ucr_pipe27_bF_buf0) );
BUFX4 BUFX4_115 ( .A(micro_hash_ucr_pipe28), .Y(micro_hash_ucr_pipe28_bF_buf3) );
BUFX4 BUFX4_116 ( .A(micro_hash_ucr_pipe28), .Y(micro_hash_ucr_pipe28_bF_buf2) );
BUFX4 BUFX4_117 ( .A(micro_hash_ucr_pipe28), .Y(micro_hash_ucr_pipe28_bF_buf1) );
BUFX4 BUFX4_118 ( .A(micro_hash_ucr_pipe28), .Y(micro_hash_ucr_pipe28_bF_buf0) );
BUFX4 BUFX4_119 ( .A(micro_hash_ucr_c_0_), .Y(micro_hash_ucr_c_0_bF_buf3_) );
BUFX4 BUFX4_120 ( .A(micro_hash_ucr_c_0_), .Y(micro_hash_ucr_c_0_bF_buf2_) );
BUFX4 BUFX4_121 ( .A(micro_hash_ucr_c_0_), .Y(micro_hash_ucr_c_0_bF_buf1_) );
BUFX4 BUFX4_122 ( .A(micro_hash_ucr_c_0_), .Y(micro_hash_ucr_c_0_bF_buf0_) );
BUFX4 BUFX4_123 ( .A(micro_hash_ucr_b_3_), .Y(micro_hash_ucr_b_3_bF_buf3_) );
BUFX4 BUFX4_124 ( .A(micro_hash_ucr_b_3_), .Y(micro_hash_ucr_b_3_bF_buf2_) );
BUFX4 BUFX4_125 ( .A(micro_hash_ucr_b_3_), .Y(micro_hash_ucr_b_3_bF_buf1_) );
BUFX4 BUFX4_126 ( .A(micro_hash_ucr_b_3_), .Y(micro_hash_ucr_b_3_bF_buf0_) );
BUFX4 BUFX4_127 ( .A(_826_), .Y(_826__bF_buf3) );
BUFX4 BUFX4_128 ( .A(_826_), .Y(_826__bF_buf2) );
BUFX4 BUFX4_129 ( .A(_826_), .Y(_826__bF_buf1) );
BUFX4 BUFX4_130 ( .A(_826_), .Y(_826__bF_buf0) );
BUFX4 BUFX4_131 ( .A(micro_hash_ucr_a_6_), .Y(micro_hash_ucr_a_6_bF_buf3_) );
BUFX4 BUFX4_132 ( .A(micro_hash_ucr_a_6_), .Y(micro_hash_ucr_a_6_bF_buf2_) );
BUFX4 BUFX4_133 ( .A(micro_hash_ucr_a_6_), .Y(micro_hash_ucr_a_6_bF_buf1_) );
BUFX4 BUFX4_134 ( .A(micro_hash_ucr_a_6_), .Y(micro_hash_ucr_a_6_bF_buf0_) );
BUFX4 BUFX4_135 ( .A(_1665_), .Y(_1665__bF_buf3) );
BUFX4 BUFX4_136 ( .A(_1665_), .Y(_1665__bF_buf2) );
BUFX4 BUFX4_137 ( .A(_1665_), .Y(_1665__bF_buf1) );
BUFX4 BUFX4_138 ( .A(_1665_), .Y(_1665__bF_buf0) );
BUFX4 BUFX4_139 ( .A(_4214_), .Y(_4214__bF_buf4) );
BUFX4 BUFX4_140 ( .A(_4214_), .Y(_4214__bF_buf3) );
BUFX4 BUFX4_141 ( .A(_4214_), .Y(_4214__bF_buf2) );
BUFX4 BUFX4_142 ( .A(_4214_), .Y(_4214__bF_buf1) );
BUFX4 BUFX4_143 ( .A(_4214_), .Y(_4214__bF_buf0) );
BUFX4 BUFX4_144 ( .A(micro_hash_ucr_b_0_), .Y(micro_hash_ucr_b_0_bF_buf3_) );
BUFX4 BUFX4_145 ( .A(micro_hash_ucr_b_0_), .Y(micro_hash_ucr_b_0_bF_buf2_) );
BUFX4 BUFX4_146 ( .A(micro_hash_ucr_b_0_), .Y(micro_hash_ucr_b_0_bF_buf1_) );
BUFX4 BUFX4_147 ( .A(micro_hash_ucr_b_0_), .Y(micro_hash_ucr_b_0_bF_buf0_) );
BUFX4 BUFX4_148 ( .A(_823_), .Y(_823__bF_buf3) );
BUFX4 BUFX4_149 ( .A(_823_), .Y(_823__bF_buf2) );
BUFX4 BUFX4_150 ( .A(_823_), .Y(_823__bF_buf1) );
BUFX4 BUFX4_151 ( .A(_823_), .Y(_823__bF_buf0) );
BUFX4 BUFX4_152 ( .A(micro_hash_ucr_a_3_), .Y(micro_hash_ucr_a_3_bF_buf3_) );
BUFX4 BUFX4_153 ( .A(micro_hash_ucr_a_3_), .Y(micro_hash_ucr_a_3_bF_buf2_) );
BUFX4 BUFX4_154 ( .A(micro_hash_ucr_a_3_), .Y(micro_hash_ucr_a_3_bF_buf1_) );
BUFX4 BUFX4_155 ( .A(micro_hash_ucr_a_3_), .Y(micro_hash_ucr_a_3_bF_buf0_) );
BUFX4 BUFX4_156 ( .A(_3138_), .Y(_3138__bF_buf3) );
BUFX4 BUFX4_157 ( .A(_3138_), .Y(_3138__bF_buf2) );
BUFX4 BUFX4_158 ( .A(_3138_), .Y(_3138__bF_buf1) );
BUFX4 BUFX4_159 ( .A(_3138_), .Y(_3138__bF_buf0) );
BUFX4 BUFX4_160 ( .A(_4211_), .Y(_4211__bF_buf4) );
BUFX4 BUFX4_161 ( .A(_4211_), .Y(_4211__bF_buf3) );
BUFX4 BUFX4_162 ( .A(_4211_), .Y(_4211__bF_buf2) );
BUFX4 BUFX4_163 ( .A(_4211_), .Y(_4211__bF_buf1) );
BUFX4 BUFX4_164 ( .A(_4211_), .Y(_4211__bF_buf0) );
BUFX4 BUFX4_165 ( .A(micro_hash_ucr_a_0_), .Y(micro_hash_ucr_a_0_bF_buf3_) );
BUFX4 BUFX4_166 ( .A(micro_hash_ucr_a_0_), .Y(micro_hash_ucr_a_0_bF_buf2_) );
BUFX4 BUFX4_167 ( .A(micro_hash_ucr_a_0_), .Y(micro_hash_ucr_a_0_bF_buf1_) );
BUFX4 BUFX4_168 ( .A(micro_hash_ucr_a_0_), .Y(micro_hash_ucr_a_0_bF_buf0_) );
CLKBUF1 CLKBUF1_1 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf83) );
CLKBUF1 CLKBUF1_2 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf82) );
CLKBUF1 CLKBUF1_3 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf81) );
CLKBUF1 CLKBUF1_4 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf80) );
CLKBUF1 CLKBUF1_5 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf79) );
CLKBUF1 CLKBUF1_6 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf78) );
CLKBUF1 CLKBUF1_7 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf77) );
CLKBUF1 CLKBUF1_8 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf76) );
CLKBUF1 CLKBUF1_9 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf75) );
CLKBUF1 CLKBUF1_10 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf74) );
CLKBUF1 CLKBUF1_11 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf73) );
CLKBUF1 CLKBUF1_12 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf72) );
CLKBUF1 CLKBUF1_13 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf71) );
CLKBUF1 CLKBUF1_14 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf70) );
CLKBUF1 CLKBUF1_15 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf69) );
CLKBUF1 CLKBUF1_16 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf68) );
CLKBUF1 CLKBUF1_17 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf67) );
CLKBUF1 CLKBUF1_18 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf66) );
CLKBUF1 CLKBUF1_19 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf65) );
CLKBUF1 CLKBUF1_20 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf64) );
CLKBUF1 CLKBUF1_21 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf63) );
CLKBUF1 CLKBUF1_22 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf62) );
CLKBUF1 CLKBUF1_23 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf61) );
CLKBUF1 CLKBUF1_24 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf60) );
CLKBUF1 CLKBUF1_25 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf59) );
CLKBUF1 CLKBUF1_26 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf58) );
CLKBUF1 CLKBUF1_27 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf57) );
CLKBUF1 CLKBUF1_28 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf56) );
CLKBUF1 CLKBUF1_29 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf55) );
CLKBUF1 CLKBUF1_30 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf54) );
CLKBUF1 CLKBUF1_31 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf53) );
CLKBUF1 CLKBUF1_32 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf52) );
CLKBUF1 CLKBUF1_33 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf51) );
CLKBUF1 CLKBUF1_34 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf50) );
CLKBUF1 CLKBUF1_35 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf49) );
CLKBUF1 CLKBUF1_36 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf48) );
CLKBUF1 CLKBUF1_37 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf47) );
CLKBUF1 CLKBUF1_38 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf46) );
CLKBUF1 CLKBUF1_39 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf45) );
CLKBUF1 CLKBUF1_40 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf44) );
CLKBUF1 CLKBUF1_41 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf43) );
CLKBUF1 CLKBUF1_42 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf42) );
CLKBUF1 CLKBUF1_43 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf41) );
CLKBUF1 CLKBUF1_44 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf40) );
CLKBUF1 CLKBUF1_45 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf39) );
CLKBUF1 CLKBUF1_46 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf38) );
CLKBUF1 CLKBUF1_47 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf37) );
CLKBUF1 CLKBUF1_48 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf36) );
CLKBUF1 CLKBUF1_49 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf35) );
CLKBUF1 CLKBUF1_50 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf34) );
CLKBUF1 CLKBUF1_51 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf33) );
CLKBUF1 CLKBUF1_52 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf32) );
CLKBUF1 CLKBUF1_53 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf31) );
CLKBUF1 CLKBUF1_54 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf30) );
CLKBUF1 CLKBUF1_55 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf29) );
CLKBUF1 CLKBUF1_56 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf28) );
CLKBUF1 CLKBUF1_57 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf27) );
CLKBUF1 CLKBUF1_58 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf26) );
CLKBUF1 CLKBUF1_59 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf25) );
CLKBUF1 CLKBUF1_60 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf24) );
CLKBUF1 CLKBUF1_61 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf23) );
CLKBUF1 CLKBUF1_62 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf22) );
CLKBUF1 CLKBUF1_63 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf21) );
CLKBUF1 CLKBUF1_64 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf20) );
CLKBUF1 CLKBUF1_65 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf19) );
CLKBUF1 CLKBUF1_66 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf18) );
CLKBUF1 CLKBUF1_67 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf17) );
CLKBUF1 CLKBUF1_68 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf16) );
CLKBUF1 CLKBUF1_69 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf15) );
CLKBUF1 CLKBUF1_70 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf14) );
CLKBUF1 CLKBUF1_71 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf13) );
CLKBUF1 CLKBUF1_72 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf12) );
CLKBUF1 CLKBUF1_73 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf11) );
CLKBUF1 CLKBUF1_74 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf10) );
CLKBUF1 CLKBUF1_75 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf9) );
CLKBUF1 CLKBUF1_76 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf8) );
CLKBUF1 CLKBUF1_77 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf7) );
CLKBUF1 CLKBUF1_78 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf6) );
CLKBUF1 CLKBUF1_79 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf5) );
CLKBUF1 CLKBUF1_80 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf4) );
CLKBUF1 CLKBUF1_81 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf3) );
CLKBUF1 CLKBUF1_82 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf2) );
CLKBUF1 CLKBUF1_83 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf1) );
CLKBUF1 CLKBUF1_84 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf0) );
BUFX4 BUFX4_169 ( .A(_2441_), .Y(_2441__bF_buf3) );
BUFX4 BUFX4_170 ( .A(_2441_), .Y(_2441__bF_buf2) );
BUFX4 BUFX4_171 ( .A(_2441_), .Y(_2441__bF_buf1) );
BUFX4 BUFX4_172 ( .A(_2441_), .Y(_2441__bF_buf0) );
BUFX4 BUFX4_173 ( .A(_2820_), .Y(_2820__bF_buf3) );
BUFX4 BUFX4_174 ( .A(_2820_), .Y(_2820__bF_buf2) );
BUFX4 BUFX4_175 ( .A(_2820_), .Y(_2820__bF_buf1) );
BUFX4 BUFX4_176 ( .A(_2820_), .Y(_2820__bF_buf0) );
BUFX4 BUFX4_177 ( .A(_4237_), .Y(_4237__bF_buf4) );
BUFX4 BUFX4_178 ( .A(_4237_), .Y(_4237__bF_buf3) );
BUFX4 BUFX4_179 ( .A(_4237_), .Y(_4237__bF_buf2) );
BUFX4 BUFX4_180 ( .A(_4237_), .Y(_4237__bF_buf1) );
BUFX4 BUFX4_181 ( .A(_4237_), .Y(_4237__bF_buf0) );
BUFX4 BUFX4_182 ( .A(_426_), .Y(_426__bF_buf3) );
BUFX4 BUFX4_183 ( .A(_426_), .Y(_426__bF_buf2) );
BUFX4 BUFX4_184 ( .A(_426_), .Y(_426__bF_buf1) );
BUFX4 BUFX4_185 ( .A(_426_), .Y(_426__bF_buf0) );
BUFX4 BUFX4_186 ( .A(_4234_), .Y(_4234__bF_buf3) );
BUFX4 BUFX4_187 ( .A(_4234_), .Y(_4234__bF_buf2) );
BUFX4 BUFX4_188 ( .A(_4234_), .Y(_4234__bF_buf1) );
BUFX4 BUFX4_189 ( .A(_4234_), .Y(_4234__bF_buf0) );
BUFX4 BUFX4_190 ( .A(_2811_), .Y(_2811__bF_buf3) );
BUFX4 BUFX4_191 ( .A(_2811_), .Y(_2811__bF_buf2) );
BUFX4 BUFX4_192 ( .A(_2811_), .Y(_2811__bF_buf1) );
BUFX4 BUFX4_193 ( .A(_2811_), .Y(_2811__bF_buf0) );
BUFX4 BUFX4_194 ( .A(_1679_), .Y(_1679__bF_buf3) );
BUFX4 BUFX4_195 ( .A(_1679_), .Y(_1679__bF_buf2) );
BUFX4 BUFX4_196 ( .A(_1679_), .Y(_1679__bF_buf1) );
BUFX4 BUFX4_197 ( .A(_1679_), .Y(_1679__bF_buf0) );
BUFX4 BUFX4_198 ( .A(_399_), .Y(_399__bF_buf3) );
BUFX4 BUFX4_199 ( .A(_399_), .Y(_399__bF_buf2) );
BUFX4 BUFX4_200 ( .A(_399_), .Y(_399__bF_buf1) );
BUFX4 BUFX4_201 ( .A(_399_), .Y(_399__bF_buf0) );
BUFX4 BUFX4_202 ( .A(_4228_), .Y(_4228__bF_buf4) );
BUFX4 BUFX4_203 ( .A(_4228_), .Y(_4228__bF_buf3) );
BUFX4 BUFX4_204 ( .A(_4228_), .Y(_4228__bF_buf2) );
BUFX4 BUFX4_205 ( .A(_4228_), .Y(_4228__bF_buf1) );
BUFX4 BUFX4_206 ( .A(_4228_), .Y(_4228__bF_buf0) );
BUFX4 BUFX4_207 ( .A(_4225_), .Y(_4225__bF_buf4) );
BUFX4 BUFX4_208 ( .A(_4225_), .Y(_4225__bF_buf3) );
BUFX4 BUFX4_209 ( .A(_4225_), .Y(_4225__bF_buf2) );
BUFX4 BUFX4_210 ( .A(_4225_), .Y(_4225__bF_buf1) );
BUFX4 BUFX4_211 ( .A(_4225_), .Y(_4225__bF_buf0) );
BUFX4 BUFX4_212 ( .A(_3246_), .Y(_3246__bF_buf3) );
BUFX4 BUFX4_213 ( .A(_3246_), .Y(_3246__bF_buf2) );
BUFX4 BUFX4_214 ( .A(_3246_), .Y(_3246__bF_buf1) );
BUFX4 BUFX4_215 ( .A(_3246_), .Y(_3246__bF_buf0) );
BUFX4 BUFX4_216 ( .A(micro_hash_ucr_pipe70), .Y(micro_hash_ucr_pipe70_bF_buf3) );
BUFX4 BUFX4_217 ( .A(micro_hash_ucr_pipe70), .Y(micro_hash_ucr_pipe70_bF_buf2) );
BUFX4 BUFX4_218 ( .A(micro_hash_ucr_pipe70), .Y(micro_hash_ucr_pipe70_bF_buf1) );
BUFX4 BUFX4_219 ( .A(micro_hash_ucr_pipe70), .Y(micro_hash_ucr_pipe70_bF_buf0) );
BUFX4 BUFX4_220 ( .A(_317_), .Y(_317__bF_buf3) );
BUFX4 BUFX4_221 ( .A(_317_), .Y(_317__bF_buf2) );
BUFX4 BUFX4_222 ( .A(_317_), .Y(_317__bF_buf1) );
BUFX4 BUFX4_223 ( .A(_317_), .Y(_317__bF_buf0) );
BUFX4 BUFX4_224 ( .A(_1673_), .Y(_1673__bF_buf3) );
BUFX4 BUFX4_225 ( .A(_1673_), .Y(_1673__bF_buf2) );
BUFX4 BUFX4_226 ( .A(_1673_), .Y(_1673__bF_buf1) );
BUFX4 BUFX4_227 ( .A(_1673_), .Y(_1673__bF_buf0) );
BUFX4 BUFX4_228 ( .A(_296_), .Y(_296__bF_buf4) );
BUFX4 BUFX4_229 ( .A(_296_), .Y(_296__bF_buf3) );
BUFX4 BUFX4_230 ( .A(_296_), .Y(_296__bF_buf2) );
BUFX4 BUFX4_231 ( .A(_296_), .Y(_296__bF_buf1) );
BUFX4 BUFX4_232 ( .A(_296_), .Y(_296__bF_buf0) );
BUFX4 BUFX4_233 ( .A(_4219_), .Y(_4219__bF_buf4) );
BUFX4 BUFX4_234 ( .A(_4219_), .Y(_4219__bF_buf3) );
BUFX4 BUFX4_235 ( .A(_4219_), .Y(_4219__bF_buf2) );
BUFX4 BUFX4_236 ( .A(_4219_), .Y(_4219__bF_buf1) );
BUFX4 BUFX4_237 ( .A(_4219_), .Y(_4219__bF_buf0) );
BUFX4 BUFX4_238 ( .A(_220_), .Y(_220__bF_buf4) );
BUFX4 BUFX4_239 ( .A(_220_), .Y(_220__bF_buf3) );
BUFX4 BUFX4_240 ( .A(_220_), .Y(_220__bF_buf2) );
BUFX4 BUFX4_241 ( .A(_220_), .Y(_220__bF_buf1) );
BUFX4 BUFX4_242 ( .A(_220_), .Y(_220__bF_buf0) );
BUFX4 BUFX4_243 ( .A(_2514_), .Y(_2514__bF_buf3) );
BUFX4 BUFX4_244 ( .A(_2514_), .Y(_2514__bF_buf2) );
BUFX4 BUFX4_245 ( .A(_2514_), .Y(_2514__bF_buf1) );
BUFX4 BUFX4_246 ( .A(_2514_), .Y(_2514__bF_buf0) );
BUFX4 BUFX4_247 ( .A(_3892_), .Y(_3892__bF_buf3) );
BUFX4 BUFX4_248 ( .A(_3892_), .Y(_3892__bF_buf2) );
BUFX4 BUFX4_249 ( .A(_3892_), .Y(_3892__bF_buf1) );
BUFX4 BUFX4_250 ( .A(_3892_), .Y(_3892__bF_buf0) );
BUFX4 BUFX4_251 ( .A(micro_hash_ucr_pipe40), .Y(micro_hash_ucr_pipe40_bF_buf4) );
BUFX4 BUFX4_252 ( .A(micro_hash_ucr_pipe40), .Y(micro_hash_ucr_pipe40_bF_buf3) );
BUFX4 BUFX4_253 ( .A(micro_hash_ucr_pipe40), .Y(micro_hash_ucr_pipe40_bF_buf2) );
BUFX4 BUFX4_254 ( .A(micro_hash_ucr_pipe40), .Y(micro_hash_ucr_pipe40_bF_buf1) );
BUFX4 BUFX4_255 ( .A(micro_hash_ucr_pipe40), .Y(micro_hash_ucr_pipe40_bF_buf0) );
BUFX4 BUFX4_256 ( .A(micro_hash_ucr_pipe41), .Y(micro_hash_ucr_pipe41_bF_buf3) );
BUFX4 BUFX4_257 ( .A(micro_hash_ucr_pipe41), .Y(micro_hash_ucr_pipe41_bF_buf2) );
BUFX4 BUFX4_258 ( .A(micro_hash_ucr_pipe41), .Y(micro_hash_ucr_pipe41_bF_buf1) );
BUFX4 BUFX4_259 ( .A(micro_hash_ucr_pipe41), .Y(micro_hash_ucr_pipe41_bF_buf0) );
BUFX4 BUFX4_260 ( .A(micro_hash_ucr_pipe42), .Y(micro_hash_ucr_pipe42_bF_buf4) );
BUFX4 BUFX4_261 ( .A(micro_hash_ucr_pipe42), .Y(micro_hash_ucr_pipe42_bF_buf3) );
BUFX4 BUFX4_262 ( .A(micro_hash_ucr_pipe42), .Y(micro_hash_ucr_pipe42_bF_buf2) );
BUFX4 BUFX4_263 ( .A(micro_hash_ucr_pipe42), .Y(micro_hash_ucr_pipe42_bF_buf1) );
BUFX4 BUFX4_264 ( .A(micro_hash_ucr_pipe42), .Y(micro_hash_ucr_pipe42_bF_buf0) );
BUFX4 BUFX4_265 ( .A(micro_hash_ucr_pipe44), .Y(micro_hash_ucr_pipe44_bF_buf3) );
BUFX4 BUFX4_266 ( .A(micro_hash_ucr_pipe44), .Y(micro_hash_ucr_pipe44_bF_buf2) );
BUFX4 BUFX4_267 ( .A(micro_hash_ucr_pipe44), .Y(micro_hash_ucr_pipe44_bF_buf1) );
BUFX4 BUFX4_268 ( .A(micro_hash_ucr_pipe44), .Y(micro_hash_ucr_pipe44_bF_buf0) );
BUFX4 BUFX4_269 ( .A(micro_hash_ucr_pipe46), .Y(micro_hash_ucr_pipe46_bF_buf4) );
BUFX4 BUFX4_270 ( .A(micro_hash_ucr_pipe46), .Y(micro_hash_ucr_pipe46_bF_buf3) );
BUFX4 BUFX4_271 ( .A(micro_hash_ucr_pipe46), .Y(micro_hash_ucr_pipe46_bF_buf2) );
BUFX4 BUFX4_272 ( .A(micro_hash_ucr_pipe46), .Y(micro_hash_ucr_pipe46_bF_buf1) );
BUFX4 BUFX4_273 ( .A(micro_hash_ucr_pipe46), .Y(micro_hash_ucr_pipe46_bF_buf0) );
BUFX4 BUFX4_274 ( .A(micro_hash_ucr_pipe48), .Y(micro_hash_ucr_pipe48_bF_buf4) );
BUFX4 BUFX4_275 ( .A(micro_hash_ucr_pipe48), .Y(micro_hash_ucr_pipe48_bF_buf3) );
BUFX4 BUFX4_276 ( .A(micro_hash_ucr_pipe48), .Y(micro_hash_ucr_pipe48_bF_buf2) );
BUFX4 BUFX4_277 ( .A(micro_hash_ucr_pipe48), .Y(micro_hash_ucr_pipe48_bF_buf1) );
BUFX4 BUFX4_278 ( .A(micro_hash_ucr_pipe48), .Y(micro_hash_ucr_pipe48_bF_buf0) );
BUFX4 BUFX4_279 ( .A(micro_hash_ucr_pipe49), .Y(micro_hash_ucr_pipe49_bF_buf3) );
BUFX4 BUFX4_280 ( .A(micro_hash_ucr_pipe49), .Y(micro_hash_ucr_pipe49_bF_buf2) );
BUFX4 BUFX4_281 ( .A(micro_hash_ucr_pipe49), .Y(micro_hash_ucr_pipe49_bF_buf1) );
BUFX4 BUFX4_282 ( .A(micro_hash_ucr_pipe49), .Y(micro_hash_ucr_pipe49_bF_buf0) );
BUFX4 BUFX4_283 ( .A(micro_hash_ucr_c_2_), .Y(micro_hash_ucr_c_2_bF_buf3_) );
BUFX4 BUFX4_284 ( .A(micro_hash_ucr_c_2_), .Y(micro_hash_ucr_c_2_bF_buf2_) );
BUFX4 BUFX4_285 ( .A(micro_hash_ucr_c_2_), .Y(micro_hash_ucr_c_2_bF_buf1_) );
BUFX4 BUFX4_286 ( .A(micro_hash_ucr_c_2_), .Y(micro_hash_ucr_c_2_bF_buf0_) );
BUFX4 BUFX4_287 ( .A(micro_hash_ucr_b_5_), .Y(micro_hash_ucr_b_5_bF_buf3_) );
BUFX4 BUFX4_288 ( .A(micro_hash_ucr_b_5_), .Y(micro_hash_ucr_b_5_bF_buf2_) );
BUFX4 BUFX4_289 ( .A(micro_hash_ucr_b_5_), .Y(micro_hash_ucr_b_5_bF_buf1_) );
BUFX4 BUFX4_290 ( .A(micro_hash_ucr_b_5_), .Y(micro_hash_ucr_b_5_bF_buf0_) );
BUFX4 BUFX4_291 ( .A(_255_), .Y(_255__bF_buf3) );
BUFX4 BUFX4_292 ( .A(_255_), .Y(_255__bF_buf2) );
BUFX4 BUFX4_293 ( .A(_255_), .Y(_255__bF_buf1) );
BUFX4 BUFX4_294 ( .A(_255_), .Y(_255__bF_buf0) );
BUFX4 BUFX4_295 ( .A(_1438_), .Y(_1438__bF_buf5) );
BUFX4 BUFX4_296 ( .A(_1438_), .Y(_1438__bF_buf4) );
BUFX4 BUFX4_297 ( .A(_1438_), .Y(_1438__bF_buf3) );
BUFX4 BUFX4_298 ( .A(_1438_), .Y(_1438__bF_buf2) );
BUFX4 BUFX4_299 ( .A(_1438_), .Y(_1438__bF_buf1) );
BUFX4 BUFX4_300 ( .A(_1438_), .Y(_1438__bF_buf0) );
BUFX4 BUFX4_301 ( .A(micro_hash_ucr_pipe12), .Y(micro_hash_ucr_pipe12_bF_buf3) );
BUFX4 BUFX4_302 ( .A(micro_hash_ucr_pipe12), .Y(micro_hash_ucr_pipe12_bF_buf2) );
BUFX4 BUFX4_303 ( .A(micro_hash_ucr_pipe12), .Y(micro_hash_ucr_pipe12_bF_buf1) );
BUFX4 BUFX4_304 ( .A(micro_hash_ucr_pipe12), .Y(micro_hash_ucr_pipe12_bF_buf0) );
BUFX4 BUFX4_305 ( .A(micro_hash_ucr_pipe18), .Y(micro_hash_ucr_pipe18_bF_buf4) );
BUFX4 BUFX4_306 ( .A(micro_hash_ucr_pipe18), .Y(micro_hash_ucr_pipe18_bF_buf3) );
BUFX4 BUFX4_307 ( .A(micro_hash_ucr_pipe18), .Y(micro_hash_ucr_pipe18_bF_buf2) );
BUFX4 BUFX4_308 ( .A(micro_hash_ucr_pipe18), .Y(micro_hash_ucr_pipe18_bF_buf1) );
BUFX4 BUFX4_309 ( .A(micro_hash_ucr_pipe18), .Y(micro_hash_ucr_pipe18_bF_buf0) );
BUFX4 BUFX4_310 ( .A(micro_hash_ucr_b_2_), .Y(micro_hash_ucr_b_2_bF_buf3_) );
BUFX4 BUFX4_311 ( .A(micro_hash_ucr_b_2_), .Y(micro_hash_ucr_b_2_bF_buf2_) );
BUFX4 BUFX4_312 ( .A(micro_hash_ucr_b_2_), .Y(micro_hash_ucr_b_2_bF_buf1_) );
BUFX4 BUFX4_313 ( .A(micro_hash_ucr_b_2_), .Y(micro_hash_ucr_b_2_bF_buf0_) );
BUFX4 BUFX4_314 ( .A(micro_hash_ucr_a_5_), .Y(micro_hash_ucr_a_5_bF_buf3_) );
BUFX4 BUFX4_315 ( .A(micro_hash_ucr_a_5_), .Y(micro_hash_ucr_a_5_bF_buf2_) );
BUFX4 BUFX4_316 ( .A(micro_hash_ucr_a_5_), .Y(micro_hash_ucr_a_5_bF_buf1_) );
BUFX4 BUFX4_317 ( .A(micro_hash_ucr_a_5_), .Y(micro_hash_ucr_a_5_bF_buf0_) );
BUFX4 BUFX4_318 ( .A(_2487_), .Y(_2487__bF_buf3) );
BUFX4 BUFX4_319 ( .A(_2487_), .Y(_2487__bF_buf2) );
BUFX4 BUFX4_320 ( .A(_2487_), .Y(_2487__bF_buf1) );
BUFX4 BUFX4_321 ( .A(_2487_), .Y(_2487__bF_buf0) );
BUFX4 BUFX4_322 ( .A(_249_), .Y(_249__bF_buf3) );
BUFX4 BUFX4_323 ( .A(_249_), .Y(_249__bF_buf2) );
BUFX4 BUFX4_324 ( .A(_249_), .Y(_249__bF_buf1) );
BUFX4 BUFX4_325 ( .A(_249_), .Y(_249__bF_buf0) );
BUFX4 BUFX4_326 ( .A(micro_hash_ucr_a_2_), .Y(micro_hash_ucr_a_2_bF_buf4_) );
BUFX4 BUFX4_327 ( .A(micro_hash_ucr_a_2_), .Y(micro_hash_ucr_a_2_bF_buf3_) );
BUFX4 BUFX4_328 ( .A(micro_hash_ucr_a_2_), .Y(micro_hash_ucr_a_2_bF_buf2_) );
BUFX4 BUFX4_329 ( .A(micro_hash_ucr_a_2_), .Y(micro_hash_ucr_a_2_bF_buf1_) );
BUFX4 BUFX4_330 ( .A(micro_hash_ucr_a_2_), .Y(micro_hash_ucr_a_2_bF_buf0_) );
BUFX4 BUFX4_331 ( .A(_4210_), .Y(_4210__bF_buf4) );
BUFX4 BUFX4_332 ( .A(_4210_), .Y(_4210__bF_buf3) );
BUFX4 BUFX4_333 ( .A(_4210_), .Y(_4210__bF_buf2) );
BUFX4 BUFX4_334 ( .A(_4210_), .Y(_4210__bF_buf1) );
BUFX4 BUFX4_335 ( .A(_4210_), .Y(_4210__bF_buf0) );
BUFX4 BUFX4_336 ( .A(_0_), .Y(_0__bF_buf8) );
BUFX4 BUFX4_337 ( .A(_0_), .Y(_0__bF_buf7) );
BUFX4 BUFX4_338 ( .A(_0_), .Y(_0__bF_buf6) );
BUFX4 BUFX4_339 ( .A(_0_), .Y(_0__bF_buf5) );
BUFX4 BUFX4_340 ( .A(_0_), .Y(_0__bF_buf4) );
BUFX4 BUFX4_341 ( .A(_0_), .Y(_0__bF_buf3) );
BUFX4 BUFX4_342 ( .A(_0_), .Y(_0__bF_buf2) );
BUFX4 BUFX4_343 ( .A(_0_), .Y(_0__bF_buf1) );
BUFX4 BUFX4_344 ( .A(_0_), .Y(_0__bF_buf0) );
BUFX4 BUFX4_345 ( .A(_4207_), .Y(_4207__bF_buf4) );
BUFX4 BUFX4_346 ( .A(_4207_), .Y(_4207__bF_buf3) );
BUFX4 BUFX4_347 ( .A(_4207_), .Y(_4207__bF_buf2) );
BUFX4 BUFX4_348 ( .A(_4207_), .Y(_4207__bF_buf1) );
BUFX4 BUFX4_349 ( .A(_4207_), .Y(_4207__bF_buf0) );
BUFX4 BUFX4_350 ( .A(_4283__hier0_bF_buf2), .Y(_4283__bF_buf42) );
BUFX4 BUFX4_351 ( .A(_4283__hier0_bF_buf2), .Y(_4283__bF_buf41) );
BUFX4 BUFX4_352 ( .A(_4283__hier0_bF_buf0), .Y(_4283__bF_buf40) );
BUFX4 BUFX4_353 ( .A(_4283__hier0_bF_buf3), .Y(_4283__bF_buf39) );
BUFX4 BUFX4_354 ( .A(_4283__hier0_bF_buf4), .Y(_4283__bF_buf38) );
BUFX4 BUFX4_355 ( .A(_4283__hier0_bF_buf2), .Y(_4283__bF_buf37) );
BUFX4 BUFX4_356 ( .A(_4283__hier0_bF_buf0), .Y(_4283__bF_buf36) );
BUFX4 BUFX4_357 ( .A(_4283__hier0_bF_buf3), .Y(_4283__bF_buf35) );
BUFX4 BUFX4_358 ( .A(_4283__hier0_bF_buf1), .Y(_4283__bF_buf34) );
BUFX4 BUFX4_359 ( .A(_4283__hier0_bF_buf5), .Y(_4283__bF_buf33) );
BUFX4 BUFX4_360 ( .A(_4283__hier0_bF_buf4), .Y(_4283__bF_buf32) );
BUFX4 BUFX4_361 ( .A(_4283__hier0_bF_buf0), .Y(_4283__bF_buf31) );
BUFX4 BUFX4_362 ( .A(_4283__hier0_bF_buf5), .Y(_4283__bF_buf30) );
BUFX4 BUFX4_363 ( .A(_4283__hier0_bF_buf3), .Y(_4283__bF_buf29) );
BUFX4 BUFX4_364 ( .A(_4283__hier0_bF_buf2), .Y(_4283__bF_buf28) );
BUFX4 BUFX4_365 ( .A(_4283__hier0_bF_buf3), .Y(_4283__bF_buf27) );
BUFX4 BUFX4_366 ( .A(_4283__hier0_bF_buf5), .Y(_4283__bF_buf26) );
BUFX4 BUFX4_367 ( .A(_4283__hier0_bF_buf0), .Y(_4283__bF_buf25) );
BUFX4 BUFX4_368 ( .A(_4283__hier0_bF_buf4), .Y(_4283__bF_buf24) );
BUFX4 BUFX4_369 ( .A(_4283__hier0_bF_buf5), .Y(_4283__bF_buf23) );
BUFX4 BUFX4_370 ( .A(_4283__hier0_bF_buf1), .Y(_4283__bF_buf22) );
BUFX4 BUFX4_371 ( .A(_4283__hier0_bF_buf4), .Y(_4283__bF_buf21) );
BUFX4 BUFX4_372 ( .A(_4283__hier0_bF_buf1), .Y(_4283__bF_buf20) );
BUFX4 BUFX4_373 ( .A(_4283__hier0_bF_buf5), .Y(_4283__bF_buf19) );
BUFX4 BUFX4_374 ( .A(_4283__hier0_bF_buf1), .Y(_4283__bF_buf18) );
BUFX4 BUFX4_375 ( .A(_4283__hier0_bF_buf4), .Y(_4283__bF_buf17) );
BUFX4 BUFX4_376 ( .A(_4283__hier0_bF_buf4), .Y(_4283__bF_buf16) );
BUFX4 BUFX4_377 ( .A(_4283__hier0_bF_buf2), .Y(_4283__bF_buf15) );
BUFX4 BUFX4_378 ( .A(_4283__hier0_bF_buf1), .Y(_4283__bF_buf14) );
BUFX4 BUFX4_379 ( .A(_4283__hier0_bF_buf5), .Y(_4283__bF_buf13) );
BUFX4 BUFX4_380 ( .A(_4283__hier0_bF_buf2), .Y(_4283__bF_buf12) );
BUFX4 BUFX4_381 ( .A(_4283__hier0_bF_buf5), .Y(_4283__bF_buf11) );
BUFX4 BUFX4_382 ( .A(_4283__hier0_bF_buf3), .Y(_4283__bF_buf10) );
BUFX4 BUFX4_383 ( .A(_4283__hier0_bF_buf0), .Y(_4283__bF_buf9) );
BUFX4 BUFX4_384 ( .A(_4283__hier0_bF_buf5), .Y(_4283__bF_buf8) );
BUFX4 BUFX4_385 ( .A(_4283__hier0_bF_buf0), .Y(_4283__bF_buf7) );
BUFX4 BUFX4_386 ( .A(_4283__hier0_bF_buf2), .Y(_4283__bF_buf6) );
BUFX4 BUFX4_387 ( .A(_4283__hier0_bF_buf1), .Y(_4283__bF_buf5) );
BUFX4 BUFX4_388 ( .A(_4283__hier0_bF_buf1), .Y(_4283__bF_buf4) );
BUFX4 BUFX4_389 ( .A(_4283__hier0_bF_buf4), .Y(_4283__bF_buf3) );
BUFX4 BUFX4_390 ( .A(_4283__hier0_bF_buf3), .Y(_4283__bF_buf2) );
BUFX4 BUFX4_391 ( .A(_4283__hier0_bF_buf3), .Y(_4283__bF_buf1) );
BUFX4 BUFX4_392 ( .A(_4283__hier0_bF_buf0), .Y(_4283__bF_buf0) );
BUFX4 BUFX4_393 ( .A(_3037_), .Y(_3037__bF_buf3) );
BUFX4 BUFX4_394 ( .A(_3037_), .Y(_3037__bF_buf2) );
BUFX4 BUFX4_395 ( .A(_3037_), .Y(_3037__bF_buf1) );
BUFX4 BUFX4_396 ( .A(_3037_), .Y(_3037__bF_buf0) );
BUFX4 BUFX4_397 ( .A(_278_), .Y(_278__bF_buf3) );
BUFX4 BUFX4_398 ( .A(_278_), .Y(_278__bF_buf2) );
BUFX4 BUFX4_399 ( .A(_278_), .Y(_278__bF_buf1) );
BUFX4 BUFX4_400 ( .A(_278_), .Y(_278__bF_buf0) );
BUFX4 BUFX4_401 ( .A(_4239_), .Y(_4239__bF_buf4) );
BUFX4 BUFX4_402 ( .A(_4239_), .Y(_4239__bF_buf3) );
BUFX4 BUFX4_403 ( .A(_4239_), .Y(_4239__bF_buf2) );
BUFX4 BUFX4_404 ( .A(_4239_), .Y(_4239__bF_buf1) );
BUFX4 BUFX4_405 ( .A(_4239_), .Y(_4239__bF_buf0) );
BUFX4 BUFX4_406 ( .A(_2190_), .Y(_2190__bF_buf4) );
BUFX4 BUFX4_407 ( .A(_2190_), .Y(_2190__bF_buf3) );
BUFX4 BUFX4_408 ( .A(_2190_), .Y(_2190__bF_buf2) );
BUFX4 BUFX4_409 ( .A(_2190_), .Y(_2190__bF_buf1) );
BUFX4 BUFX4_410 ( .A(_2190_), .Y(_2190__bF_buf0) );
BUFX4 BUFX4_411 ( .A(_4201_), .Y(_4201__bF_buf3) );
BUFX4 BUFX4_412 ( .A(_4201_), .Y(_4201__bF_buf2) );
BUFX4 BUFX4_413 ( .A(_4201_), .Y(_4201__bF_buf1) );
BUFX4 BUFX4_414 ( .A(_4201_), .Y(_4201__bF_buf0) );
BUFX4 BUFX4_415 ( .A(_4236_), .Y(_4236__bF_buf3) );
BUFX4 BUFX4_416 ( .A(_4236_), .Y(_4236__bF_buf2) );
BUFX4 BUFX4_417 ( .A(_4236_), .Y(_4236__bF_buf1) );
BUFX4 BUFX4_418 ( .A(_4236_), .Y(_4236__bF_buf0) );
BUFX4 BUFX4_419 ( .A(_3354_), .Y(_3354__bF_buf3) );
BUFX4 BUFX4_420 ( .A(_3354_), .Y(_3354__bF_buf2) );
BUFX4 BUFX4_421 ( .A(_3354_), .Y(_3354__bF_buf1) );
BUFX4 BUFX4_422 ( .A(_3354_), .Y(_3354__bF_buf0) );
BUFX4 BUFX4_423 ( .A(_845_), .Y(_845__bF_buf3) );
BUFX4 BUFX4_424 ( .A(_845_), .Y(_845__bF_buf2) );
BUFX4 BUFX4_425 ( .A(_845_), .Y(_845__bF_buf1) );
BUFX4 BUFX4_426 ( .A(_845_), .Y(_845__bF_buf0) );
BUFX4 BUFX4_427 ( .A(_425_), .Y(_425__bF_buf5) );
BUFX4 BUFX4_428 ( .A(_425_), .Y(_425__bF_buf4) );
BUFX4 BUFX4_429 ( .A(_425_), .Y(_425__bF_buf3) );
BUFX4 BUFX4_430 ( .A(_425_), .Y(_425__bF_buf2) );
BUFX4 BUFX4_431 ( .A(_425_), .Y(_425__bF_buf1) );
BUFX4 BUFX4_432 ( .A(_425_), .Y(_425__bF_buf0) );
BUFX4 BUFX4_433 ( .A(_2184_), .Y(_2184__bF_buf3) );
BUFX4 BUFX4_434 ( .A(_2184_), .Y(_2184__bF_buf2) );
BUFX4 BUFX4_435 ( .A(_2184_), .Y(_2184__bF_buf1) );
BUFX4 BUFX4_436 ( .A(_2184_), .Y(_2184__bF_buf0) );
BUFX4 BUFX4_437 ( .A(_4233_), .Y(_4233__bF_buf4) );
BUFX4 BUFX4_438 ( .A(_4233_), .Y(_4233__bF_buf3) );
BUFX4 BUFX4_439 ( .A(_4233_), .Y(_4233__bF_buf2) );
BUFX4 BUFX4_440 ( .A(_4233_), .Y(_4233__bF_buf1) );
BUFX4 BUFX4_441 ( .A(_4233_), .Y(_4233__bF_buf0) );
BUFX4 BUFX4_442 ( .A(_2813_), .Y(_2813__bF_buf3) );
BUFX4 BUFX4_443 ( .A(_2813_), .Y(_2813__bF_buf2) );
BUFX4 BUFX4_444 ( .A(_2813_), .Y(_2813__bF_buf1) );
BUFX4 BUFX4_445 ( .A(_2813_), .Y(_2813__bF_buf0) );
BUFX4 BUFX4_446 ( .A(_4230_), .Y(_4230__bF_buf4) );
BUFX4 BUFX4_447 ( .A(_4230_), .Y(_4230__bF_buf3) );
BUFX4 BUFX4_448 ( .A(_4230_), .Y(_4230__bF_buf2) );
BUFX4 BUFX4_449 ( .A(_4230_), .Y(_4230__bF_buf1) );
BUFX4 BUFX4_450 ( .A(_4230_), .Y(_4230__bF_buf0) );
BUFX4 BUFX4_451 ( .A(comparador_valid), .Y(comparador_valid_bF_buf4) );
BUFX4 BUFX4_452 ( .A(comparador_valid), .Y(comparador_valid_bF_buf3) );
BUFX4 BUFX4_453 ( .A(comparador_valid), .Y(comparador_valid_bF_buf2) );
BUFX4 BUFX4_454 ( .A(comparador_valid), .Y(comparador_valid_bF_buf1) );
BUFX4 BUFX4_455 ( .A(comparador_valid), .Y(comparador_valid_bF_buf0) );
BUFX4 BUFX4_456 ( .A(_1678_), .Y(_1678__bF_buf5) );
BUFX4 BUFX4_457 ( .A(_1678_), .Y(_1678__bF_buf4) );
BUFX4 BUFX4_458 ( .A(_1678_), .Y(_1678__bF_buf3) );
BUFX4 BUFX4_459 ( .A(_1678_), .Y(_1678__bF_buf2) );
BUFX4 BUFX4_460 ( .A(_1678_), .Y(_1678__bF_buf1) );
BUFX4 BUFX4_461 ( .A(_1678_), .Y(_1678__bF_buf0) );
BUFX4 BUFX4_462 ( .A(_742_), .Y(_742__bF_buf3) );
BUFX4 BUFX4_463 ( .A(_742_), .Y(_742__bF_buf2) );
BUFX4 BUFX4_464 ( .A(_742_), .Y(_742__bF_buf1) );
BUFX4 BUFX4_465 ( .A(_742_), .Y(_742__bF_buf0) );
BUFX4 BUFX4_466 ( .A(_131_), .Y(_131__bF_buf13) );
BUFX4 BUFX4_467 ( .A(_131_), .Y(_131__bF_buf12) );
BUFX4 BUFX4_468 ( .A(_131_), .Y(_131__bF_buf11) );
BUFX4 BUFX4_469 ( .A(_131_), .Y(_131__bF_buf10) );
BUFX4 BUFX4_470 ( .A(_131_), .Y(_131__bF_buf9) );
BUFX4 BUFX4_471 ( .A(_131_), .Y(_131__bF_buf8) );
BUFX4 BUFX4_472 ( .A(_131_), .Y(_131__bF_buf7) );
BUFX4 BUFX4_473 ( .A(_131_), .Y(_131__bF_buf6) );
BUFX4 BUFX4_474 ( .A(_131_), .Y(_131__bF_buf5) );
BUFX4 BUFX4_475 ( .A(_131_), .Y(_131__bF_buf4) );
BUFX4 BUFX4_476 ( .A(_131_), .Y(_131__bF_buf3) );
BUFX4 BUFX4_477 ( .A(_131_), .Y(_131__bF_buf2) );
BUFX4 BUFX4_478 ( .A(_131_), .Y(_131__bF_buf1) );
BUFX4 BUFX4_479 ( .A(_131_), .Y(_131__bF_buf0) );
BUFX4 BUFX4_480 ( .A(_4606_), .Y(_4606__bF_buf4) );
BUFX4 BUFX4_481 ( .A(_4606_), .Y(_4606__bF_buf3) );
BUFX4 BUFX4_482 ( .A(_4606_), .Y(_4606__bF_buf2) );
BUFX4 BUFX4_483 ( .A(_4606_), .Y(_4606__bF_buf1) );
BUFX4 BUFX4_484 ( .A(_4606_), .Y(_4606__bF_buf0) );
BUFX4 BUFX4_485 ( .A(_4224_), .Y(_4224__bF_buf4) );
BUFX4 BUFX4_486 ( .A(_4224_), .Y(_4224__bF_buf3) );
BUFX4 BUFX4_487 ( .A(_4224_), .Y(_4224__bF_buf2) );
BUFX4 BUFX4_488 ( .A(_4224_), .Y(_4224__bF_buf1) );
BUFX4 BUFX4_489 ( .A(_4224_), .Y(_4224__bF_buf0) );
BUFX4 BUFX4_490 ( .A(_4262_), .Y(_4262__bF_buf4) );
BUFX4 BUFX4_491 ( .A(_4262_), .Y(_4262__bF_buf3) );
BUFX4 BUFX4_492 ( .A(_4262_), .Y(_4262__bF_buf2) );
BUFX4 BUFX4_493 ( .A(_4262_), .Y(_4262__bF_buf1) );
BUFX4 BUFX4_494 ( .A(_4262_), .Y(_4262__bF_buf0) );
BUFX4 BUFX4_495 ( .A(_701_), .Y(_701__bF_buf4) );
BUFX4 BUFX4_496 ( .A(_701_), .Y(_701__bF_buf3) );
BUFX4 BUFX4_497 ( .A(_701_), .Y(_701__bF_buf2) );
BUFX4 BUFX4_498 ( .A(_701_), .Y(_701__bF_buf1) );
BUFX4 BUFX4_499 ( .A(_701_), .Y(_701__bF_buf0) );
BUFX4 BUFX4_500 ( .A(micro_hash_ucr_pipe60), .Y(micro_hash_ucr_pipe60_bF_buf4) );
BUFX4 BUFX4_501 ( .A(micro_hash_ucr_pipe60), .Y(micro_hash_ucr_pipe60_bF_buf3) );
BUFX4 BUFX4_502 ( .A(micro_hash_ucr_pipe60), .Y(micro_hash_ucr_pipe60_bF_buf2) );
BUFX4 BUFX4_503 ( .A(micro_hash_ucr_pipe60), .Y(micro_hash_ucr_pipe60_bF_buf1) );
BUFX4 BUFX4_504 ( .A(micro_hash_ucr_pipe60), .Y(micro_hash_ucr_pipe60_bF_buf0) );
BUFX4 BUFX4_505 ( .A(micro_hash_ucr_pipe61), .Y(micro_hash_ucr_pipe61_bF_buf3) );
BUFX4 BUFX4_506 ( .A(micro_hash_ucr_pipe61), .Y(micro_hash_ucr_pipe61_bF_buf2) );
BUFX4 BUFX4_507 ( .A(micro_hash_ucr_pipe61), .Y(micro_hash_ucr_pipe61_bF_buf1) );
BUFX4 BUFX4_508 ( .A(micro_hash_ucr_pipe61), .Y(micro_hash_ucr_pipe61_bF_buf0) );
BUFX4 BUFX4_509 ( .A(micro_hash_ucr_pipe62), .Y(micro_hash_ucr_pipe62_bF_buf3) );
BUFX4 BUFX4_510 ( .A(micro_hash_ucr_pipe62), .Y(micro_hash_ucr_pipe62_bF_buf2) );
BUFX4 BUFX4_511 ( .A(micro_hash_ucr_pipe62), .Y(micro_hash_ucr_pipe62_bF_buf1) );
BUFX4 BUFX4_512 ( .A(micro_hash_ucr_pipe62), .Y(micro_hash_ucr_pipe62_bF_buf0) );
BUFX4 BUFX4_513 ( .A(micro_hash_ucr_pipe63), .Y(micro_hash_ucr_pipe63_bF_buf3) );
BUFX4 BUFX4_514 ( .A(micro_hash_ucr_pipe63), .Y(micro_hash_ucr_pipe63_bF_buf2) );
BUFX4 BUFX4_515 ( .A(micro_hash_ucr_pipe63), .Y(micro_hash_ucr_pipe63_bF_buf1) );
BUFX4 BUFX4_516 ( .A(micro_hash_ucr_pipe63), .Y(micro_hash_ucr_pipe63_bF_buf0) );
BUFX4 BUFX4_517 ( .A(micro_hash_ucr_pipe64), .Y(micro_hash_ucr_pipe64_bF_buf4) );
BUFX4 BUFX4_518 ( .A(micro_hash_ucr_pipe64), .Y(micro_hash_ucr_pipe64_bF_buf3) );
BUFX4 BUFX4_519 ( .A(micro_hash_ucr_pipe64), .Y(micro_hash_ucr_pipe64_bF_buf2) );
BUFX4 BUFX4_520 ( .A(micro_hash_ucr_pipe64), .Y(micro_hash_ucr_pipe64_bF_buf1) );
BUFX4 BUFX4_521 ( .A(micro_hash_ucr_pipe64), .Y(micro_hash_ucr_pipe64_bF_buf0) );
BUFX4 BUFX4_522 ( .A(micro_hash_ucr_pipe65), .Y(micro_hash_ucr_pipe65_bF_buf4) );
BUFX4 BUFX4_523 ( .A(micro_hash_ucr_pipe65), .Y(micro_hash_ucr_pipe65_bF_buf3) );
BUFX4 BUFX4_524 ( .A(micro_hash_ucr_pipe65), .Y(micro_hash_ucr_pipe65_bF_buf2) );
BUFX4 BUFX4_525 ( .A(micro_hash_ucr_pipe65), .Y(micro_hash_ucr_pipe65_bF_buf1) );
BUFX4 BUFX4_526 ( .A(micro_hash_ucr_pipe65), .Y(micro_hash_ucr_pipe65_bF_buf0) );
BUFX4 BUFX4_527 ( .A(micro_hash_ucr_pipe66), .Y(micro_hash_ucr_pipe66_bF_buf4) );
BUFX4 BUFX4_528 ( .A(micro_hash_ucr_pipe66), .Y(micro_hash_ucr_pipe66_bF_buf3) );
BUFX4 BUFX4_529 ( .A(micro_hash_ucr_pipe66), .Y(micro_hash_ucr_pipe66_bF_buf2) );
BUFX4 BUFX4_530 ( .A(micro_hash_ucr_pipe66), .Y(micro_hash_ucr_pipe66_bF_buf1) );
BUFX4 BUFX4_531 ( .A(micro_hash_ucr_pipe66), .Y(micro_hash_ucr_pipe66_bF_buf0) );
BUFX4 BUFX4_532 ( .A(_1120_), .Y(_1120__bF_buf4) );
BUFX4 BUFX4_533 ( .A(_1120_), .Y(_1120__bF_buf3) );
BUFX4 BUFX4_534 ( .A(_1120_), .Y(_1120__bF_buf2) );
BUFX4 BUFX4_535 ( .A(_1120_), .Y(_1120__bF_buf1) );
BUFX4 BUFX4_536 ( .A(_1120_), .Y(_1120__bF_buf0) );
BUFX4 BUFX4_537 ( .A(micro_hash_ucr_b_7_), .Y(micro_hash_ucr_b_7_bF_buf3_) );
BUFX4 BUFX4_538 ( .A(micro_hash_ucr_b_7_), .Y(micro_hash_ucr_b_7_bF_buf2_) );
BUFX4 BUFX4_539 ( .A(micro_hash_ucr_b_7_), .Y(micro_hash_ucr_b_7_bF_buf1_) );
BUFX4 BUFX4_540 ( .A(micro_hash_ucr_b_7_), .Y(micro_hash_ucr_b_7_bF_buf0_) );
BUFX4 BUFX4_541 ( .A(_389_), .Y(_389__bF_buf3) );
BUFX4 BUFX4_542 ( .A(_389_), .Y(_389__bF_buf2) );
BUFX4 BUFX4_543 ( .A(_389_), .Y(_389__bF_buf1) );
BUFX4 BUFX4_544 ( .A(_389_), .Y(_389__bF_buf0) );
BUFX4 BUFX4_545 ( .A(_4218_), .Y(_4218__bF_buf3) );
BUFX4 BUFX4_546 ( .A(_4218_), .Y(_4218__bF_buf2) );
BUFX4 BUFX4_547 ( .A(_4218_), .Y(_4218__bF_buf1) );
BUFX4 BUFX4_548 ( .A(_4218_), .Y(_4218__bF_buf0) );
BUFX4 BUFX4_549 ( .A(micro_hash_ucr_pipe30), .Y(micro_hash_ucr_pipe30_bF_buf3) );
BUFX4 BUFX4_550 ( .A(micro_hash_ucr_pipe30), .Y(micro_hash_ucr_pipe30_bF_buf2) );
BUFX4 BUFX4_551 ( .A(micro_hash_ucr_pipe30), .Y(micro_hash_ucr_pipe30_bF_buf1) );
BUFX4 BUFX4_552 ( .A(micro_hash_ucr_pipe30), .Y(micro_hash_ucr_pipe30_bF_buf0) );
BUFX4 BUFX4_553 ( .A(micro_hash_ucr_pipe31), .Y(micro_hash_ucr_pipe31_bF_buf3) );
BUFX4 BUFX4_554 ( .A(micro_hash_ucr_pipe31), .Y(micro_hash_ucr_pipe31_bF_buf2) );
BUFX4 BUFX4_555 ( .A(micro_hash_ucr_pipe31), .Y(micro_hash_ucr_pipe31_bF_buf1) );
BUFX4 BUFX4_556 ( .A(micro_hash_ucr_pipe31), .Y(micro_hash_ucr_pipe31_bF_buf0) );
BUFX4 BUFX4_557 ( .A(micro_hash_ucr_pipe32), .Y(micro_hash_ucr_pipe32_bF_buf4) );
BUFX4 BUFX4_558 ( .A(micro_hash_ucr_pipe32), .Y(micro_hash_ucr_pipe32_bF_buf3) );
BUFX4 BUFX4_559 ( .A(micro_hash_ucr_pipe32), .Y(micro_hash_ucr_pipe32_bF_buf2) );
BUFX4 BUFX4_560 ( .A(micro_hash_ucr_pipe32), .Y(micro_hash_ucr_pipe32_bF_buf1) );
BUFX4 BUFX4_561 ( .A(micro_hash_ucr_pipe32), .Y(micro_hash_ucr_pipe32_bF_buf0) );
BUFX4 BUFX4_562 ( .A(micro_hash_ucr_pipe33), .Y(micro_hash_ucr_pipe33_bF_buf3) );
BUFX4 BUFX4_563 ( .A(micro_hash_ucr_pipe33), .Y(micro_hash_ucr_pipe33_bF_buf2) );
BUFX4 BUFX4_564 ( .A(micro_hash_ucr_pipe33), .Y(micro_hash_ucr_pipe33_bF_buf1) );
BUFX4 BUFX4_565 ( .A(micro_hash_ucr_pipe33), .Y(micro_hash_ucr_pipe33_bF_buf0) );
BUFX4 BUFX4_566 ( .A(micro_hash_ucr_pipe34), .Y(micro_hash_ucr_pipe34_bF_buf3) );
BUFX4 BUFX4_567 ( .A(micro_hash_ucr_pipe34), .Y(micro_hash_ucr_pipe34_bF_buf2) );
BUFX4 BUFX4_568 ( .A(micro_hash_ucr_pipe34), .Y(micro_hash_ucr_pipe34_bF_buf1) );
BUFX4 BUFX4_569 ( .A(micro_hash_ucr_pipe34), .Y(micro_hash_ucr_pipe34_bF_buf0) );
BUFX4 BUFX4_570 ( .A(micro_hash_ucr_pipe36), .Y(micro_hash_ucr_pipe36_bF_buf3) );
BUFX4 BUFX4_571 ( .A(micro_hash_ucr_pipe36), .Y(micro_hash_ucr_pipe36_bF_buf2) );
BUFX4 BUFX4_572 ( .A(micro_hash_ucr_pipe36), .Y(micro_hash_ucr_pipe36_bF_buf1) );
BUFX4 BUFX4_573 ( .A(micro_hash_ucr_pipe36), .Y(micro_hash_ucr_pipe36_bF_buf0) );
BUFX4 BUFX4_574 ( .A(micro_hash_ucr_pipe37), .Y(micro_hash_ucr_pipe37_bF_buf3) );
BUFX4 BUFX4_575 ( .A(micro_hash_ucr_pipe37), .Y(micro_hash_ucr_pipe37_bF_buf2) );
BUFX4 BUFX4_576 ( .A(micro_hash_ucr_pipe37), .Y(micro_hash_ucr_pipe37_bF_buf1) );
BUFX4 BUFX4_577 ( .A(micro_hash_ucr_pipe37), .Y(micro_hash_ucr_pipe37_bF_buf0) );
BUFX4 BUFX4_578 ( .A(micro_hash_ucr_pipe38), .Y(micro_hash_ucr_pipe38_bF_buf3) );
BUFX4 BUFX4_579 ( .A(micro_hash_ucr_pipe38), .Y(micro_hash_ucr_pipe38_bF_buf2) );
BUFX4 BUFX4_580 ( .A(micro_hash_ucr_pipe38), .Y(micro_hash_ucr_pipe38_bF_buf1) );
BUFX4 BUFX4_581 ( .A(micro_hash_ucr_pipe38), .Y(micro_hash_ucr_pipe38_bF_buf0) );
BUFX4 BUFX4_582 ( .A(micro_hash_ucr_c_1_), .Y(micro_hash_ucr_c_1_bF_buf3_) );
BUFX4 BUFX4_583 ( .A(micro_hash_ucr_c_1_), .Y(micro_hash_ucr_c_1_bF_buf2_) );
BUFX4 BUFX4_584 ( .A(micro_hash_ucr_c_1_), .Y(micro_hash_ucr_c_1_bF_buf1_) );
BUFX4 BUFX4_585 ( .A(micro_hash_ucr_c_1_), .Y(micro_hash_ucr_c_1_bF_buf0_) );
BUFX4 BUFX4_586 ( .A(_827_), .Y(_827__bF_buf5) );
BUFX4 BUFX4_587 ( .A(_827_), .Y(_827__bF_buf4) );
BUFX4 BUFX4_588 ( .A(_827_), .Y(_827__bF_buf3) );
BUFX4 BUFX4_589 ( .A(_827_), .Y(_827__bF_buf2) );
BUFX4 BUFX4_590 ( .A(_827_), .Y(_827__bF_buf1) );
BUFX4 BUFX4_591 ( .A(_827_), .Y(_827__bF_buf0) );
BUFX4 BUFX4_592 ( .A(micro_hash_ucr_a_7_), .Y(micro_hash_ucr_a_7_bF_buf3_) );
BUFX4 BUFX4_593 ( .A(micro_hash_ucr_a_7_), .Y(micro_hash_ucr_a_7_bF_buf2_) );
BUFX4 BUFX4_594 ( .A(micro_hash_ucr_a_7_), .Y(micro_hash_ucr_a_7_bF_buf1_) );
BUFX4 BUFX4_595 ( .A(micro_hash_ucr_a_7_), .Y(micro_hash_ucr_a_7_bF_buf0_) );
BUFX4 BUFX4_596 ( .A(_292_), .Y(_292__bF_buf12) );
BUFX4 BUFX4_597 ( .A(_292_), .Y(_292__bF_buf11) );
BUFX4 BUFX4_598 ( .A(_292_), .Y(_292__bF_buf10) );
BUFX4 BUFX4_599 ( .A(_292_), .Y(_292__bF_buf9) );
BUFX4 BUFX4_600 ( .A(_292_), .Y(_292__bF_buf8) );
BUFX4 BUFX4_601 ( .A(_292_), .Y(_292__bF_buf7) );
BUFX4 BUFX4_602 ( .A(_292_), .Y(_292__bF_buf6) );
BUFX4 BUFX4_603 ( .A(_292_), .Y(_292__bF_buf5) );
BUFX4 BUFX4_604 ( .A(_292_), .Y(_292__bF_buf4) );
BUFX4 BUFX4_605 ( .A(_292_), .Y(_292__bF_buf3) );
BUFX4 BUFX4_606 ( .A(_292_), .Y(_292__bF_buf2) );
BUFX4 BUFX4_607 ( .A(_292_), .Y(_292__bF_buf1) );
BUFX4 BUFX4_608 ( .A(_292_), .Y(_292__bF_buf0) );
BUFX4 BUFX4_609 ( .A(_4215_), .Y(_4215__bF_buf4) );
BUFX4 BUFX4_610 ( .A(_4215_), .Y(_4215__bF_buf3) );
BUFX4 BUFX4_611 ( .A(_4215_), .Y(_4215__bF_buf2) );
BUFX4 BUFX4_612 ( .A(_4215_), .Y(_4215__bF_buf1) );
BUFX4 BUFX4_613 ( .A(_4215_), .Y(_4215__bF_buf0) );
BUFX4 BUFX4_614 ( .A(micro_hash_ucr_b_1_), .Y(micro_hash_ucr_b_1_bF_buf3_) );
BUFX4 BUFX4_615 ( .A(micro_hash_ucr_b_1_), .Y(micro_hash_ucr_b_1_bF_buf2_) );
BUFX4 BUFX4_616 ( .A(micro_hash_ucr_b_1_), .Y(micro_hash_ucr_b_1_bF_buf1_) );
BUFX4 BUFX4_617 ( .A(micro_hash_ucr_b_1_), .Y(micro_hash_ucr_b_1_bF_buf0_) );
BUFX4 BUFX4_618 ( .A(_824_), .Y(_824__bF_buf3) );
BUFX4 BUFX4_619 ( .A(_824_), .Y(_824__bF_buf2) );
BUFX4 BUFX4_620 ( .A(_824_), .Y(_824__bF_buf1) );
BUFX4 BUFX4_621 ( .A(_824_), .Y(_824__bF_buf0) );
BUFX4 BUFX4_622 ( .A(micro_hash_ucr_a_4_), .Y(micro_hash_ucr_a_4_bF_buf3_) );
BUFX4 BUFX4_623 ( .A(micro_hash_ucr_a_4_), .Y(micro_hash_ucr_a_4_bF_buf2_) );
BUFX4 BUFX4_624 ( .A(micro_hash_ucr_a_4_), .Y(micro_hash_ucr_a_4_bF_buf1_) );
BUFX4 BUFX4_625 ( .A(micro_hash_ucr_a_4_), .Y(micro_hash_ucr_a_4_bF_buf0_) );
BUFX4 BUFX4_626 ( .A(_624_), .Y(_624__bF_buf3) );
BUFX4 BUFX4_627 ( .A(_624_), .Y(_624__bF_buf2) );
BUFX4 BUFX4_628 ( .A(_624_), .Y(_624__bF_buf1) );
BUFX4 BUFX4_629 ( .A(_624_), .Y(_624__bF_buf0) );
BUFX4 BUFX4_630 ( .A(_1942_), .Y(_1942__bF_buf5) );
BUFX4 BUFX4_631 ( .A(_1942_), .Y(_1942__bF_buf4) );
BUFX4 BUFX4_632 ( .A(_1942_), .Y(_1942__bF_buf3) );
BUFX4 BUFX4_633 ( .A(_1942_), .Y(_1942__bF_buf2) );
BUFX4 BUFX4_634 ( .A(_1942_), .Y(_1942__bF_buf1) );
BUFX4 BUFX4_635 ( .A(_1942_), .Y(_1942__bF_buf0) );
BUFX4 BUFX4_636 ( .A(_242_), .Y(_242__bF_buf3) );
BUFX4 BUFX4_637 ( .A(_242_), .Y(_242__bF_buf2) );
BUFX4 BUFX4_638 ( .A(_242_), .Y(_242__bF_buf1) );
BUFX4 BUFX4_639 ( .A(_242_), .Y(_242__bF_buf0) );
BUFX4 BUFX4_640 ( .A(_4241_), .Y(_4241__bF_buf3) );
BUFX4 BUFX4_641 ( .A(_4241_), .Y(_4241__bF_buf2) );
BUFX4 BUFX4_642 ( .A(_4241_), .Y(_4241__bF_buf1) );
BUFX4 BUFX4_643 ( .A(_4241_), .Y(_4241__bF_buf0) );
BUFX4 BUFX4_644 ( .A(_1078_), .Y(_1078__bF_buf3) );
BUFX4 BUFX4_645 ( .A(_1078_), .Y(_1078__bF_buf2) );
BUFX4 BUFX4_646 ( .A(_1078_), .Y(_1078__bF_buf1) );
BUFX4 BUFX4_647 ( .A(_1078_), .Y(_1078__bF_buf0) );
BUFX4 BUFX4_648 ( .A(_4238_), .Y(_4238__bF_buf3) );
BUFX4 BUFX4_649 ( .A(_4238_), .Y(_4238__bF_buf2) );
BUFX4 BUFX4_650 ( .A(_4238_), .Y(_4238__bF_buf1) );
BUFX4 BUFX4_651 ( .A(_4238_), .Y(_4238__bF_buf0) );
BUFX4 BUFX4_652 ( .A(_597_), .Y(_597__bF_buf4) );
BUFX4 BUFX4_653 ( .A(_597_), .Y(_597__bF_buf3) );
BUFX4 BUFX4_654 ( .A(_597_), .Y(_597__bF_buf2) );
BUFX4 BUFX4_655 ( .A(_597_), .Y(_597__bF_buf1) );
BUFX4 BUFX4_656 ( .A(_597_), .Y(_597__bF_buf0) );
BUFX4 BUFX4_657 ( .A(reset), .Y(reset_bF_buf5) );
BUFX4 BUFX4_658 ( .A(reset), .Y(reset_bF_buf4) );
BUFX4 BUFX4_659 ( .A(reset), .Y(reset_bF_buf3) );
BUFX4 BUFX4_660 ( .A(reset), .Y(reset_bF_buf2) );
BUFX4 BUFX4_661 ( .A(reset), .Y(reset_bF_buf1) );
BUFX4 BUFX4_662 ( .A(reset), .Y(reset_bF_buf0) );
BUFX4 BUFX4_663 ( .A(_230_), .Y(_230__bF_buf3) );
BUFX4 BUFX4_664 ( .A(_230_), .Y(_230__bF_buf2) );
BUFX4 BUFX4_665 ( .A(_230_), .Y(_230__bF_buf1) );
BUFX4 BUFX4_666 ( .A(_230_), .Y(_230__bF_buf0) );
BUFX4 BUFX4_667 ( .A(_591_), .Y(_591__bF_buf3) );
BUFX4 BUFX4_668 ( .A(_591_), .Y(_591__bF_buf2) );
BUFX4 BUFX4_669 ( .A(_591_), .Y(_591__bF_buf1) );
BUFX4 BUFX4_670 ( .A(_591_), .Y(_591__bF_buf0) );
BUFX4 BUFX4_671 ( .A(_1125_), .Y(_1125__bF_buf4) );
BUFX4 BUFX4_672 ( .A(_1125_), .Y(_1125__bF_buf3) );
BUFX4 BUFX4_673 ( .A(_1125_), .Y(_1125__bF_buf2) );
BUFX4 BUFX4_674 ( .A(_1125_), .Y(_1125__bF_buf1) );
BUFX4 BUFX4_675 ( .A(_1125_), .Y(_1125__bF_buf0) );
OAI21X1 OAI21X1_1 ( .A(_4409_), .B(_4283__bF_buf32), .C(_4408_), .Y(_4281__62_) );
NAND2X1 NAND2X1_1 ( .A(next_b_data_in_prev_63_), .B(_4283__bF_buf16), .Y(_4410_) );
MUX2X1 MUX2X1_1 ( .A(data_in[63]), .B(next_b_data_in_prev_63_), .S(_0__bF_buf0), .Y(_4411_) );
OAI21X1 OAI21X1_2 ( .A(_4411_), .B(_4283__bF_buf16), .C(_4410_), .Y(_4281__63_) );
NAND2X1 NAND2X1_2 ( .A(next_b_data_in_prev_64_), .B(_4283__bF_buf36), .Y(_4412_) );
MUX2X1 MUX2X1_2 ( .A(data_in[64]), .B(next_b_data_in_prev_64_), .S(_0__bF_buf1), .Y(_4413_) );
OAI21X1 OAI21X1_3 ( .A(_4413_), .B(_4283__bF_buf36), .C(_4412_), .Y(_4281__64_) );
NAND2X1 NAND2X1_3 ( .A(next_b_data_in_prev_65_), .B(_4283__bF_buf38), .Y(_4414_) );
MUX2X1 MUX2X1_3 ( .A(data_in[65]), .B(next_b_data_in_prev_65_), .S(_0__bF_buf6), .Y(_4415_) );
OAI21X1 OAI21X1_4 ( .A(_4415_), .B(_4283__bF_buf38), .C(_4414_), .Y(_4281__65_) );
NAND2X1 NAND2X1_4 ( .A(next_b_data_in_prev_66_), .B(_4283__bF_buf6), .Y(_4416_) );
MUX2X1 MUX2X1_4 ( .A(data_in[66]), .B(next_b_data_in_prev_66_), .S(_0__bF_buf3), .Y(_4417_) );
OAI21X1 OAI21X1_5 ( .A(_4417_), .B(_4283__bF_buf6), .C(_4416_), .Y(_4281__66_) );
NAND2X1 NAND2X1_5 ( .A(next_b_data_in_prev_67_), .B(_4283__bF_buf0), .Y(_4418_) );
MUX2X1 MUX2X1_5 ( .A(data_in[67]), .B(next_b_data_in_prev_67_), .S(_0__bF_buf1), .Y(_4419_) );
OAI21X1 OAI21X1_6 ( .A(_4419_), .B(_4283__bF_buf0), .C(_4418_), .Y(_4281__67_) );
NAND2X1 NAND2X1_6 ( .A(next_b_data_in_prev_68_), .B(_4283__bF_buf30), .Y(_4420_) );
MUX2X1 MUX2X1_6 ( .A(data_in[68]), .B(next_b_data_in_prev_68_), .S(_0__bF_buf0), .Y(_4421_) );
OAI21X1 OAI21X1_7 ( .A(_4421_), .B(_4283__bF_buf30), .C(_4420_), .Y(_4281__68_) );
NAND2X1 NAND2X1_7 ( .A(next_b_data_in_prev_69_), .B(_4283__bF_buf35), .Y(_4422_) );
MUX2X1 MUX2X1_7 ( .A(data_in[69]), .B(next_b_data_in_prev_69_), .S(_0__bF_buf5), .Y(_4423_) );
OAI21X1 OAI21X1_8 ( .A(_4423_), .B(_4283__bF_buf35), .C(_4422_), .Y(_4281__69_) );
NAND2X1 NAND2X1_8 ( .A(next_b_data_in_prev_70_), .B(_4283__bF_buf11), .Y(_4424_) );
MUX2X1 MUX2X1_8 ( .A(data_in[70]), .B(next_b_data_in_prev_70_), .S(_0__bF_buf7), .Y(_4425_) );
OAI21X1 OAI21X1_9 ( .A(_4425_), .B(_4283__bF_buf11), .C(_4424_), .Y(_4281__70_) );
NAND2X1 NAND2X1_9 ( .A(next_b_data_in_prev_71_), .B(_4283__bF_buf33), .Y(_4426_) );
MUX2X1 MUX2X1_9 ( .A(data_in[71]), .B(next_b_data_in_prev_71_), .S(_0__bF_buf4), .Y(_4427_) );
OAI21X1 OAI21X1_10 ( .A(_4427_), .B(_4283__bF_buf33), .C(_4426_), .Y(_4281__71_) );
NAND2X1 NAND2X1_10 ( .A(next_b_data_in_prev_72_), .B(_4283__bF_buf15), .Y(_4428_) );
MUX2X1 MUX2X1_10 ( .A(data_in[72]), .B(next_b_data_in_prev_72_), .S(_0__bF_buf8), .Y(_4429_) );
OAI21X1 OAI21X1_11 ( .A(_4429_), .B(_4283__bF_buf15), .C(_4428_), .Y(_4281__72_) );
NAND2X1 NAND2X1_11 ( .A(next_b_data_in_prev_73_), .B(_4283__bF_buf26), .Y(_4430_) );
MUX2X1 MUX2X1_11 ( .A(data_in[73]), .B(next_b_data_in_prev_73_), .S(_0__bF_buf7), .Y(_4431_) );
OAI21X1 OAI21X1_12 ( .A(_4431_), .B(_4283__bF_buf26), .C(_4430_), .Y(_4281__73_) );
NAND2X1 NAND2X1_12 ( .A(next_b_data_in_prev_74_), .B(_4283__bF_buf41), .Y(_4432_) );
MUX2X1 MUX2X1_12 ( .A(data_in[74]), .B(next_b_data_in_prev_74_), .S(_0__bF_buf8), .Y(_4433_) );
OAI21X1 OAI21X1_13 ( .A(_4433_), .B(_4283__bF_buf41), .C(_4432_), .Y(_4281__74_) );
NAND2X1 NAND2X1_13 ( .A(next_b_data_in_prev_75_), .B(_4283__bF_buf36), .Y(_4434_) );
MUX2X1 MUX2X1_13 ( .A(data_in[75]), .B(next_b_data_in_prev_75_), .S(_0__bF_buf1), .Y(_4435_) );
OAI21X1 OAI21X1_14 ( .A(_4435_), .B(_4283__bF_buf36), .C(_4434_), .Y(_4281__75_) );
NAND2X1 NAND2X1_14 ( .A(next_b_data_in_prev_76_), .B(_4283__bF_buf10), .Y(_4436_) );
MUX2X1 MUX2X1_14 ( .A(data_in[76]), .B(next_b_data_in_prev_76_), .S(_0__bF_buf5), .Y(_4437_) );
OAI21X1 OAI21X1_15 ( .A(_4437_), .B(_4283__bF_buf10), .C(_4436_), .Y(_4281__76_) );
NAND2X1 NAND2X1_15 ( .A(next_b_data_in_prev_77_), .B(_4283__bF_buf25), .Y(_4438_) );
MUX2X1 MUX2X1_15 ( .A(data_in[77]), .B(next_b_data_in_prev_77_), .S(_0__bF_buf1), .Y(_4439_) );
OAI21X1 OAI21X1_16 ( .A(_4439_), .B(_4283__bF_buf25), .C(_4438_), .Y(_4281__77_) );
NAND2X1 NAND2X1_16 ( .A(next_b_data_in_prev_78_), .B(_4283__bF_buf31), .Y(_4440_) );
MUX2X1 MUX2X1_16 ( .A(data_in[78]), .B(next_b_data_in_prev_78_), .S(_0__bF_buf2), .Y(_4441_) );
OAI21X1 OAI21X1_17 ( .A(_4441_), .B(_4283__bF_buf31), .C(_4440_), .Y(_4281__78_) );
NAND2X1 NAND2X1_17 ( .A(next_b_data_in_prev_79_), .B(_4283__bF_buf35), .Y(_4442_) );
MUX2X1 MUX2X1_17 ( .A(data_in[79]), .B(next_b_data_in_prev_79_), .S(_0__bF_buf5), .Y(_4443_) );
OAI21X1 OAI21X1_18 ( .A(_4443_), .B(_4283__bF_buf35), .C(_4442_), .Y(_4281__79_) );
NAND2X1 NAND2X1_18 ( .A(next_b_data_in_prev_80_), .B(_4283__bF_buf20), .Y(_4444_) );
MUX2X1 MUX2X1_18 ( .A(data_in[80]), .B(next_b_data_in_prev_80_), .S(_0__bF_buf3), .Y(_4445_) );
OAI21X1 OAI21X1_19 ( .A(_4445_), .B(_4283__bF_buf20), .C(_4444_), .Y(_4281__80_) );
NAND2X1 NAND2X1_19 ( .A(next_b_data_in_prev_81_), .B(_4283__bF_buf21), .Y(_4446_) );
MUX2X1 MUX2X1_19 ( .A(data_in[81]), .B(next_b_data_in_prev_81_), .S(_0__bF_buf0), .Y(_4447_) );
OAI21X1 OAI21X1_20 ( .A(_4447_), .B(_4283__bF_buf21), .C(_4446_), .Y(_4281__81_) );
NAND2X1 NAND2X1_20 ( .A(next_b_data_in_prev_82_), .B(_4283__bF_buf31), .Y(_4448_) );
MUX2X1 MUX2X1_20 ( .A(data_in[82]), .B(next_b_data_in_prev_82_), .S(_0__bF_buf2), .Y(_4449_) );
OAI21X1 OAI21X1_21 ( .A(_4449_), .B(_4283__bF_buf5), .C(_4448_), .Y(_4281__82_) );
NAND2X1 NAND2X1_21 ( .A(next_b_data_in_prev_83_), .B(_4283__bF_buf40), .Y(_4450_) );
MUX2X1 MUX2X1_21 ( .A(data_in[83]), .B(next_b_data_in_prev_83_), .S(_0__bF_buf1), .Y(_4451_) );
OAI21X1 OAI21X1_22 ( .A(_4451_), .B(_4283__bF_buf40), .C(_4450_), .Y(_4281__83_) );
NAND2X1 NAND2X1_22 ( .A(next_b_data_in_prev_84_), .B(_4283__bF_buf31), .Y(_4452_) );
MUX2X1 MUX2X1_22 ( .A(data_in[84]), .B(next_b_data_in_prev_84_), .S(_0__bF_buf2), .Y(_4453_) );
OAI21X1 OAI21X1_23 ( .A(_4453_), .B(_4283__bF_buf31), .C(_4452_), .Y(_4281__84_) );
NAND2X1 NAND2X1_23 ( .A(next_b_data_in_prev_85_), .B(_4283__bF_buf38), .Y(_4454_) );
MUX2X1 MUX2X1_23 ( .A(data_in[85]), .B(next_b_data_in_prev_85_), .S(_0__bF_buf6), .Y(_4455_) );
OAI21X1 OAI21X1_24 ( .A(_4455_), .B(_4283__bF_buf3), .C(_4454_), .Y(_4281__85_) );
NAND2X1 NAND2X1_24 ( .A(next_b_data_in_prev_86_), .B(_4283__bF_buf19), .Y(_4456_) );
MUX2X1 MUX2X1_24 ( .A(data_in[86]), .B(next_b_data_in_prev_86_), .S(_0__bF_buf0), .Y(_4457_) );
OAI21X1 OAI21X1_25 ( .A(_4457_), .B(_4283__bF_buf19), .C(_4456_), .Y(_4281__86_) );
NAND2X1 NAND2X1_25 ( .A(next_b_data_in_prev_87_), .B(_4283__bF_buf10), .Y(_4458_) );
MUX2X1 MUX2X1_25 ( .A(data_in[87]), .B(next_b_data_in_prev_87_), .S(_0__bF_buf5), .Y(_4459_) );
OAI21X1 OAI21X1_26 ( .A(_4459_), .B(_4283__bF_buf10), .C(_4458_), .Y(_4281__87_) );
NAND2X1 NAND2X1_26 ( .A(next_b_data_in_prev_88_), .B(_4283__bF_buf12), .Y(_4460_) );
MUX2X1 MUX2X1_26 ( .A(data_in[88]), .B(next_b_data_in_prev_88_), .S(_0__bF_buf8), .Y(_4461_) );
OAI21X1 OAI21X1_27 ( .A(_4461_), .B(_4283__bF_buf12), .C(_4460_), .Y(_4281__88_) );
NAND2X1 NAND2X1_27 ( .A(next_b_data_in_prev_89_), .B(_4283__bF_buf14), .Y(_4462_) );
MUX2X1 MUX2X1_27 ( .A(data_in[89]), .B(next_b_data_in_prev_89_), .S(_0__bF_buf2), .Y(_4463_) );
OAI21X1 OAI21X1_28 ( .A(_4463_), .B(_4283__bF_buf14), .C(_4462_), .Y(_4281__89_) );
NAND2X1 NAND2X1_28 ( .A(next_b_data_in_prev_90_), .B(_4283__bF_buf37), .Y(_4464_) );
MUX2X1 MUX2X1_28 ( .A(data_in[90]), .B(next_b_data_in_prev_90_), .S(_0__bF_buf8), .Y(_4465_) );
OAI21X1 OAI21X1_29 ( .A(_4465_), .B(_4283__bF_buf37), .C(_4464_), .Y(_4281__90_) );
NAND2X1 NAND2X1_29 ( .A(next_b_data_in_prev_91_), .B(_4283__bF_buf7), .Y(_4466_) );
MUX2X1 MUX2X1_29 ( .A(data_in[91]), .B(next_b_data_in_prev_91_), .S(_0__bF_buf1), .Y(_4467_) );
OAI21X1 OAI21X1_30 ( .A(_4467_), .B(_4283__bF_buf7), .C(_4466_), .Y(_4281__91_) );
NAND2X1 NAND2X1_30 ( .A(next_b_data_in_prev_92_), .B(_4283__bF_buf11), .Y(_4468_) );
MUX2X1 MUX2X1_30 ( .A(data_in[92]), .B(next_b_data_in_prev_92_), .S(_0__bF_buf7), .Y(_4469_) );
OAI21X1 OAI21X1_31 ( .A(_4469_), .B(_4283__bF_buf11), .C(_4468_), .Y(_4281__92_) );
NAND2X1 NAND2X1_31 ( .A(next_b_data_in_prev_93_), .B(_4283__bF_buf14), .Y(_4470_) );
MUX2X1 MUX2X1_31 ( .A(data_in[93]), .B(next_b_data_in_prev_93_), .S(_0__bF_buf2), .Y(_4471_) );
OAI21X1 OAI21X1_32 ( .A(_4471_), .B(_4283__bF_buf14), .C(_4470_), .Y(_4281__93_) );
NAND2X1 NAND2X1_32 ( .A(next_b_data_in_prev_94_), .B(_4283__bF_buf3), .Y(_4472_) );
MUX2X1 MUX2X1_32 ( .A(data_in[94]), .B(next_b_data_in_prev_94_), .S(_0__bF_buf6), .Y(_4473_) );
OAI21X1 OAI21X1_33 ( .A(_4473_), .B(_4283__bF_buf3), .C(_4472_), .Y(_4281__94_) );
NAND2X1 NAND2X1_33 ( .A(next_b_data_in_prev_95_), .B(_4283__bF_buf11), .Y(_4474_) );
MUX2X1 MUX2X1_33 ( .A(data_in[95]), .B(next_b_data_in_prev_95_), .S(_0__bF_buf0), .Y(_4475_) );
OAI21X1 OAI21X1_34 ( .A(_4475_), .B(_4283__bF_buf19), .C(_4474_), .Y(_4281__95_) );
NOR2X1 NOR2X1_1 ( .A(_4283__bF_buf28), .B(_4285_), .Y(_4282__0_) );
NOR2X1 NOR2X1_2 ( .A(_4283__bF_buf16), .B(_4287_), .Y(_4282__1_) );
NOR2X1 NOR2X1_3 ( .A(_4283__bF_buf34), .B(_4289_), .Y(_4282__2_) );
NOR2X1 NOR2X1_4 ( .A(_4283__bF_buf5), .B(_4291_), .Y(_4282__3_) );
NOR2X1 NOR2X1_5 ( .A(_4283__bF_buf20), .B(_4293_), .Y(_4282__4_) );
NOR2X1 NOR2X1_6 ( .A(_4283__bF_buf33), .B(_4295_), .Y(_4282__5_) );
NOR2X1 NOR2X1_7 ( .A(_4283__bF_buf33), .B(_4297_), .Y(_4282__6_) );
NOR2X1 NOR2X1_8 ( .A(_4283__bF_buf17), .B(_4299_), .Y(_4282__7_) );
NOR2X1 NOR2X1_9 ( .A(_4283__bF_buf21), .B(_4301_), .Y(_4282__8_) );
NOR2X1 NOR2X1_10 ( .A(_4283__bF_buf41), .B(_4303_), .Y(_4282__9_) );
NOR2X1 NOR2X1_11 ( .A(_4283__bF_buf18), .B(_4305_), .Y(_4282__10_) );
NOR2X1 NOR2X1_12 ( .A(_4283__bF_buf34), .B(_4307_), .Y(_4282__11_) );
NOR2X1 NOR2X1_13 ( .A(_4283__bF_buf24), .B(_4309_), .Y(_4282__12_) );
NOR2X1 NOR2X1_14 ( .A(_4283__bF_buf3), .B(_4311_), .Y(_4282__13_) );
NOR2X1 NOR2X1_15 ( .A(_4283__bF_buf32), .B(_4313_), .Y(_4282__14_) );
NOR2X1 NOR2X1_16 ( .A(_4283__bF_buf27), .B(_4315_), .Y(_4282__15_) );
NOR2X1 NOR2X1_17 ( .A(_4283__bF_buf40), .B(_4317_), .Y(_4282__16_) );
NOR2X1 NOR2X1_18 ( .A(_4283__bF_buf42), .B(_4319_), .Y(_4282__17_) );
NOR2X1 NOR2X1_19 ( .A(_4283__bF_buf30), .B(_4321_), .Y(_4282__18_) );
NOR2X1 NOR2X1_20 ( .A(_4283__bF_buf20), .B(_4323_), .Y(_4282__19_) );
NOR2X1 NOR2X1_21 ( .A(_4283__bF_buf30), .B(_4325_), .Y(_4282__20_) );
NOR2X1 NOR2X1_22 ( .A(_4283__bF_buf29), .B(_4327_), .Y(_4282__21_) );
NOR2X1 NOR2X1_23 ( .A(_4283__bF_buf39), .B(_4329_), .Y(_4282__22_) );
NOR2X1 NOR2X1_24 ( .A(_4283__bF_buf35), .B(_4331_), .Y(_4282__23_) );
NOR2X1 NOR2X1_25 ( .A(_4283__bF_buf38), .B(_4333_), .Y(_4282__24_) );
NOR2X1 NOR2X1_26 ( .A(_4283__bF_buf18), .B(_4335_), .Y(_4282__25_) );
NOR2X1 NOR2X1_27 ( .A(_4283__bF_buf37), .B(_4337_), .Y(_4282__26_) );
NOR2X1 NOR2X1_28 ( .A(_4283__bF_buf41), .B(_4339_), .Y(_4282__27_) );
NOR2X1 NOR2X1_29 ( .A(_4283__bF_buf23), .B(_4341_), .Y(_4282__28_) );
NOR2X1 NOR2X1_30 ( .A(_4283__bF_buf1), .B(_4343_), .Y(_4282__29_) );
NOR2X1 NOR2X1_31 ( .A(_4283__bF_buf24), .B(_4345_), .Y(_4282__30_) );
NOR2X1 NOR2X1_32 ( .A(_4283__bF_buf2), .B(_4347_), .Y(_4282__31_) );
NOR2X1 NOR2X1_33 ( .A(_4283__bF_buf25), .B(_4349_), .Y(_4282__32_) );
NOR2X1 NOR2X1_34 ( .A(_4283__bF_buf15), .B(_4351_), .Y(_4282__33_) );
NOR2X1 NOR2X1_35 ( .A(_4283__bF_buf40), .B(_4353_), .Y(_4282__34_) );
NOR2X1 NOR2X1_36 ( .A(_4283__bF_buf5), .B(_4355_), .Y(_4282__35_) );
NOR2X1 NOR2X1_37 ( .A(_4283__bF_buf17), .B(_4357_), .Y(_4282__36_) );
NOR2X1 NOR2X1_38 ( .A(_4283__bF_buf4), .B(_4359_), .Y(_4282__37_) );
NOR2X1 NOR2X1_39 ( .A(_4283__bF_buf27), .B(_4361_), .Y(_4282__38_) );
NOR2X1 NOR2X1_40 ( .A(_4283__bF_buf2), .B(_4363_), .Y(_4282__39_) );
NOR2X1 NOR2X1_41 ( .A(_4283__bF_buf14), .B(_4365_), .Y(_4282__40_) );
NOR2X1 NOR2X1_42 ( .A(_4283__bF_buf0), .B(_4367_), .Y(_4282__41_) );
NOR2X1 NOR2X1_43 ( .A(_4283__bF_buf41), .B(_4369_), .Y(_4282__42_) );
NOR2X1 NOR2X1_44 ( .A(_4283__bF_buf13), .B(_4371_), .Y(_4282__43_) );
NOR2X1 NOR2X1_45 ( .A(_4283__bF_buf4), .B(_4373_), .Y(_4282__44_) );
NOR2X1 NOR2X1_46 ( .A(_4283__bF_buf4), .B(_4375_), .Y(_4282__45_) );
NOR2X1 NOR2X1_47 ( .A(_4283__bF_buf1), .B(_4377_), .Y(_4282__46_) );
NOR2X1 NOR2X1_48 ( .A(_4283__bF_buf35), .B(_4379_), .Y(_4282__47_) );
NOR2X1 NOR2X1_49 ( .A(_4283__bF_buf4), .B(_4381_), .Y(_4282__48_) );
NOR2X1 NOR2X1_50 ( .A(_4283__bF_buf20), .B(_4383_), .Y(_4282__49_) );
NOR2X1 NOR2X1_51 ( .A(_4283__bF_buf42), .B(_4385_), .Y(_4282__50_) );
NOR2X1 NOR2X1_52 ( .A(_4283__bF_buf17), .B(_4387_), .Y(_4282__51_) );
NOR2X1 NOR2X1_53 ( .A(_4283__bF_buf24), .B(_4389_), .Y(_4282__52_) );
NOR2X1 NOR2X1_54 ( .A(_4283__bF_buf28), .B(_4391_), .Y(_4282__53_) );
NOR2X1 NOR2X1_55 ( .A(_4283__bF_buf38), .B(_4393_), .Y(_4282__54_) );
NOR2X1 NOR2X1_56 ( .A(_4283__bF_buf17), .B(_4395_), .Y(_4282__55_) );
NOR2X1 NOR2X1_57 ( .A(_4283__bF_buf38), .B(_4397_), .Y(_4282__56_) );
NOR2X1 NOR2X1_58 ( .A(_4283__bF_buf37), .B(_4399_), .Y(_4282__57_) );
NOR2X1 NOR2X1_59 ( .A(_4283__bF_buf12), .B(_4401_), .Y(_4282__58_) );
NOR2X1 NOR2X1_60 ( .A(_4283__bF_buf5), .B(_4403_), .Y(_4282__59_) );
NOR2X1 NOR2X1_61 ( .A(_4283__bF_buf18), .B(_4405_), .Y(_4282__60_) );
NOR2X1 NOR2X1_62 ( .A(_4283__bF_buf0), .B(_4407_), .Y(_4282__61_) );
NOR2X1 NOR2X1_63 ( .A(_4283__bF_buf35), .B(_4409_), .Y(_4282__62_) );
NOR2X1 NOR2X1_64 ( .A(_4283__bF_buf3), .B(_4411_), .Y(_4282__63_) );
NOR2X1 NOR2X1_65 ( .A(_4283__bF_buf14), .B(_4413_), .Y(_4282__64_) );
NOR2X1 NOR2X1_66 ( .A(_4283__bF_buf38), .B(_4415_), .Y(_4282__65_) );
NOR2X1 NOR2X1_67 ( .A(_4283__bF_buf15), .B(_4417_), .Y(_4282__66_) );
NOR2X1 NOR2X1_68 ( .A(_4283__bF_buf0), .B(_4419_), .Y(_4282__67_) );
NOR2X1 NOR2X1_69 ( .A(_4283__bF_buf16), .B(_4421_), .Y(_4282__68_) );
NOR2X1 NOR2X1_70 ( .A(_4283__bF_buf1), .B(_4423_), .Y(_4282__69_) );
NOR2X1 NOR2X1_71 ( .A(_4283__bF_buf26), .B(_4425_), .Y(_4282__70_) );
NOR2X1 NOR2X1_72 ( .A(_4283__bF_buf17), .B(_4427_), .Y(_4282__71_) );
NOR2X1 NOR2X1_73 ( .A(_4283__bF_buf15), .B(_4429_), .Y(_4282__72_) );
NOR2X1 NOR2X1_74 ( .A(_4283__bF_buf16), .B(_4431_), .Y(_4282__73_) );
NOR2X1 NOR2X1_75 ( .A(_4283__bF_buf42), .B(_4433_), .Y(_4282__74_) );
NOR2X1 NOR2X1_76 ( .A(_4283__bF_buf40), .B(_4435_), .Y(_4282__75_) );
NOR2X1 NOR2X1_77 ( .A(_4283__bF_buf10), .B(_4437_), .Y(_4282__76_) );
NOR2X1 NOR2X1_78 ( .A(_4283__bF_buf7), .B(_4439_), .Y(_4282__77_) );
NOR2X1 NOR2X1_79 ( .A(_4283__bF_buf4), .B(_4441_), .Y(_4282__78_) );
NOR2X1 NOR2X1_80 ( .A(_4283__bF_buf2), .B(_4443_), .Y(_4282__79_) );
NOR2X1 NOR2X1_81 ( .A(_4283__bF_buf28), .B(_4445_), .Y(_4282__80_) );
NOR2X1 NOR2X1_82 ( .A(_4283__bF_buf24), .B(_4447_), .Y(_4282__81_) );
NOR2X1 NOR2X1_83 ( .A(_4283__bF_buf18), .B(_4449_), .Y(_4282__82_) );
NOR2X1 NOR2X1_84 ( .A(_4283__bF_buf40), .B(_4451_), .Y(_4282__83_) );
NOR2X1 NOR2X1_85 ( .A(_4283__bF_buf4), .B(_4453_), .Y(_4282__84_) );
NOR2X1 NOR2X1_86 ( .A(_4283__bF_buf3), .B(_4455_), .Y(_4282__85_) );
NOR2X1 NOR2X1_87 ( .A(_4283__bF_buf24), .B(_4457_), .Y(_4282__86_) );
NOR2X1 NOR2X1_88 ( .A(_4283__bF_buf10), .B(_4459_), .Y(_4282__87_) );
NOR2X1 NOR2X1_89 ( .A(_4283__bF_buf12), .B(_4461_), .Y(_4282__88_) );
NOR2X1 NOR2X1_90 ( .A(_4283__bF_buf14), .B(_4463_), .Y(_4282__89_) );
NOR2X1 NOR2X1_91 ( .A(_4283__bF_buf37), .B(_4465_), .Y(_4282__90_) );
NOR2X1 NOR2X1_92 ( .A(_4283__bF_buf7), .B(_4467_), .Y(_4282__91_) );
NOR2X1 NOR2X1_93 ( .A(_4283__bF_buf16), .B(_4469_), .Y(_4282__92_) );
NOR2X1 NOR2X1_94 ( .A(_4283__bF_buf18), .B(_4471_), .Y(_4282__93_) );
NOR2X1 NOR2X1_95 ( .A(_4283__bF_buf1), .B(_4473_), .Y(_4282__94_) );
NOR2X1 NOR2X1_96 ( .A(_4283__bF_buf16), .B(_4475_), .Y(_4282__95_) );
DFFPOSX1 DFFPOSX1_1 ( .CLK(clk_bF_buf39), .D(_4282__0_), .Q(concatenador_bloque_0_) );
DFFPOSX1 DFFPOSX1_2 ( .CLK(clk_bF_buf45), .D(_4282__1_), .Q(concatenador_bloque_1_) );
DFFPOSX1 DFFPOSX1_3 ( .CLK(clk_bF_buf58), .D(_4282__2_), .Q(concatenador_bloque_2_) );
DFFPOSX1 DFFPOSX1_4 ( .CLK(clk_bF_buf38), .D(_4282__3_), .Q(concatenador_bloque_3_) );
DFFPOSX1 DFFPOSX1_5 ( .CLK(clk_bF_buf34), .D(_4282__4_), .Q(concatenador_bloque_4_) );
DFFPOSX1 DFFPOSX1_6 ( .CLK(clk_bF_buf36), .D(_4282__5_), .Q(concatenador_bloque_5_) );
DFFPOSX1 DFFPOSX1_7 ( .CLK(clk_bF_buf57), .D(_4282__6_), .Q(concatenador_bloque_6_) );
DFFPOSX1 DFFPOSX1_8 ( .CLK(clk_bF_buf78), .D(_4282__7_), .Q(concatenador_bloque_7_) );
DFFPOSX1 DFFPOSX1_9 ( .CLK(clk_bF_buf20), .D(_4282__8_), .Q(concatenador_bloque_8_) );
DFFPOSX1 DFFPOSX1_10 ( .CLK(clk_bF_buf39), .D(_4282__9_), .Q(concatenador_bloque_9_) );
DFFPOSX1 DFFPOSX1_11 ( .CLK(clk_bF_buf13), .D(_4282__10_), .Q(concatenador_bloque_10_) );
DFFPOSX1 DFFPOSX1_12 ( .CLK(clk_bF_buf38), .D(_4282__11_), .Q(concatenador_bloque_11_) );
DFFPOSX1 DFFPOSX1_13 ( .CLK(clk_bF_buf32), .D(_4282__12_), .Q(concatenador_bloque_12_) );
DFFPOSX1 DFFPOSX1_14 ( .CLK(clk_bF_buf32), .D(_4282__13_), .Q(concatenador_bloque_13_) );
DFFPOSX1 DFFPOSX1_15 ( .CLK(clk_bF_buf66), .D(_4282__14_), .Q(concatenador_bloque_14_) );
DFFPOSX1 DFFPOSX1_16 ( .CLK(clk_bF_buf65), .D(_4282__15_), .Q(concatenador_bloque_15_) );
DFFPOSX1 DFFPOSX1_17 ( .CLK(clk_bF_buf45), .D(_4282__16_), .Q(concatenador_bloque_16_) );
DFFPOSX1 DFFPOSX1_18 ( .CLK(clk_bF_buf74), .D(_4282__17_), .Q(concatenador_bloque_17_) );
DFFPOSX1 DFFPOSX1_19 ( .CLK(clk_bF_buf4), .D(_4282__18_), .Q(concatenador_bloque_18_) );
DFFPOSX1 DFFPOSX1_20 ( .CLK(clk_bF_buf38), .D(_4282__19_), .Q(concatenador_bloque_19_) );
DFFPOSX1 DFFPOSX1_21 ( .CLK(clk_bF_buf4), .D(_4282__20_), .Q(concatenador_bloque_20_) );
DFFPOSX1 DFFPOSX1_22 ( .CLK(clk_bF_buf26), .D(_4282__21_), .Q(concatenador_bloque_21_) );
DFFPOSX1 DFFPOSX1_23 ( .CLK(clk_bF_buf72), .D(_4282__22_), .Q(concatenador_bloque_22_) );
DFFPOSX1 DFFPOSX1_24 ( .CLK(clk_bF_buf37), .D(_4282__23_), .Q(concatenador_bloque_23_) );
DFFPOSX1 DFFPOSX1_25 ( .CLK(clk_bF_buf52), .D(_4282__24_), .Q(concatenador_bloque_24_) );
DFFPOSX1 DFFPOSX1_26 ( .CLK(clk_bF_buf13), .D(_4282__25_), .Q(concatenador_bloque_25_) );
DFFPOSX1 DFFPOSX1_27 ( .CLK(clk_bF_buf53), .D(_4282__26_), .Q(concatenador_bloque_26_) );
DFFPOSX1 DFFPOSX1_28 ( .CLK(clk_bF_buf53), .D(_4282__27_), .Q(concatenador_bloque_27_) );
DFFPOSX1 DFFPOSX1_29 ( .CLK(clk_bF_buf4), .D(_4282__28_), .Q(concatenador_bloque_28_) );
DFFPOSX1 DFFPOSX1_30 ( .CLK(clk_bF_buf77), .D(_4282__29_), .Q(concatenador_bloque_29_) );
DFFPOSX1 DFFPOSX1_31 ( .CLK(clk_bF_buf57), .D(_4282__30_), .Q(concatenador_bloque_30_) );
DFFPOSX1 DFFPOSX1_32 ( .CLK(clk_bF_buf66), .D(_4282__31_), .Q(concatenador_bloque_31_) );
DFFPOSX1 DFFPOSX1_33 ( .CLK(clk_bF_buf40), .D(_4282__32_), .Q(concatenador_bloque_32_) );
DFFPOSX1 DFFPOSX1_34 ( .CLK(clk_bF_buf58), .D(_4282__33_), .Q(concatenador_bloque_33_) );
DFFPOSX1 DFFPOSX1_35 ( .CLK(clk_bF_buf73), .D(_4282__34_), .Q(concatenador_bloque_34_) );
DFFPOSX1 DFFPOSX1_36 ( .CLK(clk_bF_buf13), .D(_4282__35_), .Q(concatenador_bloque_35_) );
DFFPOSX1 DFFPOSX1_37 ( .CLK(clk_bF_buf4), .D(_4282__36_), .Q(concatenador_bloque_36_) );
DFFPOSX1 DFFPOSX1_38 ( .CLK(clk_bF_buf20), .D(_4282__37_), .Q(concatenador_bloque_37_) );
DFFPOSX1 DFFPOSX1_39 ( .CLK(clk_bF_buf47), .D(_4282__38_), .Q(concatenador_bloque_38_) );
DFFPOSX1 DFFPOSX1_40 ( .CLK(clk_bF_buf37), .D(_4282__39_), .Q(concatenador_bloque_39_) );
DFFPOSX1 DFFPOSX1_41 ( .CLK(clk_bF_buf20), .D(_4282__40_), .Q(concatenador_bloque_40_) );
DFFPOSX1 DFFPOSX1_42 ( .CLK(clk_bF_buf35), .D(_4282__41_), .Q(concatenador_bloque_41_) );
DFFPOSX1 DFFPOSX1_43 ( .CLK(clk_bF_buf53), .D(_4282__42_), .Q(concatenador_bloque_42_) );
DFFPOSX1 DFFPOSX1_44 ( .CLK(clk_bF_buf61), .D(_4282__43_), .Q(concatenador_bloque_43_) );
DFFPOSX1 DFFPOSX1_45 ( .CLK(clk_bF_buf20), .D(_4282__44_), .Q(concatenador_bloque_44_) );
DFFPOSX1 DFFPOSX1_46 ( .CLK(clk_bF_buf52), .D(_4282__45_), .Q(concatenador_bloque_45_) );
DFFPOSX1 DFFPOSX1_47 ( .CLK(clk_bF_buf77), .D(_4282__46_), .Q(concatenador_bloque_46_) );
DFFPOSX1 DFFPOSX1_48 ( .CLK(clk_bF_buf26), .D(_4282__47_), .Q(concatenador_bloque_47_) );
DFFPOSX1 DFFPOSX1_49 ( .CLK(clk_bF_buf20), .D(_4282__48_), .Q(concatenador_bloque_48_) );
DFFPOSX1 DFFPOSX1_50 ( .CLK(clk_bF_buf30), .D(_4282__49_), .Q(concatenador_bloque_49_) );
DFFPOSX1 DFFPOSX1_51 ( .CLK(clk_bF_buf74), .D(_4282__50_), .Q(concatenador_bloque_50_) );
DFFPOSX1 DFFPOSX1_52 ( .CLK(clk_bF_buf38), .D(_4282__51_), .Q(concatenador_bloque_51_) );
DFFPOSX1 DFFPOSX1_53 ( .CLK(clk_bF_buf32), .D(_4282__52_), .Q(concatenador_bloque_52_) );
DFFPOSX1 DFFPOSX1_54 ( .CLK(clk_bF_buf39), .D(_4282__53_), .Q(concatenador_bloque_53_) );
DFFPOSX1 DFFPOSX1_55 ( .CLK(clk_bF_buf32), .D(_4282__54_), .Q(concatenador_bloque_54_) );
DFFPOSX1 DFFPOSX1_56 ( .CLK(clk_bF_buf4), .D(_4282__55_), .Q(concatenador_bloque_55_) );
DFFPOSX1 DFFPOSX1_57 ( .CLK(clk_bF_buf42), .D(_4282__56_), .Q(concatenador_bloque_56_) );
DFFPOSX1 DFFPOSX1_58 ( .CLK(clk_bF_buf27), .D(_4282__57_), .Q(concatenador_bloque_57_) );
DFFPOSX1 DFFPOSX1_59 ( .CLK(clk_bF_buf74), .D(_4282__58_), .Q(concatenador_bloque_58_) );
DFFPOSX1 DFFPOSX1_60 ( .CLK(clk_bF_buf13), .D(_4282__59_), .Q(concatenador_bloque_59_) );
DFFPOSX1 DFFPOSX1_61 ( .CLK(clk_bF_buf38), .D(_4282__60_), .Q(concatenador_bloque_60_) );
DFFPOSX1 DFFPOSX1_62 ( .CLK(clk_bF_buf42), .D(_4282__61_), .Q(concatenador_bloque_61_) );
DFFPOSX1 DFFPOSX1_63 ( .CLK(clk_bF_buf6), .D(_4282__62_), .Q(concatenador_bloque_62_) );
DFFPOSX1 DFFPOSX1_64 ( .CLK(clk_bF_buf66), .D(_4282__63_), .Q(concatenador_bloque_63_) );
DFFPOSX1 DFFPOSX1_65 ( .CLK(clk_bF_buf30), .D(_4282__64_), .Q(concatenador_bloque_64_) );
DFFPOSX1 DFFPOSX1_66 ( .CLK(clk_bF_buf32), .D(_4282__65_), .Q(concatenador_bloque_65_) );
DFFPOSX1 DFFPOSX1_67 ( .CLK(clk_bF_buf30), .D(_4282__66_), .Q(concatenador_bloque_66_) );
DFFPOSX1 DFFPOSX1_68 ( .CLK(clk_bF_buf36), .D(_4282__67_), .Q(concatenador_bloque_67_) );
DFFPOSX1 DFFPOSX1_69 ( .CLK(clk_bF_buf36), .D(_4282__68_), .Q(concatenador_bloque_68_) );
DFFPOSX1 DFFPOSX1_70 ( .CLK(clk_bF_buf6), .D(_4282__69_), .Q(concatenador_bloque_69_) );
DFFPOSX1 DFFPOSX1_71 ( .CLK(clk_bF_buf4), .D(_4282__70_), .Q(concatenador_bloque_70_) );
DFFPOSX1 DFFPOSX1_72 ( .CLK(clk_bF_buf78), .D(_4282__71_), .Q(concatenador_bloque_71_) );
DFFPOSX1 DFFPOSX1_73 ( .CLK(clk_bF_buf74), .D(_4282__72_), .Q(concatenador_bloque_72_) );
DFFPOSX1 DFFPOSX1_74 ( .CLK(clk_bF_buf78), .D(_4282__73_), .Q(concatenador_bloque_73_) );
DFFPOSX1 DFFPOSX1_75 ( .CLK(clk_bF_buf70), .D(_4282__74_), .Q(concatenador_bloque_74_) );
DFFPOSX1 DFFPOSX1_76 ( .CLK(clk_bF_buf73), .D(_4282__75_), .Q(concatenador_bloque_75_) );
DFFPOSX1 DFFPOSX1_77 ( .CLK(clk_bF_buf67), .D(_4282__76_), .Q(concatenador_bloque_76_) );
DFFPOSX1 DFFPOSX1_78 ( .CLK(clk_bF_buf6), .D(_4282__77_), .Q(concatenador_bloque_77_) );
DFFPOSX1 DFFPOSX1_79 ( .CLK(clk_bF_buf52), .D(_4282__78_), .Q(concatenador_bloque_78_) );
DFFPOSX1 DFFPOSX1_80 ( .CLK(clk_bF_buf37), .D(_4282__79_), .Q(concatenador_bloque_79_) );
DFFPOSX1 DFFPOSX1_81 ( .CLK(clk_bF_buf79), .D(_4282__80_), .Q(concatenador_bloque_80_) );
DFFPOSX1 DFFPOSX1_82 ( .CLK(clk_bF_buf32), .D(_4282__81_), .Q(concatenador_bloque_81_) );
DFFPOSX1 DFFPOSX1_83 ( .CLK(clk_bF_buf38), .D(_4282__82_), .Q(concatenador_bloque_82_) );
DFFPOSX1 DFFPOSX1_84 ( .CLK(clk_bF_buf35), .D(_4282__83_), .Q(concatenador_bloque_83_) );
DFFPOSX1 DFFPOSX1_85 ( .CLK(clk_bF_buf34), .D(_4282__84_), .Q(concatenador_bloque_84_) );
DFFPOSX1 DFFPOSX1_86 ( .CLK(clk_bF_buf32), .D(_4282__85_), .Q(concatenador_bloque_85_) );
DFFPOSX1 DFFPOSX1_87 ( .CLK(clk_bF_buf36), .D(_4282__86_), .Q(concatenador_bloque_86_) );
DFFPOSX1 DFFPOSX1_88 ( .CLK(clk_bF_buf65), .D(_4282__87_), .Q(concatenador_bloque_87_) );
DFFPOSX1 DFFPOSX1_89 ( .CLK(clk_bF_buf74), .D(_4282__88_), .Q(concatenador_bloque_88_) );
DFFPOSX1 DFFPOSX1_90 ( .CLK(clk_bF_buf73), .D(_4282__89_), .Q(concatenador_bloque_89_) );
DFFPOSX1 DFFPOSX1_91 ( .CLK(clk_bF_buf74), .D(_4282__90_), .Q(concatenador_bloque_90_) );
DFFPOSX1 DFFPOSX1_92 ( .CLK(clk_bF_buf36), .D(_4282__91_), .Q(concatenador_bloque_91_) );
DFFPOSX1 DFFPOSX1_93 ( .CLK(clk_bF_buf4), .D(_4282__92_), .Q(concatenador_bloque_92_) );
DFFPOSX1 DFFPOSX1_94 ( .CLK(clk_bF_buf13), .D(_4282__93_), .Q(concatenador_bloque_93_) );
DFFPOSX1 DFFPOSX1_95 ( .CLK(clk_bF_buf67), .D(_4282__94_), .Q(concatenador_bloque_94_) );
DFFPOSX1 DFFPOSX1_96 ( .CLK(clk_bF_buf57), .D(_4282__95_), .Q(concatenador_bloque_95_) );
DFFPOSX1 DFFPOSX1_97 ( .CLK(clk_bF_buf79), .D(_4281__0_), .Q(next_b_data_in_prev_0_) );
DFFPOSX1 DFFPOSX1_98 ( .CLK(clk_bF_buf78), .D(_4281__1_), .Q(next_b_data_in_prev_1_) );
DFFPOSX1 DFFPOSX1_99 ( .CLK(clk_bF_buf73), .D(_4281__2_), .Q(next_b_data_in_prev_2_) );
DFFPOSX1 DFFPOSX1_100 ( .CLK(clk_bF_buf40), .D(_4281__3_), .Q(next_b_data_in_prev_3_) );
DFFPOSX1 DFFPOSX1_101 ( .CLK(clk_bF_buf73), .D(_4281__4_), .Q(next_b_data_in_prev_4_) );
DFFPOSX1 DFFPOSX1_102 ( .CLK(clk_bF_buf61), .D(_4281__5_), .Q(next_b_data_in_prev_5_) );
DFFPOSX1 DFFPOSX1_103 ( .CLK(clk_bF_buf28), .D(_4281__6_), .Q(next_b_data_in_prev_6_) );
DFFPOSX1 DFFPOSX1_104 ( .CLK(clk_bF_buf28), .D(_4281__7_), .Q(next_b_data_in_prev_7_) );
DFFPOSX1 DFFPOSX1_105 ( .CLK(clk_bF_buf56), .D(_4281__8_), .Q(next_b_data_in_prev_8_) );
DFFPOSX1 DFFPOSX1_106 ( .CLK(clk_bF_buf58), .D(_4281__9_), .Q(next_b_data_in_prev_9_) );
DFFPOSX1 DFFPOSX1_107 ( .CLK(clk_bF_buf40), .D(_4281__10_), .Q(next_b_data_in_prev_10_) );
DFFPOSX1 DFFPOSX1_108 ( .CLK(clk_bF_buf38), .D(_4281__11_), .Q(next_b_data_in_prev_11_) );
DFFPOSX1 DFFPOSX1_109 ( .CLK(clk_bF_buf57), .D(_4281__12_), .Q(next_b_data_in_prev_12_) );
DFFPOSX1 DFFPOSX1_110 ( .CLK(clk_bF_buf56), .D(_4281__13_), .Q(next_b_data_in_prev_13_) );
DFFPOSX1 DFFPOSX1_111 ( .CLK(clk_bF_buf56), .D(_4281__14_), .Q(next_b_data_in_prev_14_) );
DFFPOSX1 DFFPOSX1_112 ( .CLK(clk_bF_buf10), .D(_4281__15_), .Q(next_b_data_in_prev_15_) );
DFFPOSX1 DFFPOSX1_113 ( .CLK(clk_bF_buf28), .D(_4281__16_), .Q(next_b_data_in_prev_16_) );
DFFPOSX1 DFFPOSX1_114 ( .CLK(clk_bF_buf53), .D(_4281__17_), .Q(next_b_data_in_prev_17_) );
DFFPOSX1 DFFPOSX1_115 ( .CLK(clk_bF_buf28), .D(_4281__18_), .Q(next_b_data_in_prev_18_) );
DFFPOSX1 DFFPOSX1_116 ( .CLK(clk_bF_buf38), .D(_4281__19_), .Q(next_b_data_in_prev_19_) );
DFFPOSX1 DFFPOSX1_117 ( .CLK(clk_bF_buf28), .D(_4281__20_), .Q(next_b_data_in_prev_20_) );
DFFPOSX1 DFFPOSX1_118 ( .CLK(clk_bF_buf56), .D(_4281__21_), .Q(next_b_data_in_prev_21_) );
DFFPOSX1 DFFPOSX1_119 ( .CLK(clk_bF_buf56), .D(_4281__22_), .Q(next_b_data_in_prev_22_) );
DFFPOSX1 DFFPOSX1_120 ( .CLK(clk_bF_buf26), .D(_4281__23_), .Q(next_b_data_in_prev_23_) );
DFFPOSX1 DFFPOSX1_121 ( .CLK(clk_bF_buf61), .D(_4281__24_), .Q(next_b_data_in_prev_24_) );
DFFPOSX1 DFFPOSX1_122 ( .CLK(clk_bF_buf73), .D(_4281__25_), .Q(next_b_data_in_prev_25_) );
DFFPOSX1 DFFPOSX1_123 ( .CLK(clk_bF_buf53), .D(_4281__26_), .Q(next_b_data_in_prev_26_) );
DFFPOSX1 DFFPOSX1_124 ( .CLK(clk_bF_buf30), .D(_4281__27_), .Q(next_b_data_in_prev_27_) );
DFFPOSX1 DFFPOSX1_125 ( .CLK(clk_bF_buf61), .D(_4281__28_), .Q(next_b_data_in_prev_28_) );
DFFPOSX1 DFFPOSX1_126 ( .CLK(clk_bF_buf37), .D(_4281__29_), .Q(next_b_data_in_prev_29_) );
DFFPOSX1 DFFPOSX1_127 ( .CLK(clk_bF_buf78), .D(_4281__30_), .Q(next_b_data_in_prev_30_) );
DFFPOSX1 DFFPOSX1_128 ( .CLK(clk_bF_buf26), .D(_4281__31_), .Q(next_b_data_in_prev_31_) );
DFFPOSX1 DFFPOSX1_129 ( .CLK(clk_bF_buf61), .D(_4281__32_), .Q(next_b_data_in_prev_32_) );
DFFPOSX1 DFFPOSX1_130 ( .CLK(clk_bF_buf58), .D(_4281__33_), .Q(next_b_data_in_prev_33_) );
DFFPOSX1 DFFPOSX1_131 ( .CLK(clk_bF_buf61), .D(_4281__34_), .Q(next_b_data_in_prev_34_) );
DFFPOSX1 DFFPOSX1_132 ( .CLK(clk_bF_buf45), .D(_4281__35_), .Q(next_b_data_in_prev_35_) );
DFFPOSX1 DFFPOSX1_133 ( .CLK(clk_bF_buf78), .D(_4281__36_), .Q(next_b_data_in_prev_36_) );
DFFPOSX1 DFFPOSX1_134 ( .CLK(clk_bF_buf56), .D(_4281__37_), .Q(next_b_data_in_prev_37_) );
DFFPOSX1 DFFPOSX1_135 ( .CLK(clk_bF_buf37), .D(_4281__38_), .Q(next_b_data_in_prev_38_) );
DFFPOSX1 DFFPOSX1_136 ( .CLK(clk_bF_buf37), .D(_4281__39_), .Q(next_b_data_in_prev_39_) );
DFFPOSX1 DFFPOSX1_137 ( .CLK(clk_bF_buf35), .D(_4281__40_), .Q(next_b_data_in_prev_40_) );
DFFPOSX1 DFFPOSX1_138 ( .CLK(clk_bF_buf61), .D(_4281__41_), .Q(next_b_data_in_prev_41_) );
DFFPOSX1 DFFPOSX1_139 ( .CLK(clk_bF_buf73), .D(_4281__42_), .Q(next_b_data_in_prev_42_) );
DFFPOSX1 DFFPOSX1_140 ( .CLK(clk_bF_buf28), .D(_4281__43_), .Q(next_b_data_in_prev_43_) );
DFFPOSX1 DFFPOSX1_141 ( .CLK(clk_bF_buf35), .D(_4281__44_), .Q(next_b_data_in_prev_44_) );
DFFPOSX1 DFFPOSX1_142 ( .CLK(clk_bF_buf35), .D(_4281__45_), .Q(next_b_data_in_prev_45_) );
DFFPOSX1 DFFPOSX1_143 ( .CLK(clk_bF_buf26), .D(_4281__46_), .Q(next_b_data_in_prev_46_) );
DFFPOSX1 DFFPOSX1_144 ( .CLK(clk_bF_buf26), .D(_4281__47_), .Q(next_b_data_in_prev_47_) );
DFFPOSX1 DFFPOSX1_145 ( .CLK(clk_bF_buf40), .D(_4281__48_), .Q(next_b_data_in_prev_48_) );
DFFPOSX1 DFFPOSX1_146 ( .CLK(clk_bF_buf73), .D(_4281__49_), .Q(next_b_data_in_prev_49_) );
DFFPOSX1 DFFPOSX1_147 ( .CLK(clk_bF_buf53), .D(_4281__50_), .Q(next_b_data_in_prev_50_) );
DFFPOSX1 DFFPOSX1_148 ( .CLK(clk_bF_buf78), .D(_4281__51_), .Q(next_b_data_in_prev_51_) );
DFFPOSX1 DFFPOSX1_149 ( .CLK(clk_bF_buf61), .D(_4281__52_), .Q(next_b_data_in_prev_52_) );
DFFPOSX1 DFFPOSX1_150 ( .CLK(clk_bF_buf58), .D(_4281__53_), .Q(next_b_data_in_prev_53_) );
DFFPOSX1 DFFPOSX1_151 ( .CLK(clk_bF_buf4), .D(_4281__54_), .Q(next_b_data_in_prev_54_) );
DFFPOSX1 DFFPOSX1_152 ( .CLK(clk_bF_buf61), .D(_4281__55_), .Q(next_b_data_in_prev_55_) );
DFFPOSX1 DFFPOSX1_153 ( .CLK(clk_bF_buf57), .D(_4281__56_), .Q(next_b_data_in_prev_56_) );
DFFPOSX1 DFFPOSX1_154 ( .CLK(clk_bF_buf53), .D(_4281__57_), .Q(next_b_data_in_prev_57_) );
DFFPOSX1 DFFPOSX1_155 ( .CLK(clk_bF_buf73), .D(_4281__58_), .Q(next_b_data_in_prev_58_) );
DFFPOSX1 DFFPOSX1_156 ( .CLK(clk_bF_buf73), .D(_4281__59_), .Q(next_b_data_in_prev_59_) );
DFFPOSX1 DFFPOSX1_157 ( .CLK(clk_bF_buf35), .D(_4281__60_), .Q(next_b_data_in_prev_60_) );
DFFPOSX1 DFFPOSX1_158 ( .CLK(clk_bF_buf40), .D(_4281__61_), .Q(next_b_data_in_prev_61_) );
DFFPOSX1 DFFPOSX1_159 ( .CLK(clk_bF_buf56), .D(_4281__62_), .Q(next_b_data_in_prev_62_) );
DFFPOSX1 DFFPOSX1_160 ( .CLK(clk_bF_buf78), .D(_4281__63_), .Q(next_b_data_in_prev_63_) );
DFFPOSX1 DFFPOSX1_161 ( .CLK(clk_bF_buf40), .D(_4281__64_), .Q(next_b_data_in_prev_64_) );
DFFPOSX1 DFFPOSX1_162 ( .CLK(clk_bF_buf57), .D(_4281__65_), .Q(next_b_data_in_prev_65_) );
DFFPOSX1 DFFPOSX1_163 ( .CLK(clk_bF_buf58), .D(_4281__66_), .Q(next_b_data_in_prev_66_) );
DFFPOSX1 DFFPOSX1_164 ( .CLK(clk_bF_buf4), .D(_4281__67_), .Q(next_b_data_in_prev_67_) );
DFFPOSX1 DFFPOSX1_165 ( .CLK(clk_bF_buf78), .D(_4281__68_), .Q(next_b_data_in_prev_68_) );
DFFPOSX1 DFFPOSX1_166 ( .CLK(clk_bF_buf26), .D(_4281__69_), .Q(next_b_data_in_prev_69_) );
DFFPOSX1 DFFPOSX1_167 ( .CLK(clk_bF_buf28), .D(_4281__70_), .Q(next_b_data_in_prev_70_) );
DFFPOSX1 DFFPOSX1_168 ( .CLK(clk_bF_buf61), .D(_4281__71_), .Q(next_b_data_in_prev_71_) );
DFFPOSX1 DFFPOSX1_169 ( .CLK(clk_bF_buf58), .D(_4281__72_), .Q(next_b_data_in_prev_72_) );
DFFPOSX1 DFFPOSX1_170 ( .CLK(clk_bF_buf28), .D(_4281__73_), .Q(next_b_data_in_prev_73_) );
DFFPOSX1 DFFPOSX1_171 ( .CLK(clk_bF_buf30), .D(_4281__74_), .Q(next_b_data_in_prev_74_) );
DFFPOSX1 DFFPOSX1_172 ( .CLK(clk_bF_buf40), .D(_4281__75_), .Q(next_b_data_in_prev_75_) );
DFFPOSX1 DFFPOSX1_173 ( .CLK(clk_bF_buf10), .D(_4281__76_), .Q(next_b_data_in_prev_76_) );
DFFPOSX1 DFFPOSX1_174 ( .CLK(clk_bF_buf40), .D(_4281__77_), .Q(next_b_data_in_prev_77_) );
DFFPOSX1 DFFPOSX1_175 ( .CLK(clk_bF_buf45), .D(_4281__78_), .Q(next_b_data_in_prev_78_) );
DFFPOSX1 DFFPOSX1_176 ( .CLK(clk_bF_buf26), .D(_4281__79_), .Q(next_b_data_in_prev_79_) );
DFFPOSX1 DFFPOSX1_177 ( .CLK(clk_bF_buf13), .D(_4281__80_), .Q(next_b_data_in_prev_80_) );
DFFPOSX1 DFFPOSX1_178 ( .CLK(clk_bF_buf57), .D(_4281__81_), .Q(next_b_data_in_prev_81_) );
DFFPOSX1 DFFPOSX1_179 ( .CLK(clk_bF_buf45), .D(_4281__82_), .Q(next_b_data_in_prev_82_) );
DFFPOSX1 DFFPOSX1_180 ( .CLK(clk_bF_buf35), .D(_4281__83_), .Q(next_b_data_in_prev_83_) );
DFFPOSX1 DFFPOSX1_181 ( .CLK(clk_bF_buf35), .D(_4281__84_), .Q(next_b_data_in_prev_84_) );
DFFPOSX1 DFFPOSX1_182 ( .CLK(clk_bF_buf57), .D(_4281__85_), .Q(next_b_data_in_prev_85_) );
DFFPOSX1 DFFPOSX1_183 ( .CLK(clk_bF_buf56), .D(_4281__86_), .Q(next_b_data_in_prev_86_) );
DFFPOSX1 DFFPOSX1_184 ( .CLK(clk_bF_buf37), .D(_4281__87_), .Q(next_b_data_in_prev_87_) );
DFFPOSX1 DFFPOSX1_185 ( .CLK(clk_bF_buf53), .D(_4281__88_), .Q(next_b_data_in_prev_88_) );
DFFPOSX1 DFFPOSX1_186 ( .CLK(clk_bF_buf35), .D(_4281__89_), .Q(next_b_data_in_prev_89_) );
DFFPOSX1 DFFPOSX1_187 ( .CLK(clk_bF_buf53), .D(_4281__90_), .Q(next_b_data_in_prev_90_) );
DFFPOSX1 DFFPOSX1_188 ( .CLK(clk_bF_buf40), .D(_4281__91_), .Q(next_b_data_in_prev_91_) );
DFFPOSX1 DFFPOSX1_189 ( .CLK(clk_bF_buf28), .D(_4281__92_), .Q(next_b_data_in_prev_92_) );
DFFPOSX1 DFFPOSX1_190 ( .CLK(clk_bF_buf45), .D(_4281__93_), .Q(next_b_data_in_prev_93_) );
DFFPOSX1 DFFPOSX1_191 ( .CLK(clk_bF_buf57), .D(_4281__94_), .Q(next_b_data_in_prev_94_) );
DFFPOSX1 DFFPOSX1_192 ( .CLK(clk_bF_buf78), .D(_4281__95_), .Q(next_b_data_in_prev_95_) );
AND2X2 AND2X2_1 ( .A(comparador_next), .B(concatenador_nonce_0_), .Y(_4604_) );
INVX1 INVX1_1 ( .A(reset_bF_buf1), .Y(_4605_) );
NOR2X1 NOR2X1_97 ( .A(_0__bF_buf5), .B(_4605_), .Y(_4606_) );
OAI21X1 OAI21X1_35 ( .A(comparador_next), .B(concatenador_nonce_0_), .C(_4606__bF_buf3), .Y(_4607_) );
NOR2X1 NOR2X1_98 ( .A(_4604_), .B(_4607_), .Y(_4476__0_) );
NAND2X1 NAND2X1_34 ( .A(concatenador_nonce_1_), .B(_4604_), .Y(_4608_) );
INVX2 INVX2_1 ( .A(_4608_), .Y(_4609_) );
OAI21X1 OAI21X1_36 ( .A(_4604_), .B(concatenador_nonce_1_), .C(_4606__bF_buf4), .Y(_4610_) );
NOR2X1 NOR2X1_99 ( .A(_4610_), .B(_4609_), .Y(_4476__1_) );
OAI21X1 OAI21X1_37 ( .A(_4609_), .B(concatenador_nonce_2_), .C(_4606__bF_buf4), .Y(_4611_) );
AOI21X1 AOI21X1_1 ( .A(concatenador_nonce_2_), .B(_4609_), .C(_4611_), .Y(_4476__2_) );
INVX2 INVX2_2 ( .A(concatenador_nonce_3_), .Y(_4612_) );
NAND2X1 NAND2X1_35 ( .A(concatenador_nonce_2_), .B(_4609_), .Y(_4613_) );
OAI21X1 OAI21X1_38 ( .A(_4613_), .B(_4612_), .C(_4606__bF_buf4), .Y(_4614_) );
AOI21X1 AOI21X1_2 ( .A(_4612_), .B(_4613_), .C(_4614_), .Y(_4476__3_) );
NAND3X1 NAND3X1_1 ( .A(concatenador_nonce_2_), .B(concatenador_nonce_3_), .C(concatenador_nonce_4_), .Y(_4615_) );
NOR2X1 NOR2X1_100 ( .A(_4615_), .B(_4608_), .Y(_4616_) );
NOR2X1 NOR2X1_101 ( .A(_4612_), .B(_4613_), .Y(_4617_) );
OAI21X1 OAI21X1_39 ( .A(_4617_), .B(concatenador_nonce_4_), .C(_4606__bF_buf4), .Y(_4618_) );
NOR2X1 NOR2X1_102 ( .A(_4616_), .B(_4618_), .Y(_4476__4_) );
AND2X2 AND2X2_2 ( .A(_4616_), .B(concatenador_nonce_5_), .Y(_4619_) );
OAI21X1 OAI21X1_40 ( .A(_4616_), .B(concatenador_nonce_5_), .C(_4606__bF_buf1), .Y(_4620_) );
NOR2X1 NOR2X1_103 ( .A(_4620_), .B(_4619_), .Y(_4476__5_) );
NOR2X1 NOR2X1_104 ( .A(concatenador_nonce_6_), .B(_4619_), .Y(_4621_) );
AND2X2 AND2X2_3 ( .A(concatenador_nonce_5_), .B(concatenador_nonce_6_), .Y(_4622_) );
NAND2X1 NAND2X1_36 ( .A(_4622_), .B(_4616_), .Y(_4623_) );
NAND2X1 NAND2X1_37 ( .A(_4606__bF_buf1), .B(_4623_), .Y(_4624_) );
NOR2X1 NOR2X1_105 ( .A(_4624_), .B(_4621_), .Y(_4476__6_) );
INVX2 INVX2_3 ( .A(_4623_), .Y(_4625_) );
OAI21X1 OAI21X1_41 ( .A(_4625_), .B(concatenador_nonce_7_), .C(_4606__bF_buf3), .Y(_4626_) );
AOI21X1 AOI21X1_3 ( .A(concatenador_nonce_7_), .B(_4625_), .C(_4626_), .Y(_4476__7_) );
AOI21X1 AOI21X1_4 ( .A(concatenador_nonce_7_), .B(_4625_), .C(concatenador_nonce_8_), .Y(_4627_) );
INVX1 INVX1_2 ( .A(_4615_), .Y(_4477_) );
NAND2X1 NAND2X1_38 ( .A(concatenador_nonce_5_), .B(concatenador_nonce_6_), .Y(_4478_) );
NAND2X1 NAND2X1_39 ( .A(concatenador_nonce_7_), .B(concatenador_nonce_8_), .Y(_4479_) );
NOR2X1 NOR2X1_106 ( .A(_4478_), .B(_4479_), .Y(_4480_) );
NAND2X1 NAND2X1_40 ( .A(_4477_), .B(_4480_), .Y(_4481_) );
OAI21X1 OAI21X1_42 ( .A(_4481_), .B(_4608_), .C(_4606__bF_buf3), .Y(_4482_) );
NOR2X1 NOR2X1_107 ( .A(_4482_), .B(_4627_), .Y(_4476__8_) );
NOR2X1 NOR2X1_108 ( .A(_4608_), .B(_4481_), .Y(_4483_) );
OAI21X1 OAI21X1_43 ( .A(_4483_), .B(concatenador_nonce_9_), .C(_4606__bF_buf0), .Y(_4484_) );
AOI21X1 AOI21X1_5 ( .A(concatenador_nonce_9_), .B(_4483_), .C(_4484_), .Y(_4476__9_) );
AOI21X1 AOI21X1_6 ( .A(concatenador_nonce_9_), .B(_4483_), .C(concatenador_nonce_10_), .Y(_4485_) );
AND2X2 AND2X2_4 ( .A(_4480_), .B(_4477_), .Y(_4486_) );
NAND2X1 NAND2X1_41 ( .A(_4609_), .B(_4486_), .Y(_4487_) );
NAND2X1 NAND2X1_42 ( .A(concatenador_nonce_9_), .B(concatenador_nonce_10_), .Y(_4488_) );
OAI21X1 OAI21X1_44 ( .A(_4487_), .B(_4488_), .C(_4606__bF_buf0), .Y(_4489_) );
NOR2X1 NOR2X1_109 ( .A(_4485_), .B(_4489_), .Y(_4476__10_) );
AND2X2 AND2X2_5 ( .A(concatenador_nonce_9_), .B(concatenador_nonce_10_), .Y(_4490_) );
NAND2X1 NAND2X1_43 ( .A(_4490_), .B(_4483_), .Y(_4491_) );
INVX1 INVX1_3 ( .A(_4491_), .Y(_4492_) );
OAI21X1 OAI21X1_45 ( .A(_4492_), .B(concatenador_nonce_11_), .C(_4606__bF_buf0), .Y(_4493_) );
INVX1 INVX1_4 ( .A(concatenador_nonce_11_), .Y(_4494_) );
NOR2X1 NOR2X1_110 ( .A(_4494_), .B(_4491_), .Y(_4495_) );
NOR2X1 NOR2X1_111 ( .A(_4495_), .B(_4493_), .Y(_4476__11_) );
OAI21X1 OAI21X1_46 ( .A(_4495_), .B(concatenador_nonce_12_), .C(_4606__bF_buf0), .Y(_4496_) );
AOI21X1 AOI21X1_7 ( .A(concatenador_nonce_12_), .B(_4495_), .C(_4496_), .Y(_4476__12_) );
AND2X2 AND2X2_6 ( .A(concatenador_nonce_11_), .B(concatenador_nonce_12_), .Y(_4497_) );
NAND2X1 NAND2X1_44 ( .A(_4490_), .B(_4497_), .Y(_4498_) );
NOR2X1 NOR2X1_112 ( .A(_4498_), .B(_4487_), .Y(_4499_) );
OAI21X1 OAI21X1_47 ( .A(_4499_), .B(concatenador_nonce_13_), .C(_4606__bF_buf4), .Y(_4500_) );
AOI21X1 AOI21X1_8 ( .A(concatenador_nonce_13_), .B(_4499_), .C(_4500_), .Y(_4476__13_) );
INVX4 INVX4_1 ( .A(_4606__bF_buf3), .Y(_4501_) );
INVX1 INVX1_5 ( .A(concatenador_nonce_14_), .Y(_4502_) );
NAND2X1 NAND2X1_45 ( .A(concatenador_nonce_13_), .B(_4499_), .Y(_4503_) );
NOR2X1 NOR2X1_113 ( .A(_4502_), .B(_4503_), .Y(_4504_) );
AOI21X1 AOI21X1_9 ( .A(concatenador_nonce_13_), .B(_4499_), .C(concatenador_nonce_14_), .Y(_4505_) );
NOR3X1 NOR3X1_1 ( .A(_4501_), .B(_4505_), .C(_4504_), .Y(_4476__14_) );
AND2X2 AND2X2_7 ( .A(concatenador_nonce_13_), .B(concatenador_nonce_14_), .Y(_4506_) );
NAND3X1 NAND3X1_2 ( .A(_4490_), .B(_4497_), .C(_4506_), .Y(_4507_) );
NOR2X1 NOR2X1_114 ( .A(_4507_), .B(_4487_), .Y(_4508_) );
OAI21X1 OAI21X1_48 ( .A(_4508_), .B(concatenador_nonce_15_), .C(_4606__bF_buf3), .Y(_4509_) );
AOI21X1 AOI21X1_10 ( .A(concatenador_nonce_15_), .B(_4508_), .C(_4509_), .Y(_4476__15_) );
INVX1 INVX1_6 ( .A(concatenador_nonce_15_), .Y(_4510_) );
INVX1 INVX1_7 ( .A(concatenador_nonce_16_), .Y(_4511_) );
OR2X2 OR2X2_1 ( .A(_4487_), .B(_4507_), .Y(_4512_) );
NOR3X1 NOR3X1_2 ( .A(_4510_), .B(_4511_), .C(_4512_), .Y(_4513_) );
AOI21X1 AOI21X1_11 ( .A(concatenador_nonce_15_), .B(_4508_), .C(concatenador_nonce_16_), .Y(_4514_) );
NOR3X1 NOR3X1_3 ( .A(_4501_), .B(_4514_), .C(_4513_), .Y(_4476__16_) );
INVX1 INVX1_8 ( .A(concatenador_nonce_17_), .Y(_4515_) );
NAND2X1 NAND2X1_46 ( .A(concatenador_nonce_15_), .B(concatenador_nonce_16_), .Y(_4516_) );
OR2X2 OR2X2_2 ( .A(_4507_), .B(_4516_), .Y(_4517_) );
OAI21X1 OAI21X1_49 ( .A(_4487_), .B(_4517_), .C(_4515_), .Y(_4518_) );
AND2X2 AND2X2_8 ( .A(_4518_), .B(_4606__bF_buf0), .Y(_4519_) );
NOR2X1 NOR2X1_115 ( .A(_4516_), .B(_4507_), .Y(_4520_) );
NAND3X1 NAND3X1_3 ( .A(concatenador_nonce_17_), .B(_4520_), .C(_4483_), .Y(_4521_) );
AND2X2 AND2X2_9 ( .A(_4519_), .B(_4521_), .Y(_4476__17_) );
INVX1 INVX1_9 ( .A(concatenador_nonce_18_), .Y(_4522_) );
NOR2X1 NOR2X1_116 ( .A(_4522_), .B(_4521_), .Y(_4523_) );
AND2X2 AND2X2_10 ( .A(_4521_), .B(_4522_), .Y(_4524_) );
NOR3X1 NOR3X1_4 ( .A(_4523_), .B(_4501_), .C(_4524_), .Y(_4476__18_) );
INVX2 INVX2_4 ( .A(comparador_next), .Y(_4525_) );
NAND2X1 NAND2X1_47 ( .A(concatenador_nonce_0_), .B(concatenador_nonce_1_), .Y(_4526_) );
NOR3X1 NOR3X1_5 ( .A(_4526_), .B(_4478_), .C(_4479_), .Y(_4527_) );
NAND2X1 NAND2X1_48 ( .A(concatenador_nonce_17_), .B(concatenador_nonce_18_), .Y(_4528_) );
INVX1 INVX1_10 ( .A(_4528_), .Y(_4529_) );
NAND3X1 NAND3X1_4 ( .A(_4477_), .B(_4529_), .C(_4527_), .Y(_4530_) );
NOR3X1 NOR3X1_6 ( .A(_4525_), .B(_4530_), .C(_4517_), .Y(_4531_) );
OAI21X1 OAI21X1_50 ( .A(_4531_), .B(concatenador_nonce_19_), .C(_4606__bF_buf1), .Y(_4532_) );
AND2X2 AND2X2_11 ( .A(_4531_), .B(concatenador_nonce_19_), .Y(_4533_) );
NOR2X1 NOR2X1_117 ( .A(_4532_), .B(_4533_), .Y(_4476__19_) );
NOR2X1 NOR2X1_118 ( .A(concatenador_nonce_20_), .B(_4533_), .Y(_4534_) );
NAND3X1 NAND3X1_5 ( .A(concatenador_nonce_12_), .B(concatenador_nonce_13_), .C(concatenador_nonce_14_), .Y(_4535_) );
NOR2X1 NOR2X1_119 ( .A(_4516_), .B(_4535_), .Y(_4536_) );
INVX1 INVX1_11 ( .A(_4536_), .Y(_4537_) );
NAND3X1 NAND3X1_6 ( .A(concatenador_nonce_11_), .B(concatenador_nonce_17_), .C(concatenador_nonce_18_), .Y(_4538_) );
INVX1 INVX1_12 ( .A(_4538_), .Y(_4539_) );
NOR2X1 NOR2X1_120 ( .A(_4526_), .B(_4488_), .Y(_4540_) );
NAND2X1 NAND2X1_49 ( .A(_4539_), .B(_4540_), .Y(_4541_) );
NOR3X1 NOR3X1_7 ( .A(_4481_), .B(_4541_), .C(_4537_), .Y(_4542_) );
NAND2X1 NAND2X1_50 ( .A(concatenador_nonce_19_), .B(concatenador_nonce_20_), .Y(_4543_) );
INVX1 INVX1_13 ( .A(_4543_), .Y(_4544_) );
NAND3X1 NAND3X1_7 ( .A(comparador_next), .B(_4544_), .C(_4542_), .Y(_4545_) );
NAND2X1 NAND2X1_51 ( .A(_4606__bF_buf2), .B(_4545_), .Y(_4546_) );
NOR2X1 NOR2X1_121 ( .A(_4546_), .B(_4534_), .Y(_4476__20_) );
AND2X2 AND2X2_12 ( .A(_4540_), .B(_4539_), .Y(_4547_) );
NAND3X1 NAND3X1_8 ( .A(_4536_), .B(_4486_), .C(_4547_), .Y(_4548_) );
NOR3X1 NOR3X1_8 ( .A(_4525_), .B(_4543_), .C(_4548_), .Y(_4549_) );
OAI21X1 OAI21X1_51 ( .A(_4549_), .B(concatenador_nonce_21_), .C(_4606__bF_buf2), .Y(_4550_) );
AOI21X1 AOI21X1_12 ( .A(concatenador_nonce_21_), .B(_4549_), .C(_4550_), .Y(_4476__21_) );
INVX1 INVX1_14 ( .A(concatenador_nonce_21_), .Y(_4551_) );
INVX1 INVX1_15 ( .A(concatenador_nonce_22_), .Y(_4552_) );
NOR3X1 NOR3X1_9 ( .A(_4551_), .B(_4552_), .C(_4545_), .Y(_4553_) );
AOI21X1 AOI21X1_13 ( .A(concatenador_nonce_21_), .B(_4549_), .C(concatenador_nonce_22_), .Y(_4554_) );
NOR3X1 NOR3X1_10 ( .A(_4553_), .B(_4501_), .C(_4554_), .Y(_4476__22_) );
AND2X2 AND2X2_13 ( .A(concatenador_nonce_0_), .B(concatenador_nonce_1_), .Y(_4555_) );
AND2X2 AND2X2_14 ( .A(concatenador_nonce_7_), .B(concatenador_nonce_8_), .Y(_4556_) );
NAND3X1 NAND3X1_9 ( .A(_4555_), .B(_4622_), .C(_4556_), .Y(_4557_) );
NOR3X1 NOR3X1_11 ( .A(_4615_), .B(_4528_), .C(_4557_), .Y(_4558_) );
NAND3X1 NAND3X1_10 ( .A(comparador_next), .B(_4520_), .C(_4558_), .Y(_4559_) );
NAND2X1 NAND2X1_52 ( .A(concatenador_nonce_21_), .B(concatenador_nonce_22_), .Y(_4560_) );
OR2X2 OR2X2_3 ( .A(_4543_), .B(_4560_), .Y(_4561_) );
NOR2X1 NOR2X1_122 ( .A(_4561_), .B(_4559_), .Y(_4562_) );
OAI21X1 OAI21X1_52 ( .A(_4562_), .B(concatenador_nonce_23_), .C(_4606__bF_buf2), .Y(_4563_) );
AOI21X1 AOI21X1_14 ( .A(concatenador_nonce_23_), .B(_4553_), .C(_4563_), .Y(_4476__23_) );
NAND2X1 NAND2X1_53 ( .A(concatenador_nonce_23_), .B(concatenador_nonce_24_), .Y(_4564_) );
OR2X2 OR2X2_4 ( .A(_4561_), .B(_4564_), .Y(_4565_) );
NOR2X1 NOR2X1_123 ( .A(_4565_), .B(_4559_), .Y(_4566_) );
AOI21X1 AOI21X1_15 ( .A(concatenador_nonce_23_), .B(_4562_), .C(concatenador_nonce_24_), .Y(_4567_) );
NOR3X1 NOR3X1_12 ( .A(_4501_), .B(_4566_), .C(_4567_), .Y(_4476__24_) );
INVX1 INVX1_16 ( .A(concatenador_nonce_25_), .Y(_4568_) );
NOR3X1 NOR3X1_13 ( .A(_4568_), .B(_4565_), .C(_4559_), .Y(_4569_) );
OAI21X1 OAI21X1_53 ( .A(_4566_), .B(concatenador_nonce_25_), .C(_4606__bF_buf1), .Y(_4570_) );
NOR2X1 NOR2X1_124 ( .A(_4569_), .B(_4570_), .Y(_4476__25_) );
INVX1 INVX1_17 ( .A(_4565_), .Y(_4571_) );
NAND2X1 NAND2X1_54 ( .A(_4571_), .B(_4531_), .Y(_4572_) );
OAI21X1 OAI21X1_54 ( .A(_4572_), .B(_4568_), .C(concatenador_nonce_26_), .Y(_4573_) );
INVX1 INVX1_18 ( .A(concatenador_nonce_26_), .Y(_4574_) );
NAND2X1 NAND2X1_55 ( .A(_4574_), .B(_4569_), .Y(_4575_) );
AOI21X1 AOI21X1_16 ( .A(_4575_), .B(_4573_), .C(_4501_), .Y(_4476__26_) );
INVX2 INVX2_5 ( .A(concatenador_nonce_27_), .Y(_4576_) );
NAND2X1 NAND2X1_56 ( .A(concatenador_nonce_25_), .B(concatenador_nonce_26_), .Y(_4577_) );
OR2X2 OR2X2_5 ( .A(_4565_), .B(_4577_), .Y(_4578_) );
NOR3X1 NOR3X1_14 ( .A(_4578_), .B(_4576_), .C(_4559_), .Y(_4579_) );
OAI21X1 OAI21X1_55 ( .A(_4559_), .B(_4578_), .C(_4576_), .Y(_4580_) );
NAND2X1 NAND2X1_57 ( .A(_4606__bF_buf1), .B(_4580_), .Y(_4581_) );
NOR2X1 NOR2X1_125 ( .A(_4579_), .B(_4581_), .Y(_4476__27_) );
NOR2X1 NOR2X1_126 ( .A(_4577_), .B(_4565_), .Y(_4582_) );
NAND2X1 NAND2X1_58 ( .A(_4582_), .B(_4531_), .Y(_4583_) );
OAI21X1 OAI21X1_56 ( .A(_4583_), .B(_4576_), .C(concatenador_nonce_28_), .Y(_4584_) );
INVX1 INVX1_19 ( .A(concatenador_nonce_28_), .Y(_4585_) );
NAND2X1 NAND2X1_59 ( .A(_4585_), .B(_4579_), .Y(_4586_) );
AOI21X1 AOI21X1_17 ( .A(_4584_), .B(_4586_), .C(_4501_), .Y(_4476__28_) );
INVX1 INVX1_20 ( .A(concatenador_nonce_29_), .Y(_4587_) );
NAND3X1 NAND3X1_11 ( .A(concatenador_nonce_22_), .B(concatenador_nonce_23_), .C(concatenador_nonce_24_), .Y(_4588_) );
OR2X2 OR2X2_6 ( .A(_4588_), .B(_4577_), .Y(_4589_) );
NOR2X1 NOR2X1_127 ( .A(_4576_), .B(_4585_), .Y(_4590_) );
NOR2X1 NOR2X1_128 ( .A(_4525_), .B(_4551_), .Y(_4591_) );
NAND3X1 NAND3X1_12 ( .A(_4544_), .B(_4590_), .C(_4591_), .Y(_4592_) );
OR2X2 OR2X2_7 ( .A(_4592_), .B(_4589_), .Y(_4593_) );
OAI21X1 OAI21X1_57 ( .A(_4548_), .B(_4593_), .C(_4587_), .Y(_4594_) );
NAND2X1 NAND2X1_60 ( .A(_4606__bF_buf2), .B(_4594_), .Y(_4595_) );
NOR3X1 NOR3X1_15 ( .A(_4593_), .B(_4587_), .C(_4548_), .Y(_4596_) );
NOR2X1 NOR2X1_129 ( .A(_4596_), .B(_4595_), .Y(_4476__29_) );
OAI21X1 OAI21X1_58 ( .A(_4596_), .B(concatenador_nonce_30_), .C(_4606__bF_buf2), .Y(_4597_) );
AOI21X1 AOI21X1_18 ( .A(concatenador_nonce_30_), .B(_4596_), .C(_4597_), .Y(_4476__30_) );
INVX1 INVX1_21 ( .A(concatenador_nonce_30_), .Y(_4598_) );
INVX1 INVX1_22 ( .A(concatenador_nonce_31_), .Y(_4599_) );
NOR2X1 NOR2X1_130 ( .A(_4589_), .B(_4592_), .Y(_4600_) );
NAND3X1 NAND3X1_13 ( .A(concatenador_nonce_29_), .B(_4600_), .C(_4542_), .Y(_4601_) );
NOR3X1 NOR3X1_16 ( .A(_4598_), .B(_4599_), .C(_4601_), .Y(_4602_) );
AOI21X1 AOI21X1_19 ( .A(concatenador_nonce_30_), .B(_4596_), .C(concatenador_nonce_31_), .Y(_4603_) );
NOR3X1 NOR3X1_17 ( .A(_4602_), .B(_4501_), .C(_4603_), .Y(_4476__31_) );
DFFPOSX1 DFFPOSX1_193 ( .CLK(clk_bF_buf72), .D(_4476__0_), .Q(concatenador_nonce_0_) );
DFFPOSX1 DFFPOSX1_194 ( .CLK(clk_bF_buf72), .D(_4476__1_), .Q(concatenador_nonce_1_) );
DFFPOSX1 DFFPOSX1_195 ( .CLK(clk_bF_buf7), .D(_4476__2_), .Q(concatenador_nonce_2_) );
DFFPOSX1 DFFPOSX1_196 ( .CLK(clk_bF_buf69), .D(_4476__3_), .Q(concatenador_nonce_3_) );
DFFPOSX1 DFFPOSX1_197 ( .CLK(clk_bF_buf7), .D(_4476__4_), .Q(concatenador_nonce_4_) );
DFFPOSX1 DFFPOSX1_198 ( .CLK(clk_bF_buf22), .D(_4476__5_), .Q(concatenador_nonce_5_) );
DFFPOSX1 DFFPOSX1_199 ( .CLK(clk_bF_buf22), .D(_4476__6_), .Q(concatenador_nonce_6_) );
DFFPOSX1 DFFPOSX1_200 ( .CLK(clk_bF_buf22), .D(_4476__7_), .Q(concatenador_nonce_7_) );
DFFPOSX1 DFFPOSX1_201 ( .CLK(clk_bF_buf72), .D(_4476__8_), .Q(concatenador_nonce_8_) );
DFFPOSX1 DFFPOSX1_202 ( .CLK(clk_bF_buf67), .D(_4476__9_), .Q(concatenador_nonce_9_) );
DFFPOSX1 DFFPOSX1_203 ( .CLK(clk_bF_buf67), .D(_4476__10_), .Q(concatenador_nonce_10_) );
DFFPOSX1 DFFPOSX1_204 ( .CLK(clk_bF_buf67), .D(_4476__11_), .Q(concatenador_nonce_11_) );
DFFPOSX1 DFFPOSX1_205 ( .CLK(clk_bF_buf67), .D(_4476__12_), .Q(concatenador_nonce_12_) );
DFFPOSX1 DFFPOSX1_206 ( .CLK(clk_bF_buf7), .D(_4476__13_), .Q(concatenador_nonce_13_) );
DFFPOSX1 DFFPOSX1_207 ( .CLK(clk_bF_buf72), .D(_4476__14_), .Q(concatenador_nonce_14_) );
DFFPOSX1 DFFPOSX1_208 ( .CLK(clk_bF_buf72), .D(_4476__15_), .Q(concatenador_nonce_15_) );
DFFPOSX1 DFFPOSX1_209 ( .CLK(clk_bF_buf22), .D(_4476__16_), .Q(concatenador_nonce_16_) );
DFFPOSX1 DFFPOSX1_210 ( .CLK(clk_bF_buf67), .D(_4476__17_), .Q(concatenador_nonce_17_) );
DFFPOSX1 DFFPOSX1_211 ( .CLK(clk_bF_buf72), .D(_4476__18_), .Q(concatenador_nonce_18_) );
DFFPOSX1 DFFPOSX1_212 ( .CLK(clk_bF_buf65), .D(_4476__19_), .Q(concatenador_nonce_19_) );
DFFPOSX1 DFFPOSX1_213 ( .CLK(clk_bF_buf17), .D(_4476__20_), .Q(concatenador_nonce_20_) );
DFFPOSX1 DFFPOSX1_214 ( .CLK(clk_bF_buf50), .D(_4476__21_), .Q(concatenador_nonce_21_) );
DFFPOSX1 DFFPOSX1_215 ( .CLK(clk_bF_buf17), .D(_4476__22_), .Q(concatenador_nonce_22_) );
DFFPOSX1 DFFPOSX1_216 ( .CLK(clk_bF_buf50), .D(_4476__23_), .Q(concatenador_nonce_23_) );
DFFPOSX1 DFFPOSX1_217 ( .CLK(clk_bF_buf50), .D(_4476__24_), .Q(concatenador_nonce_24_) );
DFFPOSX1 DFFPOSX1_218 ( .CLK(clk_bF_buf49), .D(_4476__25_), .Q(concatenador_nonce_25_) );
DFFPOSX1 DFFPOSX1_219 ( .CLK(clk_bF_buf49), .D(_4476__26_), .Q(concatenador_nonce_26_) );
DFFPOSX1 DFFPOSX1_220 ( .CLK(clk_bF_buf49), .D(_4476__27_), .Q(concatenador_nonce_27_) );
DFFPOSX1 DFFPOSX1_221 ( .CLK(clk_bF_buf49), .D(_4476__28_), .Q(concatenador_nonce_28_) );
DFFPOSX1 DFFPOSX1_222 ( .CLK(clk_bF_buf49), .D(_4476__29_), .Q(concatenador_nonce_29_) );
DFFPOSX1 DFFPOSX1_223 ( .CLK(clk_bF_buf17), .D(_4476__30_), .Q(concatenador_nonce_30_) );
DFFPOSX1 DFFPOSX1_224 ( .CLK(clk_bF_buf17), .D(_4476__31_), .Q(concatenador_nonce_31_) );
INVX1 INVX1_23 ( .A(comparador_valid_bF_buf3), .Y(_4647_) );
NAND2X1 NAND2X1_61 ( .A(reset_bF_buf5), .B(_4647_), .Y(_4628_) );
NAND3X1 NAND3X1_14 ( .A(comparador_valid_bF_buf2), .B(reset_bF_buf0), .C(concatenador_nonce_0_), .Y(_4648_) );
INVX1 INVX1_24 ( .A(_4648_), .Y(_4629__0_) );
NAND3X1 NAND3X1_15 ( .A(comparador_valid_bF_buf1), .B(reset_bF_buf0), .C(concatenador_nonce_1_), .Y(_4649_) );
INVX1 INVX1_25 ( .A(_4649_), .Y(_4629__1_) );
NAND3X1 NAND3X1_16 ( .A(comparador_valid_bF_buf3), .B(reset_bF_buf5), .C(concatenador_nonce_2_), .Y(_4650_) );
INVX1 INVX1_26 ( .A(_4650_), .Y(_4629__2_) );
NAND3X1 NAND3X1_17 ( .A(comparador_valid_bF_buf3), .B(reset_bF_buf5), .C(concatenador_nonce_3_), .Y(_4651_) );
INVX1 INVX1_27 ( .A(_4651_), .Y(_4629__3_) );
NAND3X1 NAND3X1_18 ( .A(comparador_valid_bF_buf3), .B(reset_bF_buf5), .C(concatenador_nonce_4_), .Y(_4652_) );
INVX1 INVX1_28 ( .A(_4652_), .Y(_4629__4_) );
NAND3X1 NAND3X1_19 ( .A(comparador_valid_bF_buf2), .B(reset_bF_buf4), .C(concatenador_nonce_5_), .Y(_4653_) );
INVX1 INVX1_29 ( .A(_4653_), .Y(_4629__5_) );
NAND3X1 NAND3X1_20 ( .A(comparador_valid_bF_buf2), .B(reset_bF_buf0), .C(concatenador_nonce_6_), .Y(_4654_) );
INVX1 INVX1_30 ( .A(_4654_), .Y(_4629__6_) );
NAND3X1 NAND3X1_21 ( .A(comparador_valid_bF_buf2), .B(reset_bF_buf4), .C(concatenador_nonce_7_), .Y(_4655_) );
INVX1 INVX1_31 ( .A(_4655_), .Y(_4629__7_) );
NAND3X1 NAND3X1_22 ( .A(comparador_valid_bF_buf1), .B(reset_bF_buf3), .C(concatenador_nonce_8_), .Y(_4656_) );
INVX1 INVX1_32 ( .A(_4656_), .Y(_4629__8_) );
NAND3X1 NAND3X1_23 ( .A(comparador_valid_bF_buf3), .B(reset_bF_buf5), .C(concatenador_nonce_9_), .Y(_4657_) );
INVX1 INVX1_33 ( .A(_4657_), .Y(_4629__9_) );
NAND3X1 NAND3X1_24 ( .A(comparador_valid_bF_buf3), .B(reset_bF_buf1), .C(concatenador_nonce_10_), .Y(_4658_) );
INVX1 INVX1_34 ( .A(_4658_), .Y(_4629__10_) );
NAND3X1 NAND3X1_25 ( .A(comparador_valid_bF_buf3), .B(reset_bF_buf5), .C(concatenador_nonce_11_), .Y(_4659_) );
INVX1 INVX1_35 ( .A(_4659_), .Y(_4629__11_) );
NAND3X1 NAND3X1_26 ( .A(comparador_valid_bF_buf0), .B(reset_bF_buf1), .C(concatenador_nonce_12_), .Y(_4660_) );
INVX1 INVX1_36 ( .A(_4660_), .Y(_4629__12_) );
NAND3X1 NAND3X1_27 ( .A(comparador_valid_bF_buf0), .B(reset_bF_buf3), .C(concatenador_nonce_13_), .Y(_4661_) );
INVX1 INVX1_37 ( .A(_4661_), .Y(_4629__13_) );
NAND3X1 NAND3X1_28 ( .A(comparador_valid_bF_buf1), .B(reset_bF_buf3), .C(concatenador_nonce_14_), .Y(_4662_) );
INVX1 INVX1_38 ( .A(_4662_), .Y(_4629__14_) );
NAND3X1 NAND3X1_29 ( .A(comparador_valid_bF_buf0), .B(reset_bF_buf3), .C(concatenador_nonce_15_), .Y(_4630_) );
INVX1 INVX1_39 ( .A(_4630_), .Y(_4629__15_) );
NAND3X1 NAND3X1_30 ( .A(comparador_valid_bF_buf2), .B(reset_bF_buf0), .C(concatenador_nonce_16_), .Y(_4631_) );
INVX1 INVX1_40 ( .A(_4631_), .Y(_4629__16_) );
NAND3X1 NAND3X1_31 ( .A(comparador_valid_bF_buf0), .B(reset_bF_buf1), .C(concatenador_nonce_17_), .Y(_4632_) );
INVX1 INVX1_41 ( .A(_4632_), .Y(_4629__17_) );
NAND3X1 NAND3X1_32 ( .A(comparador_valid_bF_buf0), .B(reset_bF_buf3), .C(concatenador_nonce_18_), .Y(_4633_) );
INVX1 INVX1_42 ( .A(_4633_), .Y(_4629__18_) );
NAND3X1 NAND3X1_33 ( .A(comparador_valid_bF_buf1), .B(reset_bF_buf0), .C(concatenador_nonce_19_), .Y(_4634_) );
INVX1 INVX1_43 ( .A(_4634_), .Y(_4629__19_) );
NAND3X1 NAND3X1_34 ( .A(comparador_valid_bF_buf4), .B(reset_bF_buf4), .C(concatenador_nonce_20_), .Y(_4635_) );
INVX1 INVX1_44 ( .A(_4635_), .Y(_4629__20_) );
NAND3X1 NAND3X1_35 ( .A(comparador_valid_bF_buf4), .B(reset_bF_buf2), .C(concatenador_nonce_21_), .Y(_4636_) );
INVX1 INVX1_45 ( .A(_4636_), .Y(_4629__21_) );
NAND3X1 NAND3X1_36 ( .A(comparador_valid_bF_buf4), .B(reset_bF_buf2), .C(concatenador_nonce_22_), .Y(_4637_) );
INVX1 INVX1_46 ( .A(_4637_), .Y(_4629__22_) );
NAND3X1 NAND3X1_37 ( .A(comparador_valid_bF_buf4), .B(reset_bF_buf2), .C(concatenador_nonce_23_), .Y(_4638_) );
INVX1 INVX1_47 ( .A(_4638_), .Y(_4629__23_) );
NAND3X1 NAND3X1_38 ( .A(comparador_valid_bF_buf4), .B(reset_bF_buf4), .C(concatenador_nonce_24_), .Y(_4639_) );
INVX1 INVX1_48 ( .A(_4639_), .Y(_4629__24_) );
NAND3X1 NAND3X1_39 ( .A(comparador_valid_bF_buf1), .B(reset_bF_buf3), .C(concatenador_nonce_25_), .Y(_4640_) );
INVX1 INVX1_49 ( .A(_4640_), .Y(_4629__25_) );
NAND3X1 NAND3X1_40 ( .A(comparador_valid_bF_buf0), .B(reset_bF_buf1), .C(concatenador_nonce_26_), .Y(_4641_) );
INVX1 INVX1_50 ( .A(_4641_), .Y(_4629__26_) );
NAND3X1 NAND3X1_41 ( .A(comparador_valid_bF_buf1), .B(reset_bF_buf0), .C(concatenador_nonce_27_), .Y(_4642_) );
INVX1 INVX1_51 ( .A(_4642_), .Y(_4629__27_) );
NAND3X1 NAND3X1_42 ( .A(comparador_valid_bF_buf2), .B(reset_bF_buf4), .C(concatenador_nonce_28_), .Y(_4643_) );
INVX1 INVX1_52 ( .A(_4643_), .Y(_4629__28_) );
NAND3X1 NAND3X1_43 ( .A(comparador_valid_bF_buf2), .B(reset_bF_buf4), .C(concatenador_nonce_29_), .Y(_4644_) );
INVX1 INVX1_53 ( .A(_4644_), .Y(_4629__29_) );
NAND3X1 NAND3X1_44 ( .A(comparador_valid_bF_buf4), .B(reset_bF_buf2), .C(concatenador_nonce_30_), .Y(_4645_) );
INVX1 INVX1_54 ( .A(_4645_), .Y(_4629__30_) );
NAND3X1 NAND3X1_45 ( .A(comparador_valid_bF_buf4), .B(reset_bF_buf2), .C(concatenador_nonce_31_), .Y(_4646_) );
INVX1 INVX1_55 ( .A(_4646_), .Y(_4629__31_) );
DFFPOSX1 DFFPOSX1_225 ( .CLK(clk_bF_buf65), .D(_4629__0_), .Q(_1__0_) );
DFFPOSX1 DFFPOSX1_226 ( .CLK(clk_bF_buf65), .D(_4629__1_), .Q(_1__1_) );
DFFPOSX1 DFFPOSX1_227 ( .CLK(clk_bF_buf67), .D(_4629__2_), .Q(_1__2_) );
DFFPOSX1 DFFPOSX1_228 ( .CLK(clk_bF_buf37), .D(_4629__3_), .Q(_1__3_) );
DFFPOSX1 DFFPOSX1_229 ( .CLK(clk_bF_buf37), .D(_4629__4_), .Q(_1__4_) );
DFFPOSX1 DFFPOSX1_230 ( .CLK(clk_bF_buf49), .D(_4629__5_), .Q(_1__5_) );
DFFPOSX1 DFFPOSX1_231 ( .CLK(clk_bF_buf65), .D(_4629__6_), .Q(_1__6_) );
DFFPOSX1 DFFPOSX1_232 ( .CLK(clk_bF_buf49), .D(_4629__7_), .Q(_1__7_) );
DFFPOSX1 DFFPOSX1_233 ( .CLK(clk_bF_buf65), .D(_4629__8_), .Q(_1__8_) );
DFFPOSX1 DFFPOSX1_234 ( .CLK(clk_bF_buf56), .D(_4629__9_), .Q(_1__9_) );
DFFPOSX1 DFFPOSX1_235 ( .CLK(clk_bF_buf10), .D(_4629__10_), .Q(_1__10_) );
DFFPOSX1 DFFPOSX1_236 ( .CLK(clk_bF_buf26), .D(_4629__11_), .Q(_1__11_) );
DFFPOSX1 DFFPOSX1_237 ( .CLK(clk_bF_buf10), .D(_4629__12_), .Q(_1__12_) );
DFFPOSX1 DFFPOSX1_238 ( .CLK(clk_bF_buf10), .D(_4629__13_), .Q(_1__13_) );
DFFPOSX1 DFFPOSX1_239 ( .CLK(clk_bF_buf72), .D(_4629__14_), .Q(_1__14_) );
DFFPOSX1 DFFPOSX1_240 ( .CLK(clk_bF_buf10), .D(_4629__15_), .Q(_1__15_) );
DFFPOSX1 DFFPOSX1_241 ( .CLK(clk_bF_buf72), .D(_4629__16_), .Q(_1__16_) );
DFFPOSX1 DFFPOSX1_242 ( .CLK(clk_bF_buf10), .D(_4629__17_), .Q(_1__17_) );
DFFPOSX1 DFFPOSX1_243 ( .CLK(clk_bF_buf10), .D(_4629__18_), .Q(_1__18_) );
DFFPOSX1 DFFPOSX1_244 ( .CLK(clk_bF_buf65), .D(_4629__19_), .Q(_1__19_) );
DFFPOSX1 DFFPOSX1_245 ( .CLK(clk_bF_buf17), .D(_4629__20_), .Q(_1__20_) );
DFFPOSX1 DFFPOSX1_246 ( .CLK(clk_bF_buf15), .D(_4629__21_), .Q(_1__21_) );
DFFPOSX1 DFFPOSX1_247 ( .CLK(clk_bF_buf15), .D(_4629__22_), .Q(_1__22_) );
DFFPOSX1 DFFPOSX1_248 ( .CLK(clk_bF_buf15), .D(_4629__23_), .Q(_1__23_) );
DFFPOSX1 DFFPOSX1_249 ( .CLK(clk_bF_buf17), .D(_4629__24_), .Q(_1__24_) );
DFFPOSX1 DFFPOSX1_250 ( .CLK(clk_bF_buf65), .D(_4629__25_), .Q(_1__25_) );
DFFPOSX1 DFFPOSX1_251 ( .CLK(clk_bF_buf10), .D(_4629__26_), .Q(_1__26_) );
DFFPOSX1 DFFPOSX1_252 ( .CLK(clk_bF_buf65), .D(_4629__27_), .Q(_1__27_) );
DFFPOSX1 DFFPOSX1_253 ( .CLK(clk_bF_buf49), .D(_4629__28_), .Q(_1__28_) );
DFFPOSX1 DFFPOSX1_254 ( .CLK(clk_bF_buf49), .D(_4629__29_), .Q(_1__29_) );
DFFPOSX1 DFFPOSX1_255 ( .CLK(clk_bF_buf17), .D(_4629__30_), .Q(_1__30_) );
DFFPOSX1 DFFPOSX1_256 ( .CLK(clk_bF_buf15), .D(_4629__31_), .Q(_1__31_) );
DFFPOSX1 DFFPOSX1_257 ( .CLK(clk_bF_buf66), .D(_4628_), .Q(_0_) );
BUFX2 BUFX2_1 ( .A(_0__bF_buf7), .Y(finished) );
BUFX2 BUFX2_2 ( .A(_1__0_), .Y(nonce_out[0]) );
BUFX2 BUFX2_3 ( .A(_1__1_), .Y(nonce_out[1]) );
BUFX2 BUFX2_4 ( .A(_1__2_), .Y(nonce_out[2]) );
BUFX2 BUFX2_5 ( .A(_1__3_), .Y(nonce_out[3]) );
BUFX2 BUFX2_6 ( .A(_1__4_), .Y(nonce_out[4]) );
BUFX2 BUFX2_7 ( .A(_1__5_), .Y(nonce_out[5]) );
BUFX2 BUFX2_8 ( .A(_1__6_), .Y(nonce_out[6]) );
BUFX2 BUFX2_9 ( .A(_1__7_), .Y(nonce_out[7]) );
BUFX2 BUFX2_10 ( .A(_1__8_), .Y(nonce_out[8]) );
BUFX2 BUFX2_11 ( .A(_1__9_), .Y(nonce_out[9]) );
BUFX2 BUFX2_12 ( .A(_1__10_), .Y(nonce_out[10]) );
BUFX2 BUFX2_13 ( .A(_1__11_), .Y(nonce_out[11]) );
BUFX2 BUFX2_14 ( .A(_1__12_), .Y(nonce_out[12]) );
BUFX2 BUFX2_15 ( .A(_1__13_), .Y(nonce_out[13]) );
BUFX2 BUFX2_16 ( .A(_1__14_), .Y(nonce_out[14]) );
BUFX2 BUFX2_17 ( .A(_1__15_), .Y(nonce_out[15]) );
BUFX2 BUFX2_18 ( .A(_1__16_), .Y(nonce_out[16]) );
BUFX2 BUFX2_19 ( .A(_1__17_), .Y(nonce_out[17]) );
BUFX2 BUFX2_20 ( .A(_1__18_), .Y(nonce_out[18]) );
BUFX2 BUFX2_21 ( .A(_1__19_), .Y(nonce_out[19]) );
BUFX2 BUFX2_22 ( .A(_1__20_), .Y(nonce_out[20]) );
BUFX2 BUFX2_23 ( .A(_1__21_), .Y(nonce_out[21]) );
BUFX2 BUFX2_24 ( .A(_1__22_), .Y(nonce_out[22]) );
BUFX2 BUFX2_25 ( .A(_1__23_), .Y(nonce_out[23]) );
BUFX2 BUFX2_26 ( .A(_1__24_), .Y(nonce_out[24]) );
BUFX2 BUFX2_27 ( .A(_1__25_), .Y(nonce_out[25]) );
BUFX2 BUFX2_28 ( .A(_1__26_), .Y(nonce_out[26]) );
BUFX2 BUFX2_29 ( .A(_1__27_), .Y(nonce_out[27]) );
BUFX2 BUFX2_30 ( .A(_1__28_), .Y(nonce_out[28]) );
BUFX2 BUFX2_31 ( .A(_1__29_), .Y(nonce_out[29]) );
BUFX2 BUFX2_32 ( .A(_1__30_), .Y(nonce_out[30]) );
BUFX2 BUFX2_33 ( .A(_1__31_), .Y(nonce_out[31]) );
INVX4 INVX4_2 ( .A(target[7]), .Y(_54_) );
INVX2 INVX2_6 ( .A(target[6]), .Y(_55_) );
OAI22X1 OAI22X1_1 ( .A(_54_), .B(H_23_), .C(_55_), .D(H_22_), .Y(_56_) );
INVX1 INVX1_56 ( .A(H_23_), .Y(_57_) );
INVX1 INVX1_57 ( .A(H_22_), .Y(_58_) );
OAI22X1 OAI22X1_2 ( .A(_57_), .B(target[7]), .C(target[6]), .D(_58_), .Y(_59_) );
NOR2X1 NOR2X1_131 ( .A(_56_), .B(_59_), .Y(_60_) );
INVX1 INVX1_58 ( .A(H_21_), .Y(_61_) );
INVX1 INVX1_59 ( .A(H_20_), .Y(_62_) );
AOI22X1 AOI22X1_1 ( .A(_61_), .B(target[5]), .C(target[4]), .D(_62_), .Y(_63_) );
INVX2 INVX2_7 ( .A(target[4]), .Y(_64_) );
NOR2X1 NOR2X1_132 ( .A(target[5]), .B(_61_), .Y(_65_) );
AOI21X1 AOI21X1_20 ( .A(_64_), .B(H_20_), .C(_65_), .Y(_66_) );
NAND3X1 NAND3X1_46 ( .A(_63_), .B(_66_), .C(_60_), .Y(_67_) );
INVX2 INVX2_8 ( .A(target[3]), .Y(_68_) );
INVX2 INVX2_9 ( .A(target[2]), .Y(_69_) );
OAI22X1 OAI22X1_3 ( .A(_68_), .B(H_19_), .C(_69_), .D(H_18_), .Y(_70_) );
INVX2 INVX2_10 ( .A(H_19_), .Y(_71_) );
INVX1 INVX1_60 ( .A(H_18_), .Y(_72_) );
OAI22X1 OAI22X1_4 ( .A(_71_), .B(target[3]), .C(target[2]), .D(_72_), .Y(_73_) );
NOR2X1 NOR2X1_133 ( .A(_70_), .B(_73_), .Y(_74_) );
INVX1 INVX1_61 ( .A(H_17_), .Y(_75_) );
NAND2X1 NAND2X1_62 ( .A(target[1]), .B(_75_), .Y(_76_) );
NOR2X1 NOR2X1_134 ( .A(target[1]), .B(_75_), .Y(_77_) );
INVX1 INVX1_62 ( .A(H_16_), .Y(_78_) );
NOR2X1 NOR2X1_135 ( .A(target[0]), .B(_78_), .Y(_79_) );
OAI21X1 OAI21X1_59 ( .A(_77_), .B(_79_), .C(_76_), .Y(_80_) );
NAND2X1 NAND2X1_63 ( .A(target[3]), .B(_71_), .Y(_81_) );
NAND2X1 NAND2X1_64 ( .A(target[2]), .B(_72_), .Y(_82_) );
NOR2X1 NOR2X1_136 ( .A(target[3]), .B(_71_), .Y(_83_) );
OAI21X1 OAI21X1_60 ( .A(_83_), .B(_82_), .C(_81_), .Y(_84_) );
AOI21X1 AOI21X1_21 ( .A(_80_), .B(_74_), .C(_84_), .Y(_85_) );
NOR2X1 NOR2X1_137 ( .A(_65_), .B(_63_), .Y(_86_) );
AOI22X1 AOI22X1_2 ( .A(_57_), .B(target[7]), .C(target[6]), .D(_58_), .Y(_87_) );
AOI21X1 AOI21X1_22 ( .A(H_23_), .B(_54_), .C(_87_), .Y(_88_) );
AOI21X1 AOI21X1_23 ( .A(_86_), .B(_60_), .C(_88_), .Y(_89_) );
OAI21X1 OAI21X1_61 ( .A(_85_), .B(_67_), .C(_89_), .Y(_90_) );
INVX1 INVX1_63 ( .A(H_14_), .Y(_91_) );
OAI22X1 OAI22X1_5 ( .A(_54_), .B(H_15_), .C(target[6]), .D(_91_), .Y(_92_) );
INVX2 INVX2_11 ( .A(H_15_), .Y(_93_) );
OAI22X1 OAI22X1_6 ( .A(_55_), .B(H_14_), .C(target[7]), .D(_93_), .Y(_94_) );
NOR2X1 NOR2X1_138 ( .A(_92_), .B(_94_), .Y(_95_) );
XNOR2X1 XNOR2X1_1 ( .A(target[5]), .B(H_13_), .Y(_96_) );
XNOR2X1 XNOR2X1_2 ( .A(target[4]), .B(H_12_), .Y(_97_) );
NAND3X1 NAND3X1_47 ( .A(_96_), .B(_97_), .C(_95_), .Y(_98_) );
NOR2X1 NOR2X1_139 ( .A(target[3]), .B(H_11_), .Y(_99_) );
INVX1 INVX1_64 ( .A(_99_), .Y(_100_) );
NAND2X1 NAND2X1_65 ( .A(target[3]), .B(H_11_), .Y(_101_) );
XOR2X1 XOR2X1_1 ( .A(target[2]), .B(H_10_), .Y(_102_) );
AOI21X1 AOI21X1_24 ( .A(_100_), .B(_101_), .C(_102_), .Y(_103_) );
INVX1 INVX1_65 ( .A(H_9_), .Y(_104_) );
NAND2X1 NAND2X1_66 ( .A(target[1]), .B(_104_), .Y(_105_) );
INVX1 INVX1_66 ( .A(H_8_), .Y(_106_) );
NOR2X1 NOR2X1_140 ( .A(target[0]), .B(_106_), .Y(_107_) );
NOR2X1 NOR2X1_141 ( .A(target[1]), .B(_104_), .Y(_108_) );
OAI21X1 OAI21X1_62 ( .A(_107_), .B(_108_), .C(_105_), .Y(_109_) );
INVX1 INVX1_67 ( .A(H_11_), .Y(_110_) );
NAND2X1 NAND2X1_67 ( .A(target[3]), .B(_110_), .Y(_111_) );
NOR2X1 NOR2X1_142 ( .A(target[3]), .B(_110_), .Y(_112_) );
OR2X2 OR2X2_8 ( .A(_69_), .B(H_10_), .Y(_113_) );
OAI21X1 OAI21X1_63 ( .A(_113_), .B(_112_), .C(_111_), .Y(_114_) );
AOI21X1 AOI21X1_25 ( .A(_109_), .B(_103_), .C(_114_), .Y(_115_) );
INVX1 INVX1_68 ( .A(H_13_), .Y(_116_) );
NAND2X1 NAND2X1_68 ( .A(target[5]), .B(_116_), .Y(_117_) );
NOR2X1 NOR2X1_143 ( .A(target[5]), .B(_116_), .Y(_118_) );
OR2X2 OR2X2_9 ( .A(_64_), .B(H_12_), .Y(_119_) );
OAI21X1 OAI21X1_64 ( .A(_119_), .B(_118_), .C(_117_), .Y(_120_) );
NAND2X1 NAND2X1_69 ( .A(target[7]), .B(_93_), .Y(_121_) );
NAND2X1 NAND2X1_70 ( .A(H_15_), .B(_54_), .Y(_122_) );
INVX1 INVX1_69 ( .A(_122_), .Y(_123_) );
NAND2X1 NAND2X1_71 ( .A(target[6]), .B(_91_), .Y(_124_) );
OAI21X1 OAI21X1_65 ( .A(_123_), .B(_124_), .C(_121_), .Y(_4_) );
AOI21X1 AOI21X1_26 ( .A(_95_), .B(_120_), .C(_4_), .Y(_5_) );
OAI21X1 OAI21X1_66 ( .A(_115_), .B(_98_), .C(_5_), .Y(_6_) );
AOI22X1 AOI22X1_3 ( .A(_54_), .B(H_23_), .C(_55_), .D(H_22_), .Y(_7_) );
NAND2X1 NAND2X1_72 ( .A(_87_), .B(_7_), .Y(_8_) );
INVX1 INVX1_70 ( .A(target[5]), .Y(_9_) );
NAND2X1 NAND2X1_73 ( .A(H_21_), .B(_9_), .Y(_10_) );
NAND2X1 NAND2X1_74 ( .A(H_20_), .B(_64_), .Y(_11_) );
NAND3X1 NAND3X1_48 ( .A(_10_), .B(_11_), .C(_63_), .Y(_12_) );
NOR2X1 NOR2X1_144 ( .A(_8_), .B(_12_), .Y(_13_) );
AOI22X1 AOI22X1_4 ( .A(_55_), .B(H_14_), .C(target[7]), .D(_93_), .Y(_14_) );
NAND3X1 NAND3X1_49 ( .A(_122_), .B(_124_), .C(_14_), .Y(_15_) );
NAND2X1 NAND2X1_75 ( .A(_96_), .B(_97_), .Y(_16_) );
NOR2X1 NOR2X1_145 ( .A(_16_), .B(_15_), .Y(_17_) );
INVX1 INVX1_71 ( .A(_101_), .Y(_18_) );
XNOR2X1 XNOR2X1_3 ( .A(target[2]), .B(H_10_), .Y(_19_) );
OAI21X1 OAI21X1_67 ( .A(_99_), .B(_18_), .C(_19_), .Y(_20_) );
INVX1 INVX1_72 ( .A(target[0]), .Y(_21_) );
NAND2X1 NAND2X1_76 ( .A(H_8_), .B(_21_), .Y(_22_) );
XNOR2X1 XNOR2X1_4 ( .A(target[1]), .B(H_9_), .Y(_23_) );
NAND2X1 NAND2X1_77 ( .A(target[0]), .B(_106_), .Y(_24_) );
NAND3X1 NAND3X1_50 ( .A(_22_), .B(_24_), .C(_23_), .Y(_25_) );
NOR2X1 NOR2X1_146 ( .A(_20_), .B(_25_), .Y(_26_) );
AOI22X1 AOI22X1_5 ( .A(_68_), .B(H_19_), .C(_69_), .D(H_18_), .Y(_27_) );
NAND3X1 NAND3X1_51 ( .A(_81_), .B(_82_), .C(_27_), .Y(_28_) );
XNOR2X1 XNOR2X1_5 ( .A(target[1]), .B(H_17_), .Y(_29_) );
XNOR2X1 XNOR2X1_6 ( .A(target[0]), .B(H_16_), .Y(_30_) );
NAND2X1 NAND2X1_78 ( .A(_29_), .B(_30_), .Y(_31_) );
NOR2X1 NOR2X1_147 ( .A(_31_), .B(_28_), .Y(_32_) );
AOI22X1 AOI22X1_6 ( .A(_13_), .B(_32_), .C(_26_), .D(_17_), .Y(_33_) );
NAND3X1 NAND3X1_52 ( .A(_90_), .B(_33_), .C(_6_), .Y(_34_) );
NAND2X1 NAND2X1_79 ( .A(comparador_valid_hash), .B(reset_bF_buf2), .Y(_35_) );
NOR2X1 NOR2X1_148 ( .A(_35_), .B(_34_), .Y(_3_) );
INVX2 INVX2_12 ( .A(target[1]), .Y(_36_) );
NOR2X1 NOR2X1_149 ( .A(H_9_), .B(_36_), .Y(_37_) );
NAND2X1 NAND2X1_80 ( .A(H_9_), .B(_36_), .Y(_38_) );
AOI21X1 AOI21X1_27 ( .A(_22_), .B(_38_), .C(_37_), .Y(_39_) );
NOR2X1 NOR2X1_150 ( .A(_39_), .B(_20_), .Y(_40_) );
OAI21X1 OAI21X1_68 ( .A(_40_), .B(_114_), .C(_17_), .Y(_41_) );
AOI22X1 AOI22X1_7 ( .A(_17_), .B(_26_), .C(_41_), .D(_5_), .Y(_42_) );
NOR2X1 NOR2X1_151 ( .A(H_17_), .B(_36_), .Y(_43_) );
NAND2X1 NAND2X1_81 ( .A(H_17_), .B(_36_), .Y(_44_) );
NAND2X1 NAND2X1_82 ( .A(H_16_), .B(_21_), .Y(_45_) );
AOI21X1 AOI21X1_28 ( .A(_44_), .B(_45_), .C(_43_), .Y(_46_) );
INVX1 INVX1_73 ( .A(_81_), .Y(_47_) );
NOR2X1 NOR2X1_152 ( .A(H_18_), .B(_69_), .Y(_48_) );
NAND2X1 NAND2X1_83 ( .A(H_19_), .B(_68_), .Y(_49_) );
AOI21X1 AOI21X1_29 ( .A(_49_), .B(_48_), .C(_47_), .Y(_50_) );
OAI21X1 OAI21X1_69 ( .A(_28_), .B(_46_), .C(_50_), .Y(_51_) );
NAND2X1 NAND2X1_84 ( .A(_13_), .B(_51_), .Y(_52_) );
AOI22X1 AOI22X1_8 ( .A(_13_), .B(_32_), .C(_52_), .D(_89_), .Y(_53_) );
AOI21X1 AOI21X1_30 ( .A(_53_), .B(_42_), .C(_35_), .Y(_2_) );
DFFPOSX1 DFFPOSX1_258 ( .CLK(clk_bF_buf15), .D(_2_), .Q(comparador_next) );
DFFPOSX1 DFFPOSX1_259 ( .CLK(clk_bF_buf15), .D(_3_), .Q(comparador_valid) );
DFFPOSX1 DFFPOSX1_260 ( .CLK(clk_bF_buf69), .D(concatenador_nonce_0_), .Q(concatenador_data_out_0_) );
DFFPOSX1 DFFPOSX1_261 ( .CLK(clk_bF_buf69), .D(concatenador_nonce_1_), .Q(concatenador_data_out_1_) );
DFFPOSX1 DFFPOSX1_262 ( .CLK(clk_bF_buf82), .D(concatenador_nonce_2_), .Q(concatenador_data_out_2_) );
DFFPOSX1 DFFPOSX1_263 ( .CLK(clk_bF_buf77), .D(concatenador_nonce_3_), .Q(concatenador_data_out_3_) );
DFFPOSX1 DFFPOSX1_264 ( .CLK(clk_bF_buf82), .D(concatenador_nonce_4_), .Q(concatenador_data_out_4_) );
DFFPOSX1 DFFPOSX1_265 ( .CLK(clk_bF_buf69), .D(concatenador_nonce_5_), .Q(concatenador_data_out_5_) );
DFFPOSX1 DFFPOSX1_266 ( .CLK(clk_bF_buf12), .D(concatenador_nonce_6_), .Q(concatenador_data_out_6_) );
DFFPOSX1 DFFPOSX1_267 ( .CLK(clk_bF_buf59), .D(concatenador_nonce_7_), .Q(concatenador_data_out_7_) );
DFFPOSX1 DFFPOSX1_268 ( .CLK(clk_bF_buf7), .D(concatenador_nonce_8_), .Q(concatenador_data_out_8_) );
DFFPOSX1 DFFPOSX1_269 ( .CLK(clk_bF_buf77), .D(concatenador_nonce_9_), .Q(concatenador_data_out_9_) );
DFFPOSX1 DFFPOSX1_270 ( .CLK(clk_bF_buf82), .D(concatenador_nonce_10_), .Q(concatenador_data_out_10_) );
DFFPOSX1 DFFPOSX1_271 ( .CLK(clk_bF_buf66), .D(concatenador_nonce_11_), .Q(concatenador_data_out_11_) );
DFFPOSX1 DFFPOSX1_272 ( .CLK(clk_bF_buf77), .D(concatenador_nonce_12_), .Q(concatenador_data_out_12_) );
DFFPOSX1 DFFPOSX1_273 ( .CLK(clk_bF_buf7), .D(concatenador_nonce_13_), .Q(concatenador_data_out_13_) );
DFFPOSX1 DFFPOSX1_274 ( .CLK(clk_bF_buf7), .D(concatenador_nonce_14_), .Q(concatenador_data_out_14_) );
DFFPOSX1 DFFPOSX1_275 ( .CLK(clk_bF_buf22), .D(concatenador_nonce_15_), .Q(concatenador_data_out_15_) );
DFFPOSX1 DFFPOSX1_276 ( .CLK(clk_bF_buf69), .D(concatenador_nonce_16_), .Q(concatenador_data_out_16_) );
DFFPOSX1 DFFPOSX1_277 ( .CLK(clk_bF_buf77), .D(concatenador_nonce_17_), .Q(concatenador_data_out_17_) );
DFFPOSX1 DFFPOSX1_278 ( .CLK(clk_bF_buf82), .D(concatenador_nonce_18_), .Q(concatenador_data_out_18_) );
DFFPOSX1 DFFPOSX1_279 ( .CLK(clk_bF_buf7), .D(concatenador_nonce_19_), .Q(concatenador_data_out_19_) );
DFFPOSX1 DFFPOSX1_280 ( .CLK(clk_bF_buf69), .D(concatenador_nonce_20_), .Q(concatenador_data_out_20_) );
DFFPOSX1 DFFPOSX1_281 ( .CLK(clk_bF_buf50), .D(concatenador_nonce_21_), .Q(concatenador_data_out_21_) );
DFFPOSX1 DFFPOSX1_282 ( .CLK(clk_bF_buf50), .D(concatenador_nonce_22_), .Q(concatenador_data_out_22_) );
DFFPOSX1 DFFPOSX1_283 ( .CLK(clk_bF_buf17), .D(concatenador_nonce_23_), .Q(concatenador_data_out_23_) );
DFFPOSX1 DFFPOSX1_284 ( .CLK(clk_bF_buf59), .D(concatenador_nonce_24_), .Q(concatenador_data_out_24_) );
DFFPOSX1 DFFPOSX1_285 ( .CLK(clk_bF_buf8), .D(concatenador_nonce_25_), .Q(concatenador_data_out_25_) );
DFFPOSX1 DFFPOSX1_286 ( .CLK(clk_bF_buf47), .D(concatenador_nonce_26_), .Q(concatenador_data_out_26_) );
DFFPOSX1 DFFPOSX1_287 ( .CLK(clk_bF_buf47), .D(concatenador_nonce_27_), .Q(concatenador_data_out_27_) );
DFFPOSX1 DFFPOSX1_288 ( .CLK(clk_bF_buf22), .D(concatenador_nonce_28_), .Q(concatenador_data_out_28_) );
DFFPOSX1 DFFPOSX1_289 ( .CLK(clk_bF_buf50), .D(concatenador_nonce_29_), .Q(concatenador_data_out_29_) );
DFFPOSX1 DFFPOSX1_290 ( .CLK(clk_bF_buf17), .D(concatenador_nonce_30_), .Q(concatenador_data_out_30_) );
DFFPOSX1 DFFPOSX1_291 ( .CLK(clk_bF_buf15), .D(concatenador_nonce_31_), .Q(concatenador_data_out_31_) );
DFFPOSX1 DFFPOSX1_292 ( .CLK(clk_bF_buf39), .D(concatenador_bloque_0_), .Q(concatenador_data_out_32_) );
DFFPOSX1 DFFPOSX1_293 ( .CLK(clk_bF_buf64), .D(concatenador_bloque_1_), .Q(concatenador_data_out_33_) );
DFFPOSX1 DFFPOSX1_294 ( .CLK(clk_bF_buf79), .D(concatenador_bloque_2_), .Q(concatenador_data_out_34_) );
DFFPOSX1 DFFPOSX1_295 ( .CLK(clk_bF_buf34), .D(concatenador_bloque_3_), .Q(concatenador_data_out_35_) );
DFFPOSX1 DFFPOSX1_296 ( .CLK(clk_bF_buf34), .D(concatenador_bloque_4_), .Q(concatenador_data_out_36_) );
DFFPOSX1 DFFPOSX1_297 ( .CLK(clk_bF_buf42), .D(concatenador_bloque_5_), .Q(concatenador_data_out_37_) );
DFFPOSX1 DFFPOSX1_298 ( .CLK(clk_bF_buf42), .D(concatenador_bloque_6_), .Q(concatenador_data_out_38_) );
DFFPOSX1 DFFPOSX1_299 ( .CLK(clk_bF_buf32), .D(concatenador_bloque_7_), .Q(concatenador_data_out_39_) );
DFFPOSX1 DFFPOSX1_300 ( .CLK(clk_bF_buf54), .D(concatenador_bloque_8_), .Q(concatenador_data_out_40_) );
DFFPOSX1 DFFPOSX1_301 ( .CLK(clk_bF_buf39), .D(concatenador_bloque_9_), .Q(concatenador_data_out_41_) );
DFFPOSX1 DFFPOSX1_302 ( .CLK(clk_bF_buf34), .D(concatenador_bloque_10_), .Q(concatenador_data_out_42_) );
DFFPOSX1 DFFPOSX1_303 ( .CLK(clk_bF_buf30), .D(concatenador_bloque_11_), .Q(concatenador_data_out_43_) );
DFFPOSX1 DFFPOSX1_304 ( .CLK(clk_bF_buf52), .D(concatenador_bloque_12_), .Q(concatenador_data_out_44_) );
DFFPOSX1 DFFPOSX1_305 ( .CLK(clk_bF_buf66), .D(concatenador_bloque_13_), .Q(concatenador_data_out_45_) );
DFFPOSX1 DFFPOSX1_306 ( .CLK(clk_bF_buf82), .D(concatenador_bloque_14_), .Q(concatenador_data_out_46_) );
DFFPOSX1 DFFPOSX1_307 ( .CLK(clk_bF_buf22), .D(concatenador_bloque_15_), .Q(concatenador_data_out_47_) );
DFFPOSX1 DFFPOSX1_308 ( .CLK(clk_bF_buf60), .D(concatenador_bloque_16_), .Q(concatenador_data_out_48_) );
DFFPOSX1 DFFPOSX1_309 ( .CLK(clk_bF_buf74), .D(concatenador_bloque_17_), .Q(concatenador_data_out_49_) );
DFFPOSX1 DFFPOSX1_310 ( .CLK(clk_bF_buf36), .D(concatenador_bloque_18_), .Q(concatenador_data_out_50_) );
DFFPOSX1 DFFPOSX1_311 ( .CLK(clk_bF_buf79), .D(concatenador_bloque_19_), .Q(concatenador_data_out_51_) );
DFFPOSX1 DFFPOSX1_312 ( .CLK(clk_bF_buf36), .D(concatenador_bloque_20_), .Q(concatenador_data_out_52_) );
DFFPOSX1 DFFPOSX1_313 ( .CLK(clk_bF_buf66), .D(concatenador_bloque_21_), .Q(concatenador_data_out_53_) );
DFFPOSX1 DFFPOSX1_314 ( .CLK(clk_bF_buf72), .D(concatenador_bloque_22_), .Q(concatenador_data_out_54_) );
DFFPOSX1 DFFPOSX1_315 ( .CLK(clk_bF_buf22), .D(concatenador_bloque_23_), .Q(concatenador_data_out_55_) );
DFFPOSX1 DFFPOSX1_316 ( .CLK(clk_bF_buf54), .D(concatenador_bloque_24_), .Q(concatenador_data_out_56_) );
DFFPOSX1 DFFPOSX1_317 ( .CLK(clk_bF_buf55), .D(concatenador_bloque_25_), .Q(concatenador_data_out_57_) );
DFFPOSX1 DFFPOSX1_318 ( .CLK(clk_bF_buf74), .D(concatenador_bloque_26_), .Q(concatenador_data_out_58_) );
DFFPOSX1 DFFPOSX1_319 ( .CLK(clk_bF_buf44), .D(concatenador_bloque_27_), .Q(concatenador_data_out_59_) );
DFFPOSX1 DFFPOSX1_320 ( .CLK(clk_bF_buf36), .D(concatenador_bloque_28_), .Q(concatenador_data_out_60_) );
DFFPOSX1 DFFPOSX1_321 ( .CLK(clk_bF_buf47), .D(concatenador_bloque_29_), .Q(concatenador_data_out_61_) );
DFFPOSX1 DFFPOSX1_322 ( .CLK(clk_bF_buf32), .D(concatenador_bloque_30_), .Q(concatenador_data_out_62_) );
DFFPOSX1 DFFPOSX1_323 ( .CLK(clk_bF_buf77), .D(concatenador_bloque_31_), .Q(concatenador_data_out_63_) );
DFFPOSX1 DFFPOSX1_324 ( .CLK(clk_bF_buf45), .D(concatenador_bloque_32_), .Q(concatenador_data_out_64_) );
DFFPOSX1 DFFPOSX1_325 ( .CLK(clk_bF_buf58), .D(concatenador_bloque_33_), .Q(concatenador_data_out_65_) );
DFFPOSX1 DFFPOSX1_326 ( .CLK(clk_bF_buf74), .D(concatenador_bloque_34_), .Q(concatenador_data_out_66_) );
DFFPOSX1 DFFPOSX1_327 ( .CLK(clk_bF_buf34), .D(concatenador_bloque_35_), .Q(concatenador_data_out_67_) );
DFFPOSX1 DFFPOSX1_328 ( .CLK(clk_bF_buf20), .D(concatenador_bloque_36_), .Q(concatenador_data_out_68_) );
DFFPOSX1 DFFPOSX1_329 ( .CLK(clk_bF_buf52), .D(concatenador_bloque_37_), .Q(concatenador_data_out_69_) );
DFFPOSX1 DFFPOSX1_330 ( .CLK(clk_bF_buf82), .D(concatenador_bloque_38_), .Q(concatenador_data_out_70_) );
DFFPOSX1 DFFPOSX1_331 ( .CLK(clk_bF_buf67), .D(concatenador_bloque_39_), .Q(concatenador_data_out_71_) );
DFFPOSX1 DFFPOSX1_332 ( .CLK(clk_bF_buf34), .D(concatenador_bloque_40_), .Q(concatenador_data_out_72_) );
DFFPOSX1 DFFPOSX1_333 ( .CLK(clk_bF_buf45), .D(concatenador_bloque_41_), .Q(concatenador_data_out_73_) );
DFFPOSX1 DFFPOSX1_334 ( .CLK(clk_bF_buf70), .D(concatenador_bloque_42_), .Q(concatenador_data_out_74_) );
DFFPOSX1 DFFPOSX1_335 ( .CLK(clk_bF_buf13), .D(concatenador_bloque_43_), .Q(concatenador_data_out_75_) );
DFFPOSX1 DFFPOSX1_336 ( .CLK(clk_bF_buf20), .D(concatenador_bloque_44_), .Q(concatenador_data_out_76_) );
DFFPOSX1 DFFPOSX1_337 ( .CLK(clk_bF_buf52), .D(concatenador_bloque_45_), .Q(concatenador_data_out_77_) );
DFFPOSX1 DFFPOSX1_338 ( .CLK(clk_bF_buf82), .D(concatenador_bloque_46_), .Q(concatenador_data_out_78_) );
DFFPOSX1 DFFPOSX1_339 ( .CLK(clk_bF_buf77), .D(concatenador_bloque_47_), .Q(concatenador_data_out_79_) );
DFFPOSX1 DFFPOSX1_340 ( .CLK(clk_bF_buf60), .D(concatenador_bloque_48_), .Q(concatenador_data_out_80_) );
DFFPOSX1 DFFPOSX1_341 ( .CLK(clk_bF_buf55), .D(concatenador_bloque_49_), .Q(concatenador_data_out_81_) );
DFFPOSX1 DFFPOSX1_342 ( .CLK(clk_bF_buf27), .D(concatenador_bloque_50_), .Q(concatenador_data_out_82_) );
DFFPOSX1 DFFPOSX1_343 ( .CLK(clk_bF_buf30), .D(concatenador_bloque_51_), .Q(concatenador_data_out_83_) );
DFFPOSX1 DFFPOSX1_344 ( .CLK(clk_bF_buf42), .D(concatenador_bloque_52_), .Q(concatenador_data_out_84_) );
DFFPOSX1 DFFPOSX1_345 ( .CLK(clk_bF_buf39), .D(concatenador_bloque_53_), .Q(concatenador_data_out_85_) );
DFFPOSX1 DFFPOSX1_346 ( .CLK(clk_bF_buf42), .D(concatenador_bloque_54_), .Q(concatenador_data_out_86_) );
DFFPOSX1 DFFPOSX1_347 ( .CLK(clk_bF_buf77), .D(concatenador_bloque_55_), .Q(concatenador_data_out_87_) );
DFFPOSX1 DFFPOSX1_348 ( .CLK(clk_bF_buf16), .D(concatenador_bloque_56_), .Q(concatenador_data_out_88_) );
DFFPOSX1 DFFPOSX1_349 ( .CLK(clk_bF_buf27), .D(concatenador_bloque_57_), .Q(concatenador_data_out_89_) );
DFFPOSX1 DFFPOSX1_350 ( .CLK(clk_bF_buf27), .D(concatenador_bloque_58_), .Q(concatenador_data_out_90_) );
DFFPOSX1 DFFPOSX1_351 ( .CLK(clk_bF_buf13), .D(concatenador_bloque_59_), .Q(concatenador_data_out_91_) );
DFFPOSX1 DFFPOSX1_352 ( .CLK(clk_bF_buf79), .D(concatenador_bloque_60_), .Q(concatenador_data_out_92_) );
DFFPOSX1 DFFPOSX1_353 ( .CLK(clk_bF_buf52), .D(concatenador_bloque_61_), .Q(concatenador_data_out_93_) );
DFFPOSX1 DFFPOSX1_354 ( .CLK(clk_bF_buf47), .D(concatenador_bloque_62_), .Q(concatenador_data_out_94_) );
DFFPOSX1 DFFPOSX1_355 ( .CLK(clk_bF_buf66), .D(concatenador_bloque_63_), .Q(concatenador_data_out_95_) );
DFFPOSX1 DFFPOSX1_356 ( .CLK(clk_bF_buf74), .D(concatenador_bloque_64_), .Q(concatenador_data_out_96_) );
DFFPOSX1 DFFPOSX1_357 ( .CLK(clk_bF_buf64), .D(concatenador_bloque_65_), .Q(concatenador_data_out_97_) );
DFFPOSX1 DFFPOSX1_358 ( .CLK(clk_bF_buf44), .D(concatenador_bloque_66_), .Q(concatenador_data_out_98_) );
DFFPOSX1 DFFPOSX1_359 ( .CLK(clk_bF_buf20), .D(concatenador_bloque_67_), .Q(concatenador_data_out_99_) );
DFFPOSX1 DFFPOSX1_360 ( .CLK(clk_bF_buf42), .D(concatenador_bloque_68_), .Q(concatenador_data_out_100_) );
DFFPOSX1 DFFPOSX1_361 ( .CLK(clk_bF_buf16), .D(concatenador_bloque_69_), .Q(concatenador_data_out_101_) );
DFFPOSX1 DFFPOSX1_362 ( .CLK(clk_bF_buf42), .D(concatenador_bloque_70_), .Q(concatenador_data_out_102_) );
DFFPOSX1 DFFPOSX1_363 ( .CLK(clk_bF_buf66), .D(concatenador_bloque_71_), .Q(concatenador_data_out_103_) );
DFFPOSX1 DFFPOSX1_364 ( .CLK(clk_bF_buf27), .D(concatenador_bloque_72_), .Q(concatenador_data_out_104_) );
DFFPOSX1 DFFPOSX1_365 ( .CLK(clk_bF_buf36), .D(concatenador_bloque_73_), .Q(concatenador_data_out_105_) );
DFFPOSX1 DFFPOSX1_366 ( .CLK(clk_bF_buf27), .D(concatenador_bloque_74_), .Q(concatenador_data_out_106_) );
DFFPOSX1 DFFPOSX1_367 ( .CLK(clk_bF_buf58), .D(concatenador_bloque_75_), .Q(concatenador_data_out_107_) );
DFFPOSX1 DFFPOSX1_368 ( .CLK(clk_bF_buf67), .D(concatenador_bloque_76_), .Q(concatenador_data_out_108_) );
DFFPOSX1 DFFPOSX1_369 ( .CLK(clk_bF_buf6), .D(concatenador_bloque_77_), .Q(concatenador_data_out_109_) );
DFFPOSX1 DFFPOSX1_370 ( .CLK(clk_bF_buf52), .D(concatenador_bloque_78_), .Q(concatenador_data_out_110_) );
DFFPOSX1 DFFPOSX1_371 ( .CLK(clk_bF_buf77), .D(concatenador_bloque_79_), .Q(concatenador_data_out_111_) );
DFFPOSX1 DFFPOSX1_372 ( .CLK(clk_bF_buf60), .D(concatenador_bloque_80_), .Q(concatenador_data_out_112_) );
DFFPOSX1 DFFPOSX1_373 ( .CLK(clk_bF_buf52), .D(concatenador_bloque_81_), .Q(concatenador_data_out_113_) );
DFFPOSX1 DFFPOSX1_374 ( .CLK(clk_bF_buf30), .D(concatenador_bloque_82_), .Q(concatenador_data_out_114_) );
DFFPOSX1 DFFPOSX1_375 ( .CLK(clk_bF_buf79), .D(concatenador_bloque_83_), .Q(concatenador_data_out_115_) );
DFFPOSX1 DFFPOSX1_376 ( .CLK(clk_bF_buf34), .D(concatenador_bloque_84_), .Q(concatenador_data_out_116_) );
DFFPOSX1 DFFPOSX1_377 ( .CLK(clk_bF_buf47), .D(concatenador_bloque_85_), .Q(concatenador_data_out_117_) );
DFFPOSX1 DFFPOSX1_378 ( .CLK(clk_bF_buf6), .D(concatenador_bloque_86_), .Q(concatenador_data_out_118_) );
DFFPOSX1 DFFPOSX1_379 ( .CLK(clk_bF_buf22), .D(concatenador_bloque_87_), .Q(concatenador_data_out_119_) );
DFFPOSX1 DFFPOSX1_380 ( .CLK(clk_bF_buf70), .D(concatenador_bloque_88_), .Q(concatenador_data_out_120_) );
DFFPOSX1 DFFPOSX1_381 ( .CLK(clk_bF_buf38), .D(concatenador_bloque_89_), .Q(concatenador_data_out_121_) );
DFFPOSX1 DFFPOSX1_382 ( .CLK(clk_bF_buf0), .D(concatenador_bloque_90_), .Q(concatenador_data_out_122_) );
DFFPOSX1 DFFPOSX1_383 ( .CLK(clk_bF_buf45), .D(concatenador_bloque_91_), .Q(concatenador_data_out_123_) );
DFFPOSX1 DFFPOSX1_384 ( .CLK(clk_bF_buf42), .D(concatenador_bloque_92_), .Q(concatenador_data_out_124_) );
DFFPOSX1 DFFPOSX1_385 ( .CLK(clk_bF_buf20), .D(concatenador_bloque_93_), .Q(concatenador_data_out_125_) );
DFFPOSX1 DFFPOSX1_386 ( .CLK(clk_bF_buf69), .D(concatenador_bloque_94_), .Q(concatenador_data_out_126_) );
DFFPOSX1 DFFPOSX1_387 ( .CLK(clk_bF_buf66), .D(concatenador_bloque_95_), .Q(concatenador_data_out_127_) );
INVX8 INVX8_1 ( .A(micro_hash_ucr_pipe68), .Y(_4199_) );
INVX8 INVX8_2 ( .A(micro_hash_ucr_c_3_bF_buf3_), .Y(_4200_) );
INVX8 INVX8_3 ( .A(micro_hash_ucr_pipe67), .Y(_4201_) );
NOR2X1 NOR2X1_153 ( .A(_4200_), .B(_4201__bF_buf2), .Y(_4202_) );
NAND2X1 NAND2X1_85 ( .A(micro_hash_ucr_c_3_bF_buf2_), .B(micro_hash_ucr_pipe63_bF_buf2), .Y(_4203_) );
INVX8 INVX8_4 ( .A(micro_hash_ucr_pipe63_bF_buf1), .Y(_4204_) );
INVX8 INVX8_5 ( .A(micro_hash_ucr_b_7_bF_buf3_), .Y(_4205_) );
NAND2X1 NAND2X1_86 ( .A(micro_hash_ucr_pipe62_bF_buf3), .B(_4205_), .Y(_4206_) );
INVX8 INVX8_6 ( .A(micro_hash_ucr_pipe62_bF_buf2), .Y(_4207_) );
INVX8 INVX8_7 ( .A(micro_hash_ucr_pipe61_bF_buf2), .Y(_4208_) );
NOR2X1 NOR2X1_154 ( .A(micro_hash_ucr_c_3_bF_buf1_), .B(_4208_), .Y(_4209_) );
INVX8 INVX8_8 ( .A(micro_hash_ucr_pipe60_bF_buf4), .Y(_4210_) );
INVX8 INVX8_9 ( .A(micro_hash_ucr_pipe58_bF_buf0), .Y(_4211_) );
INVX8 INVX8_10 ( .A(micro_hash_ucr_pipe57_bF_buf0), .Y(_4212_) );
NAND2X1 NAND2X1_87 ( .A(micro_hash_ucr_b_7_bF_buf2_), .B(micro_hash_ucr_pipe54_bF_buf2), .Y(_4213_) );
INVX8 INVX8_11 ( .A(micro_hash_ucr_pipe52_bF_buf2), .Y(_4214_) );
INVX8 INVX8_12 ( .A(micro_hash_ucr_pipe50_bF_buf0), .Y(_4215_) );
NAND2X1 NAND2X1_88 ( .A(micro_hash_ucr_c_3_bF_buf0_), .B(micro_hash_ucr_pipe49_bF_buf3), .Y(_4216_) );
INVX8 INVX8_13 ( .A(micro_hash_ucr_pipe48_bF_buf3), .Y(_4217_) );
INVX8 INVX8_14 ( .A(micro_hash_ucr_pipe46_bF_buf2), .Y(_4218_) );
INVX8 INVX8_15 ( .A(micro_hash_ucr_pipe44_bF_buf2), .Y(_4219_) );
INVX8 INVX8_16 ( .A(micro_hash_ucr_pipe42_bF_buf1), .Y(_4220_) );
NAND2X1 NAND2X1_89 ( .A(micro_hash_ucr_c_3_bF_buf3_), .B(micro_hash_ucr_pipe41_bF_buf1), .Y(_4221_) );
NAND2X1 NAND2X1_90 ( .A(micro_hash_ucr_c_3_bF_buf2_), .B(micro_hash_ucr_pipe39), .Y(_4222_) );
NAND2X1 NAND2X1_91 ( .A(micro_hash_ucr_c_3_bF_buf1_), .B(micro_hash_ucr_pipe37_bF_buf0), .Y(_4223_) );
INVX8 INVX8_17 ( .A(micro_hash_ucr_pipe36_bF_buf1), .Y(_4224_) );
INVX8 INVX8_18 ( .A(micro_hash_ucr_pipe34_bF_buf2), .Y(_4225_) );
INVX8 INVX8_19 ( .A(micro_hash_ucr_pipe32_bF_buf3), .Y(_4226_) );
NAND2X1 NAND2X1_92 ( .A(micro_hash_ucr_c_3_bF_buf0_), .B(micro_hash_ucr_pipe31_bF_buf1), .Y(_4227_) );
INVX8 INVX8_20 ( .A(micro_hash_ucr_pipe30_bF_buf2), .Y(_4228_) );
INVX8 INVX8_21 ( .A(micro_hash_ucr_pipe27_bF_buf1), .Y(_4229_) );
INVX8 INVX8_22 ( .A(micro_hash_ucr_pipe26_bF_buf1), .Y(_4230_) );
NOR2X1 NOR2X1_155 ( .A(_4205_), .B(_4230__bF_buf2), .Y(_4231_) );
NAND2X1 NAND2X1_93 ( .A(micro_hash_ucr_c_3_bF_buf3_), .B(micro_hash_ucr_pipe25_bF_buf3), .Y(_4232_) );
INVX8 INVX8_23 ( .A(micro_hash_ucr_pipe24_bF_buf0), .Y(_4233_) );
INVX8 INVX8_24 ( .A(micro_hash_ucr_pipe23), .Y(_4234_) );
NOR2X1 NOR2X1_156 ( .A(micro_hash_ucr_c_3_bF_buf2_), .B(_4234__bF_buf2), .Y(_4235_) );
INVX8 INVX8_25 ( .A(micro_hash_ucr_pipe21), .Y(_4236_) );
INVX8 INVX8_26 ( .A(micro_hash_ucr_pipe20_bF_buf3), .Y(_4237_) );
INVX8 INVX8_27 ( .A(micro_hash_ucr_pipe17), .Y(_4238_) );
INVX8 INVX8_28 ( .A(micro_hash_ucr_pipe16), .Y(_4239_) );
INVX8 INVX8_29 ( .A(micro_hash_ucr_pipe15), .Y(_4240_) );
INVX8 INVX8_30 ( .A(micro_hash_ucr_pipe14), .Y(_4241_) );
INVX4 INVX4_3 ( .A(micro_hash_ucr_pipe13), .Y(_4242_) );
INVX8 INVX8_31 ( .A(micro_hash_ucr_pipe10), .Y(_4243_) );
NOR2X1 NOR2X1_157 ( .A(micro_hash_ucr_pipe11), .B(_4243_), .Y(_4244_) );
OAI21X1 OAI21X1_70 ( .A(_4244_), .B(micro_hash_ucr_pipe12_bF_buf0), .C(_4242_), .Y(_4245_) );
NAND2X1 NAND2X1_94 ( .A(_4241__bF_buf3), .B(_4245_), .Y(_4246_) );
NAND2X1 NAND2X1_95 ( .A(_4240_), .B(_4246_), .Y(_4247_) );
NAND2X1 NAND2X1_96 ( .A(_4239__bF_buf3), .B(_4247_), .Y(_4248_) );
AOI21X1 AOI21X1_31 ( .A(_4238__bF_buf1), .B(_4248_), .C(micro_hash_ucr_pipe18_bF_buf1), .Y(_4249_) );
OAI21X1 OAI21X1_71 ( .A(_4249_), .B(micro_hash_ucr_pipe19), .C(_4237__bF_buf2), .Y(_4250_) );
AOI21X1 AOI21X1_32 ( .A(_4236__bF_buf0), .B(_4250_), .C(micro_hash_ucr_pipe22_bF_buf0), .Y(_4251_) );
INVX4 INVX4_4 ( .A(micro_hash_ucr_pipe6), .Y(_4252_) );
NOR2X1 NOR2X1_158 ( .A(micro_hash_ucr_pipe8), .B(_4252_), .Y(_4253_) );
INVX2 INVX2_13 ( .A(micro_hash_ucr_pipe7), .Y(_4254_) );
INVX4 INVX4_5 ( .A(micro_hash_ucr_pipe9), .Y(_4255_) );
OAI21X1 OAI21X1_72 ( .A(_4254_), .B(micro_hash_ucr_pipe8), .C(_4255_), .Y(_4256_) );
OAI21X1 OAI21X1_73 ( .A(_4256_), .B(_4253_), .C(_4243_), .Y(_4257_) );
INVX8 INVX8_32 ( .A(micro_hash_ucr_pipe12_bF_buf0), .Y(_4258_) );
NAND2X1 NAND2X1_97 ( .A(_4258_), .B(_4241__bF_buf0), .Y(_4259_) );
NOR2X1 NOR2X1_159 ( .A(_4259_), .B(_4257_), .Y(_4260_) );
NAND2X1 NAND2X1_98 ( .A(_4239__bF_buf1), .B(_4260_), .Y(_4261_) );
INVX8 INVX8_33 ( .A(micro_hash_ucr_pipe22_bF_buf3), .Y(_4262_) );
NOR2X1 NOR2X1_160 ( .A(micro_hash_ucr_pipe18_bF_buf0), .B(micro_hash_ucr_pipe20_bF_buf0), .Y(_4263_) );
NAND2X1 NAND2X1_99 ( .A(_4262__bF_buf4), .B(_4263_), .Y(_4264_) );
OAI21X1 OAI21X1_74 ( .A(_4261_), .B(_4264_), .C(_4205_), .Y(_4265_) );
NAND2X1 NAND2X1_100 ( .A(_4254_), .B(_4255_), .Y(_4266_) );
INVX2 INVX2_14 ( .A(_4266_), .Y(_4267_) );
INVX1 INVX1_74 ( .A(_4253_), .Y(_4268_) );
NOR2X1 NOR2X1_161 ( .A(H_15_), .B(_4268_), .Y(_4269_) );
NOR2X1 NOR2X1_162 ( .A(micro_hash_ucr_pipe19), .B(micro_hash_ucr_pipe21), .Y(_4270_) );
NOR2X1 NOR2X1_163 ( .A(micro_hash_ucr_pipe13), .B(micro_hash_ucr_pipe15), .Y(_4271_) );
NOR2X1 NOR2X1_164 ( .A(micro_hash_ucr_pipe11), .B(_4256_), .Y(_4272_) );
NAND2X1 NAND2X1_101 ( .A(_4271_), .B(_4272_), .Y(_4273_) );
NOR2X1 NOR2X1_165 ( .A(micro_hash_ucr_pipe17), .B(_4273_), .Y(_4274_) );
NAND2X1 NAND2X1_102 ( .A(_4270_), .B(_4274_), .Y(_4275_) );
AOI22X1 AOI22X1_9 ( .A(_4267_), .B(_4269_), .C(_4275_), .D(_4200_), .Y(_4276_) );
INVX4 INVX4_6 ( .A(micro_hash_ucr_pipe11), .Y(_4277_) );
OAI21X1 OAI21X1_75 ( .A(_4277_), .B(micro_hash_ucr_pipe12_bF_buf1), .C(_4242_), .Y(_4278_) );
NAND2X1 NAND2X1_103 ( .A(_4241__bF_buf0), .B(_4278_), .Y(_4279_) );
INVX1 INVX1_75 ( .A(_4279_), .Y(_4280_) );
OAI21X1 OAI21X1_76 ( .A(_4280_), .B(micro_hash_ucr_pipe15), .C(_4239__bF_buf0), .Y(_205_) );
AOI21X1 AOI21X1_33 ( .A(_4238__bF_buf1), .B(_205_), .C(micro_hash_ucr_pipe18_bF_buf1), .Y(_206_) );
OAI21X1 OAI21X1_77 ( .A(_206_), .B(micro_hash_ucr_pipe19), .C(_4237__bF_buf2), .Y(_207_) );
NAND2X1 NAND2X1_104 ( .A(_4236__bF_buf0), .B(_207_), .Y(_208_) );
NOR2X1 NOR2X1_166 ( .A(micro_hash_ucr_pipe22_bF_buf0), .B(_4200_), .Y(_209_) );
AOI22X1 AOI22X1_10 ( .A(_4265_), .B(_4276_), .C(_208_), .D(_209_), .Y(_210_) );
OAI21X1 OAI21X1_78 ( .A(_4251_), .B(_4205_), .C(_210_), .Y(_211_) );
NOR2X1 NOR2X1_167 ( .A(micro_hash_ucr_pipe23), .B(_211_), .Y(_212_) );
OAI21X1 OAI21X1_79 ( .A(_212_), .B(_4235_), .C(_4233__bF_buf3), .Y(_213_) );
OAI21X1 OAI21X1_80 ( .A(micro_hash_ucr_b_7_bF_buf1_), .B(_4233__bF_buf2), .C(_213_), .Y(_214_) );
OR2X2 OR2X2_10 ( .A(_214_), .B(micro_hash_ucr_pipe25_bF_buf3), .Y(_215_) );
AOI21X1 AOI21X1_34 ( .A(_4232_), .B(_215_), .C(micro_hash_ucr_pipe26_bF_buf3), .Y(_216_) );
OAI21X1 OAI21X1_81 ( .A(_216_), .B(_4231_), .C(_4229_), .Y(_217_) );
AOI21X1 AOI21X1_35 ( .A(micro_hash_ucr_c_3_bF_buf1_), .B(micro_hash_ucr_pipe27_bF_buf3), .C(micro_hash_ucr_pipe28_bF_buf0), .Y(_218_) );
INVX8 INVX8_34 ( .A(micro_hash_ucr_pipe29), .Y(_219_) );
INVX8 INVX8_35 ( .A(micro_hash_ucr_pipe28_bF_buf3), .Y(_220_) );
OAI21X1 OAI21X1_82 ( .A(_220__bF_buf4), .B(micro_hash_ucr_b_7_bF_buf0_), .C(_219_), .Y(_221_) );
AOI21X1 AOI21X1_36 ( .A(_218_), .B(_217_), .C(_221_), .Y(_222_) );
OAI21X1 OAI21X1_83 ( .A(_4200_), .B(_219_), .C(_4228__bF_buf2), .Y(_223_) );
OAI22X1 OAI22X1_7 ( .A(micro_hash_ucr_b_7_bF_buf3_), .B(_4228__bF_buf2), .C(_222_), .D(_223_), .Y(_224_) );
OAI21X1 OAI21X1_84 ( .A(_224_), .B(micro_hash_ucr_pipe31_bF_buf1), .C(_4227_), .Y(_225_) );
NAND2X1 NAND2X1_105 ( .A(_4226__bF_buf3), .B(_225_), .Y(_226_) );
OAI21X1 OAI21X1_85 ( .A(_4205_), .B(_4226__bF_buf3), .C(_226_), .Y(_227_) );
NAND2X1 NAND2X1_106 ( .A(micro_hash_ucr_pipe33_bF_buf3), .B(_4200_), .Y(_228_) );
OAI21X1 OAI21X1_86 ( .A(_227_), .B(micro_hash_ucr_pipe33_bF_buf3), .C(_228_), .Y(_229_) );
INVX8 INVX8_36 ( .A(micro_hash_ucr_pipe35), .Y(_230_) );
OAI21X1 OAI21X1_87 ( .A(_4225__bF_buf2), .B(micro_hash_ucr_b_7_bF_buf2_), .C(_230__bF_buf3), .Y(_231_) );
AOI21X1 AOI21X1_37 ( .A(_4225__bF_buf2), .B(_229_), .C(_231_), .Y(_232_) );
OAI21X1 OAI21X1_88 ( .A(_4200_), .B(_230__bF_buf3), .C(_4224__bF_buf0), .Y(_233_) );
OAI22X1 OAI22X1_8 ( .A(micro_hash_ucr_b_7_bF_buf1_), .B(_4224__bF_buf0), .C(_232_), .D(_233_), .Y(_234_) );
OAI21X1 OAI21X1_89 ( .A(_234_), .B(micro_hash_ucr_pipe37_bF_buf0), .C(_4223_), .Y(_235_) );
NAND2X1 NAND2X1_107 ( .A(micro_hash_ucr_pipe38_bF_buf1), .B(_4205_), .Y(_236_) );
OAI21X1 OAI21X1_90 ( .A(_235_), .B(micro_hash_ucr_pipe38_bF_buf1), .C(_236_), .Y(_237_) );
OAI21X1 OAI21X1_91 ( .A(_237_), .B(micro_hash_ucr_pipe39), .C(_4222_), .Y(_238_) );
NAND2X1 NAND2X1_108 ( .A(micro_hash_ucr_pipe40_bF_buf0), .B(_4205_), .Y(_239_) );
OAI21X1 OAI21X1_92 ( .A(_238_), .B(micro_hash_ucr_pipe40_bF_buf2), .C(_239_), .Y(_240_) );
OAI21X1 OAI21X1_93 ( .A(_240_), .B(micro_hash_ucr_pipe41_bF_buf1), .C(_4221_), .Y(_241_) );
INVX8 INVX8_37 ( .A(micro_hash_ucr_pipe43), .Y(_242_) );
OAI21X1 OAI21X1_94 ( .A(_4205_), .B(_4220__bF_buf3), .C(_242__bF_buf3), .Y(_243_) );
AOI21X1 AOI21X1_38 ( .A(_4220__bF_buf3), .B(_241_), .C(_243_), .Y(_244_) );
OAI21X1 OAI21X1_95 ( .A(_242__bF_buf3), .B(micro_hash_ucr_c_3_bF_buf0_), .C(_4219__bF_buf4), .Y(_245_) );
OAI22X1 OAI22X1_9 ( .A(_4205_), .B(_4219__bF_buf4), .C(_244_), .D(_245_), .Y(_246_) );
NAND2X1 NAND2X1_109 ( .A(micro_hash_ucr_pipe45), .B(_4200_), .Y(_247_) );
OAI21X1 OAI21X1_96 ( .A(_246_), .B(micro_hash_ucr_pipe45), .C(_247_), .Y(_248_) );
INVX8 INVX8_38 ( .A(micro_hash_ucr_pipe47), .Y(_249_) );
OAI21X1 OAI21X1_97 ( .A(_4218__bF_buf1), .B(micro_hash_ucr_b_7_bF_buf0_), .C(_249__bF_buf2), .Y(_250_) );
AOI21X1 AOI21X1_39 ( .A(_4218__bF_buf1), .B(_248_), .C(_250_), .Y(_251_) );
OAI21X1 OAI21X1_98 ( .A(_4200_), .B(_249__bF_buf0), .C(_4217__bF_buf0), .Y(_252_) );
OAI22X1 OAI22X1_10 ( .A(micro_hash_ucr_b_7_bF_buf3_), .B(_4217__bF_buf2), .C(_251_), .D(_252_), .Y(_253_) );
OAI21X1 OAI21X1_99 ( .A(_253_), .B(micro_hash_ucr_pipe49_bF_buf3), .C(_4216_), .Y(_254_) );
INVX8 INVX8_39 ( .A(micro_hash_ucr_pipe51), .Y(_255_) );
OAI21X1 OAI21X1_100 ( .A(_4205_), .B(_4215__bF_buf3), .C(_255__bF_buf3), .Y(_256_) );
AOI21X1 AOI21X1_40 ( .A(_4215__bF_buf3), .B(_254_), .C(_256_), .Y(_257_) );
OAI21X1 OAI21X1_101 ( .A(_255__bF_buf3), .B(micro_hash_ucr_c_3_bF_buf3_), .C(_4214__bF_buf1), .Y(_258_) );
OAI22X1 OAI22X1_11 ( .A(_4205_), .B(_4214__bF_buf1), .C(_257_), .D(_258_), .Y(_259_) );
NAND2X1 NAND2X1_110 ( .A(micro_hash_ucr_pipe53_bF_buf2), .B(_4200_), .Y(_260_) );
OAI21X1 OAI21X1_102 ( .A(_259_), .B(micro_hash_ucr_pipe53_bF_buf2), .C(_260_), .Y(_261_) );
OAI21X1 OAI21X1_103 ( .A(_261_), .B(micro_hash_ucr_pipe54_bF_buf2), .C(_4213_), .Y(_262_) );
NAND2X1 NAND2X1_111 ( .A(micro_hash_ucr_pipe55), .B(_4200_), .Y(_263_) );
OAI21X1 OAI21X1_104 ( .A(_262_), .B(micro_hash_ucr_pipe55), .C(_263_), .Y(_264_) );
AOI21X1 AOI21X1_41 ( .A(micro_hash_ucr_b_7_bF_buf2_), .B(micro_hash_ucr_pipe56_bF_buf3), .C(micro_hash_ucr_pipe57_bF_buf3), .Y(_265_) );
OAI21X1 OAI21X1_105 ( .A(_264_), .B(micro_hash_ucr_pipe56_bF_buf3), .C(_265_), .Y(_266_) );
OAI21X1 OAI21X1_106 ( .A(micro_hash_ucr_c_3_bF_buf2_), .B(_4212_), .C(_266_), .Y(_267_) );
AND2X2 AND2X2_15 ( .A(_267_), .B(_4211__bF_buf4), .Y(_268_) );
INVX8 INVX8_40 ( .A(micro_hash_ucr_pipe59), .Y(_269_) );
OAI21X1 OAI21X1_107 ( .A(_4211__bF_buf4), .B(micro_hash_ucr_b_7_bF_buf1_), .C(_269_), .Y(_270_) );
AOI21X1 AOI21X1_42 ( .A(micro_hash_ucr_c_3_bF_buf1_), .B(micro_hash_ucr_pipe59), .C(micro_hash_ucr_pipe60_bF_buf2), .Y(_271_) );
OAI21X1 OAI21X1_108 ( .A(_268_), .B(_270_), .C(_271_), .Y(_272_) );
OAI21X1 OAI21X1_109 ( .A(micro_hash_ucr_b_7_bF_buf0_), .B(_4210__bF_buf4), .C(_272_), .Y(_273_) );
AND2X2 AND2X2_16 ( .A(_273_), .B(_4208_), .Y(_274_) );
OAI21X1 OAI21X1_110 ( .A(_274_), .B(_4209_), .C(_4207__bF_buf3), .Y(_275_) );
NAND3X1 NAND3X1_53 ( .A(_4204_), .B(_4206_), .C(_275_), .Y(_276_) );
AOI21X1 AOI21X1_43 ( .A(_4203_), .B(_276_), .C(micro_hash_ucr_pipe64_bF_buf2), .Y(_277_) );
INVX8 INVX8_41 ( .A(micro_hash_ucr_pipe64_bF_buf0), .Y(_278_) );
INVX2 INVX2_15 ( .A(micro_hash_ucr_pipe65_bF_buf1), .Y(_279_) );
OAI21X1 OAI21X1_111 ( .A(_4205_), .B(_278__bF_buf2), .C(_279_), .Y(_280_) );
AOI21X1 AOI21X1_44 ( .A(micro_hash_ucr_pipe65_bF_buf3), .B(_4200_), .C(micro_hash_ucr_pipe66_bF_buf3), .Y(_281_) );
OAI21X1 OAI21X1_112 ( .A(_277_), .B(_280_), .C(_281_), .Y(_282_) );
NAND2X1 NAND2X1_112 ( .A(micro_hash_ucr_b_7_bF_buf3_), .B(micro_hash_ucr_pipe66_bF_buf3), .Y(_283_) );
AOI21X1 AOI21X1_45 ( .A(_283_), .B(_282_), .C(micro_hash_ucr_pipe67), .Y(_284_) );
OAI21X1 OAI21X1_113 ( .A(_284_), .B(_4202_), .C(_4199__bF_buf4), .Y(_285_) );
AOI21X1 AOI21X1_46 ( .A(micro_hash_ucr_b_7_bF_buf2_), .B(micro_hash_ucr_pipe68), .C(micro_hash_ucr_pipe69), .Y(_286_) );
INVX8 INVX8_42 ( .A(micro_hash_ucr_pipe69), .Y(_287_) );
INVX1 INVX1_76 ( .A(_0__bF_buf5), .Y(_288_) );
NAND2X1 NAND2X1_113 ( .A(reset_bF_buf1), .B(_288_), .Y(_289_) );
NOR2X1 NOR2X1_168 ( .A(comparador_next), .B(_289_), .Y(_131_) );
OAI21X1 OAI21X1_114 ( .A(micro_hash_ucr_c_3_bF_buf0_), .B(_287_), .C(_131__bF_buf10), .Y(_290_) );
AOI21X1 AOI21X1_47 ( .A(_286_), .B(_285_), .C(_290_), .Y(_127__7_) );
INVX1 INVX1_77 ( .A(micro_hash_ucr_k_0_), .Y(_291_) );
INVX8 INVX8_43 ( .A(_131__bF_buf11), .Y(_292_) );
NOR2X1 NOR2X1_169 ( .A(micro_hash_ucr_pipe40_bF_buf3), .B(micro_hash_ucr_pipe7), .Y(_293_) );
AOI21X1 AOI21X1_48 ( .A(_291_), .B(_293_), .C(_292__bF_buf1), .Y(_130__0_) );
NAND2X1 NAND2X1_114 ( .A(micro_hash_ucr_k_1_), .B(_293_), .Y(_294_) );
NOR2X1 NOR2X1_170 ( .A(_294_), .B(_292__bF_buf1), .Y(_130__1_) );
NAND2X1 NAND2X1_115 ( .A(micro_hash_ucr_k_2_), .B(_293_), .Y(_295_) );
NOR2X1 NOR2X1_171 ( .A(_295_), .B(_292__bF_buf6), .Y(_130__2_) );
INVX8 INVX8_44 ( .A(micro_hash_ucr_pipe40_bF_buf4), .Y(_296_) );
OAI21X1 OAI21X1_115 ( .A(micro_hash_ucr_pipe7), .B(micro_hash_ucr_k_3_), .C(_296__bF_buf4), .Y(_297_) );
NOR2X1 NOR2X1_172 ( .A(_297_), .B(_292__bF_buf5), .Y(_130__3_) );
OAI21X1 OAI21X1_116 ( .A(micro_hash_ucr_pipe7), .B(micro_hash_ucr_k_4_), .C(_296__bF_buf4), .Y(_298_) );
NOR2X1 NOR2X1_173 ( .A(_298_), .B(_292__bF_buf10), .Y(_130__4_) );
INVX2 INVX2_16 ( .A(micro_hash_ucr_k_5_), .Y(_299_) );
OAI21X1 OAI21X1_117 ( .A(_299_), .B(micro_hash_ucr_pipe7), .C(_296__bF_buf4), .Y(_300_) );
AND2X2 AND2X2_17 ( .A(_131__bF_buf10), .B(_300_), .Y(_130__5_) );
NAND2X1 NAND2X1_116 ( .A(micro_hash_ucr_k_6_), .B(_293_), .Y(_301_) );
NOR2X1 NOR2X1_174 ( .A(_301_), .B(_292__bF_buf10), .Y(_130__6_) );
INVX1 INVX1_78 ( .A(micro_hash_ucr_k_7_), .Y(_302_) );
AOI21X1 AOI21X1_49 ( .A(_302_), .B(_293_), .C(_292__bF_buf10), .Y(_130__7_) );
NOR2X1 NOR2X1_175 ( .A(micro_hash_ucr_b_0_bF_buf3_), .B(micro_hash_ucr_a_0_bF_buf3_), .Y(_303_) );
INVX8 INVX8_45 ( .A(micro_hash_ucr_pipe49_bF_buf2), .Y(_304_) );
NOR2X1 NOR2X1_176 ( .A(micro_hash_ucr_pipe53_bF_buf2), .B(micro_hash_ucr_pipe55), .Y(_305_) );
NAND3X1 NAND3X1_54 ( .A(_304_), .B(_255__bF_buf1), .C(_305_), .Y(_306_) );
NOR2X1 NOR2X1_177 ( .A(micro_hash_ucr_pipe65_bF_buf3), .B(micro_hash_ucr_pipe67), .Y(_307_) );
NOR2X1 NOR2X1_178 ( .A(micro_hash_ucr_pipe61_bF_buf1), .B(micro_hash_ucr_pipe63_bF_buf2), .Y(_308_) );
INVX1 INVX1_79 ( .A(_308_), .Y(_309_) );
NOR2X1 NOR2X1_179 ( .A(micro_hash_ucr_pipe57_bF_buf3), .B(micro_hash_ucr_pipe59), .Y(_310_) );
INVX1 INVX1_80 ( .A(_310_), .Y(_311_) );
NOR2X1 NOR2X1_180 ( .A(_309_), .B(_311_), .Y(_312_) );
NAND2X1 NAND2X1_117 ( .A(_307_), .B(_312_), .Y(_313_) );
NOR2X1 NOR2X1_181 ( .A(_306_), .B(_313_), .Y(_314_) );
OAI21X1 OAI21X1_118 ( .A(_314_), .B(_303_), .C(_287_), .Y(_315_) );
INVX1 INVX1_81 ( .A(micro_hash_ucr_x_0_), .Y(_316_) );
INVX8 INVX8_46 ( .A(micro_hash_ucr_pipe31_bF_buf0), .Y(_317_) );
INVX8 INVX8_47 ( .A(micro_hash_ucr_pipe33_bF_buf0), .Y(_318_) );
NOR2X1 NOR2X1_182 ( .A(micro_hash_ucr_pipe27_bF_buf3), .B(micro_hash_ucr_pipe29), .Y(_319_) );
AND2X2 AND2X2_18 ( .A(_4267_), .B(_319_), .Y(_320_) );
NAND3X1 NAND3X1_55 ( .A(_317__bF_buf1), .B(_318_), .C(_320_), .Y(_321_) );
NOR2X1 NOR2X1_183 ( .A(micro_hash_ucr_pipe11), .B(micro_hash_ucr_pipe17), .Y(_322_) );
AND2X2 AND2X2_19 ( .A(_4271_), .B(_322_), .Y(_323_) );
NOR2X1 NOR2X1_184 ( .A(micro_hash_ucr_pipe23), .B(micro_hash_ucr_pipe25_bF_buf3), .Y(_324_) );
AND2X2 AND2X2_20 ( .A(_4270_), .B(_230__bF_buf3), .Y(_325_) );
NAND3X1 NAND3X1_56 ( .A(_324_), .B(_325_), .C(_323_), .Y(_326_) );
NOR2X1 NOR2X1_185 ( .A(_326_), .B(_321_), .Y(_327_) );
AND2X2 AND2X2_21 ( .A(_327_), .B(_316_), .Y(_328_) );
NOR2X1 NOR2X1_186 ( .A(micro_hash_ucr_pipe37_bF_buf0), .B(micro_hash_ucr_pipe39), .Y(_329_) );
INVX8 INVX8_48 ( .A(micro_hash_ucr_b_0_bF_buf2_), .Y(_330_) );
INVX8 INVX8_49 ( .A(micro_hash_ucr_a_0_bF_buf2_), .Y(_331_) );
NOR2X1 NOR2X1_187 ( .A(_330_), .B(_331_), .Y(_332_) );
NOR2X1 NOR2X1_188 ( .A(_303_), .B(_332_), .Y(_333_) );
OAI21X1 OAI21X1_119 ( .A(_327_), .B(_333_), .C(_329_), .Y(_334_) );
INVX1 INVX1_82 ( .A(_329_), .Y(_335_) );
INVX8 INVX8_50 ( .A(micro_hash_ucr_pipe45), .Y(_336_) );
NOR2X1 NOR2X1_189 ( .A(micro_hash_ucr_pipe41_bF_buf1), .B(micro_hash_ucr_pipe43), .Y(_337_) );
NAND3X1 NAND3X1_57 ( .A(_336_), .B(_249__bF_buf2), .C(_337_), .Y(_338_) );
AOI21X1 AOI21X1_50 ( .A(_335_), .B(_333_), .C(_338_), .Y(_339_) );
OAI21X1 OAI21X1_120 ( .A(_328_), .B(_334_), .C(_339_), .Y(_340_) );
INVX1 INVX1_83 ( .A(_314_), .Y(_341_) );
AOI21X1 AOI21X1_51 ( .A(_303_), .B(_338_), .C(_341_), .Y(_342_) );
AOI21X1 AOI21X1_52 ( .A(_342_), .B(_340_), .C(_315_), .Y(_343_) );
NOR2X1 NOR2X1_190 ( .A(micro_hash_ucr_pipe69), .B(_292__bF_buf5), .Y(_344_) );
INVX4 INVX4_7 ( .A(_344_), .Y(_345_) );
OAI21X1 OAI21X1_121 ( .A(micro_hash_ucr_b_0_bF_buf1_), .B(micro_hash_ucr_a_0_bF_buf1_), .C(_131__bF_buf10), .Y(_346_) );
AOI21X1 AOI21X1_53 ( .A(_345_), .B(_346_), .C(_343_), .Y(_204__0_) );
NAND2X1 NAND2X1_118 ( .A(_317__bF_buf1), .B(_318_), .Y(_347_) );
NAND2X1 NAND2X1_119 ( .A(_323_), .B(_4267_), .Y(_348_) );
NOR2X1 NOR2X1_191 ( .A(_347_), .B(_348_), .Y(_349_) );
NAND2X1 NAND2X1_120 ( .A(_4234__bF_buf1), .B(_4270_), .Y(_350_) );
NOR2X1 NOR2X1_192 ( .A(micro_hash_ucr_pipe35), .B(micro_hash_ucr_pipe37_bF_buf0), .Y(_351_) );
NOR2X1 NOR2X1_193 ( .A(micro_hash_ucr_pipe25_bF_buf3), .B(micro_hash_ucr_pipe39), .Y(_352_) );
NAND3X1 NAND3X1_58 ( .A(_319_), .B(_351_), .C(_352_), .Y(_353_) );
NOR2X1 NOR2X1_194 ( .A(_350_), .B(_353_), .Y(_354_) );
NAND2X1 NAND2X1_121 ( .A(_354_), .B(_349_), .Y(_355_) );
INVX4 INVX4_8 ( .A(_355_), .Y(_356_) );
AOI21X1 AOI21X1_54 ( .A(micro_hash_ucr_b_1_bF_buf3_), .B(micro_hash_ucr_a_1_), .C(_356_), .Y(_357_) );
NOR2X1 NOR2X1_195 ( .A(_306_), .B(_338_), .Y(_358_) );
NAND2X1 NAND2X1_122 ( .A(_287_), .B(_307_), .Y(_359_) );
NOR2X1 NOR2X1_196 ( .A(_309_), .B(_359_), .Y(_360_) );
INVX1 INVX1_84 ( .A(_360_), .Y(_361_) );
NOR2X1 NOR2X1_197 ( .A(_311_), .B(_361_), .Y(_362_) );
NAND2X1 NAND2X1_123 ( .A(_358_), .B(_362_), .Y(_363_) );
OAI22X1 OAI22X1_12 ( .A(micro_hash_ucr_b_1_bF_buf2_), .B(micro_hash_ucr_a_1_), .C(_357_), .D(_363_), .Y(_364_) );
INVX2 INVX2_17 ( .A(_363_), .Y(_365_) );
NAND3X1 NAND3X1_59 ( .A(micro_hash_ucr_x_1_), .B(_356_), .C(_365_), .Y(_366_) );
AOI21X1 AOI21X1_55 ( .A(_366_), .B(_364_), .C(_292__bF_buf5), .Y(_204__1_) );
AOI21X1 AOI21X1_56 ( .A(micro_hash_ucr_b_2_bF_buf3_), .B(micro_hash_ucr_a_2_bF_buf4_), .C(_356_), .Y(_367_) );
OAI22X1 OAI22X1_13 ( .A(micro_hash_ucr_b_2_bF_buf2_), .B(micro_hash_ucr_a_2_bF_buf3_), .C(_367_), .D(_363_), .Y(_368_) );
NAND3X1 NAND3X1_60 ( .A(micro_hash_ucr_x_2_), .B(_356_), .C(_365_), .Y(_369_) );
AOI21X1 AOI21X1_57 ( .A(_369_), .B(_368_), .C(_292__bF_buf5), .Y(_204__2_) );
AOI21X1 AOI21X1_58 ( .A(micro_hash_ucr_b_3_bF_buf3_), .B(micro_hash_ucr_a_3_bF_buf3_), .C(_356_), .Y(_370_) );
OAI22X1 OAI22X1_14 ( .A(micro_hash_ucr_b_3_bF_buf2_), .B(micro_hash_ucr_a_3_bF_buf2_), .C(_370_), .D(_363_), .Y(_371_) );
NOR2X1 NOR2X1_198 ( .A(micro_hash_ucr_pipe33_bF_buf3), .B(micro_hash_ucr_pipe35), .Y(_372_) );
AND2X2 AND2X2_22 ( .A(_329_), .B(_372_), .Y(_373_) );
NOR2X1 NOR2X1_199 ( .A(micro_hash_ucr_pipe17), .B(micro_hash_ucr_pipe31_bF_buf3), .Y(_374_) );
NAND3X1 NAND3X1_61 ( .A(_4271_), .B(_374_), .C(_373_), .Y(_375_) );
NAND3X1 NAND3X1_62 ( .A(_4234__bF_buf1), .B(_4270_), .C(_320_), .Y(_376_) );
NOR2X1 NOR2X1_200 ( .A(_375_), .B(_376_), .Y(_377_) );
NOR2X1 NOR2X1_201 ( .A(micro_hash_ucr_pipe11), .B(micro_hash_ucr_pipe25_bF_buf3), .Y(_378_) );
NAND3X1 NAND3X1_63 ( .A(_287_), .B(micro_hash_ucr_x_3_), .C(_378_), .Y(_379_) );
NOR2X1 NOR2X1_202 ( .A(_379_), .B(_313_), .Y(_380_) );
NAND3X1 NAND3X1_64 ( .A(_358_), .B(_380_), .C(_377_), .Y(_381_) );
AOI21X1 AOI21X1_59 ( .A(_381_), .B(_371_), .C(_292__bF_buf7), .Y(_204__3_) );
AOI21X1 AOI21X1_60 ( .A(micro_hash_ucr_b_4_), .B(micro_hash_ucr_a_4_bF_buf3_), .C(_356_), .Y(_382_) );
OAI22X1 OAI22X1_15 ( .A(micro_hash_ucr_b_4_), .B(micro_hash_ucr_a_4_bF_buf2_), .C(_382_), .D(_363_), .Y(_383_) );
NAND2X1 NAND2X1_124 ( .A(micro_hash_ucr_x_4_), .B(_287_), .Y(_384_) );
NOR2X1 NOR2X1_203 ( .A(_384_), .B(_313_), .Y(_385_) );
NAND3X1 NAND3X1_65 ( .A(_358_), .B(_385_), .C(_356_), .Y(_386_) );
AOI21X1 AOI21X1_61 ( .A(_386_), .B(_383_), .C(_292__bF_buf5), .Y(_204__4_) );
XNOR2X1 XNOR2X1_7 ( .A(micro_hash_ucr_b_5_bF_buf3_), .B(micro_hash_ucr_a_5_bF_buf3_), .Y(_387_) );
OAI21X1 OAI21X1_122 ( .A(_363_), .B(_355_), .C(_387_), .Y(_388_) );
INVX8 INVX8_51 ( .A(micro_hash_ucr_pipe25_bF_buf1), .Y(_389_) );
NAND3X1 NAND3X1_66 ( .A(_389__bF_buf0), .B(_317__bF_buf1), .C(_319_), .Y(_390_) );
NOR2X1 NOR2X1_204 ( .A(_335_), .B(_390_), .Y(_391_) );
INVX2 INVX2_18 ( .A(micro_hash_ucr_x_5_), .Y(_392_) );
NAND2X1 NAND2X1_125 ( .A(_4234__bF_buf1), .B(_392_), .Y(_393_) );
NAND3X1 NAND3X1_67 ( .A(_4270_), .B(_372_), .C(_323_), .Y(_394_) );
NOR2X1 NOR2X1_205 ( .A(_393_), .B(_394_), .Y(_395_) );
NAND2X1 NAND2X1_126 ( .A(_391_), .B(_395_), .Y(_396_) );
OAI21X1 OAI21X1_123 ( .A(_4266_), .B(_396_), .C(_388_), .Y(_397_) );
OAI21X1 OAI21X1_124 ( .A(micro_hash_ucr_b_5_bF_buf2_), .B(micro_hash_ucr_a_5_bF_buf2_), .C(_363_), .Y(_398_) );
AOI21X1 AOI21X1_62 ( .A(_398_), .B(_397_), .C(_292__bF_buf5), .Y(_204__5_) );
INVX8 INVX8_52 ( .A(micro_hash_ucr_b_6_bF_buf3_), .Y(_399_) );
INVX4 INVX4_9 ( .A(micro_hash_ucr_a_6_bF_buf3_), .Y(_400_) );
NAND2X1 NAND2X1_127 ( .A(_399__bF_buf2), .B(_400_), .Y(_401_) );
AOI21X1 AOI21X1_63 ( .A(micro_hash_ucr_b_6_bF_buf2_), .B(micro_hash_ucr_a_6_bF_buf2_), .C(_356_), .Y(_402_) );
INVX1 INVX1_85 ( .A(_313_), .Y(_403_) );
NAND2X1 NAND2X1_128 ( .A(_358_), .B(_403_), .Y(_404_) );
OAI21X1 OAI21X1_125 ( .A(_402_), .B(_404_), .C(_401_), .Y(_405_) );
INVX1 INVX1_86 ( .A(_358_), .Y(_406_) );
NAND2X1 NAND2X1_129 ( .A(micro_hash_ucr_x_6_), .B(_403_), .Y(_407_) );
NOR2X1 NOR2X1_206 ( .A(_406_), .B(_407_), .Y(_408_) );
AOI21X1 AOI21X1_64 ( .A(_356_), .B(_408_), .C(micro_hash_ucr_pipe69), .Y(_409_) );
OAI21X1 OAI21X1_126 ( .A(_287_), .B(_401_), .C(_131__bF_buf10), .Y(_410_) );
AOI21X1 AOI21X1_65 ( .A(_409_), .B(_405_), .C(_410_), .Y(_204__6_) );
NOR2X1 NOR2X1_207 ( .A(micro_hash_ucr_b_7_bF_buf1_), .B(micro_hash_ucr_a_7_bF_buf3_), .Y(_411_) );
AOI21X1 AOI21X1_66 ( .A(_349_), .B(_365_), .C(_411_), .Y(_412_) );
INVX1 INVX1_87 ( .A(micro_hash_ucr_x_7_), .Y(_413_) );
NAND2X1 NAND2X1_130 ( .A(_413_), .B(_354_), .Y(_414_) );
NOR2X1 NOR2X1_208 ( .A(_414_), .B(_412_), .Y(_415_) );
NAND3X1 NAND3X1_68 ( .A(micro_hash_ucr_b_7_bF_buf0_), .B(micro_hash_ucr_a_7_bF_buf2_), .C(_312_), .Y(_416_) );
NOR2X1 NOR2X1_209 ( .A(_359_), .B(_416_), .Y(_417_) );
AOI21X1 AOI21X1_67 ( .A(_358_), .B(_417_), .C(_411_), .Y(_418_) );
AOI21X1 AOI21X1_68 ( .A(_411_), .B(_363_), .C(_292__bF_buf5), .Y(_419_) );
OAI21X1 OAI21X1_127 ( .A(_356_), .B(_418_), .C(_419_), .Y(_420_) );
NOR2X1 NOR2X1_210 ( .A(_420_), .B(_415_), .Y(_204__7_) );
INVX1 INVX1_88 ( .A(micro_hash_ucr_Wx_200_), .Y(_421_) );
NOR2X1 NOR2X1_211 ( .A(micro_hash_ucr_k_0_), .B(micro_hash_ucr_x_0_), .Y(_422_) );
NOR2X1 NOR2X1_212 ( .A(_291_), .B(_316_), .Y(_423_) );
OAI21X1 OAI21X1_128 ( .A(_423_), .B(_422_), .C(_421_), .Y(_424_) );
NOR2X1 NOR2X1_213 ( .A(_422_), .B(_423_), .Y(_425_) );
INVX8 INVX8_53 ( .A(_425__bF_buf5), .Y(_426_) );
NOR2X1 NOR2X1_214 ( .A(_421_), .B(_426__bF_buf0), .Y(_427_) );
INVX1 INVX1_89 ( .A(_427_), .Y(_428_) );
NAND2X1 NAND2X1_131 ( .A(_424_), .B(_428_), .Y(_429_) );
NOR2X1 NOR2X1_215 ( .A(micro_hash_ucr_Wx_24_), .B(_425__bF_buf1), .Y(_430_) );
INVX2 INVX2_19 ( .A(micro_hash_ucr_Wx_24_), .Y(_431_) );
NOR2X1 NOR2X1_216 ( .A(_431_), .B(_426__bF_buf3), .Y(_432_) );
OAI21X1 OAI21X1_129 ( .A(_432_), .B(_430_), .C(micro_hash_ucr_pipe14), .Y(_433_) );
NOR2X1 NOR2X1_217 ( .A(micro_hash_ucr_Wx_8_), .B(_425__bF_buf1), .Y(_434_) );
NAND2X1 NAND2X1_132 ( .A(micro_hash_ucr_Wx_8_), .B(_425__bF_buf1), .Y(_435_) );
INVX2 INVX2_20 ( .A(_435_), .Y(_436_) );
OAI21X1 OAI21X1_130 ( .A(_436_), .B(_434_), .C(micro_hash_ucr_pipe10), .Y(_437_) );
INVX4 INVX4_10 ( .A(micro_hash_ucr_pipe8), .Y(_438_) );
NAND2X1 NAND2X1_133 ( .A(micro_hash_ucr_Wx_0_), .B(_425__bF_buf1), .Y(_439_) );
INVX2 INVX2_21 ( .A(_439_), .Y(_440_) );
NOR2X1 NOR2X1_218 ( .A(_438_), .B(_440_), .Y(_441_) );
OAI21X1 OAI21X1_131 ( .A(micro_hash_ucr_Wx_0_), .B(_425__bF_buf1), .C(_441_), .Y(_442_) );
INVX2 INVX2_22 ( .A(H_16_), .Y(_443_) );
NAND2X1 NAND2X1_134 ( .A(micro_hash_ucr_pipe6), .B(_443_), .Y(_444_) );
OAI21X1 OAI21X1_132 ( .A(micro_hash_ucr_c_0_bF_buf3_), .B(micro_hash_ucr_pipe6), .C(_444_), .Y(_445_) );
OAI21X1 OAI21X1_133 ( .A(micro_hash_ucr_pipe8), .B(_445_), .C(_442_), .Y(_446_) );
OAI21X1 OAI21X1_134 ( .A(_446_), .B(micro_hash_ucr_pipe10), .C(_437_), .Y(_447_) );
NAND2X1 NAND2X1_135 ( .A(micro_hash_ucr_Wx_16_), .B(_425__bF_buf1), .Y(_448_) );
INVX2 INVX2_23 ( .A(micro_hash_ucr_Wx_16_), .Y(_449_) );
OAI21X1 OAI21X1_135 ( .A(_423_), .B(_422_), .C(_449_), .Y(_450_) );
NAND3X1 NAND3X1_69 ( .A(micro_hash_ucr_pipe12_bF_buf2), .B(_450_), .C(_448_), .Y(_451_) );
OAI21X1 OAI21X1_136 ( .A(_447_), .B(micro_hash_ucr_pipe12_bF_buf2), .C(_451_), .Y(_452_) );
OAI21X1 OAI21X1_137 ( .A(_452_), .B(micro_hash_ucr_pipe14), .C(_433_), .Y(_453_) );
NAND2X1 NAND2X1_136 ( .A(_4239__bF_buf2), .B(_453_), .Y(_454_) );
INVX2 INVX2_24 ( .A(micro_hash_ucr_Wx_32_), .Y(_455_) );
NOR2X1 NOR2X1_219 ( .A(_455_), .B(_426__bF_buf3), .Y(_456_) );
NOR2X1 NOR2X1_220 ( .A(micro_hash_ucr_Wx_32_), .B(_425__bF_buf1), .Y(_457_) );
OAI21X1 OAI21X1_138 ( .A(_456_), .B(_457_), .C(micro_hash_ucr_pipe16), .Y(_458_) );
NAND2X1 NAND2X1_137 ( .A(_458_), .B(_454_), .Y(_459_) );
NOR2X1 NOR2X1_221 ( .A(micro_hash_ucr_pipe18_bF_buf3), .B(_459_), .Y(_460_) );
INVX2 INVX2_25 ( .A(micro_hash_ucr_Wx_40_), .Y(_461_) );
NOR2X1 NOR2X1_222 ( .A(_461_), .B(_426__bF_buf3), .Y(_462_) );
OAI21X1 OAI21X1_139 ( .A(_425__bF_buf0), .B(micro_hash_ucr_Wx_40_), .C(micro_hash_ucr_pipe18_bF_buf3), .Y(_463_) );
OAI21X1 OAI21X1_140 ( .A(_462_), .B(_463_), .C(_4237__bF_buf1), .Y(_464_) );
OR2X2 OR2X2_11 ( .A(_460_), .B(_464_), .Y(_465_) );
NOR2X1 NOR2X1_223 ( .A(micro_hash_ucr_Wx_48_), .B(_425__bF_buf0), .Y(_466_) );
INVX2 INVX2_26 ( .A(micro_hash_ucr_Wx_48_), .Y(_467_) );
NOR2X1 NOR2X1_224 ( .A(_467_), .B(_426__bF_buf3), .Y(_468_) );
OAI21X1 OAI21X1_141 ( .A(_468_), .B(_466_), .C(micro_hash_ucr_pipe20_bF_buf1), .Y(_469_) );
AND2X2 AND2X2_23 ( .A(_465_), .B(_469_), .Y(_470_) );
INVX2 INVX2_27 ( .A(micro_hash_ucr_Wx_56_), .Y(_471_) );
NOR2X1 NOR2X1_225 ( .A(_471_), .B(_426__bF_buf3), .Y(_472_) );
NOR2X1 NOR2X1_226 ( .A(micro_hash_ucr_Wx_56_), .B(_425__bF_buf0), .Y(_473_) );
OAI21X1 OAI21X1_142 ( .A(_472_), .B(_473_), .C(micro_hash_ucr_pipe22_bF_buf1), .Y(_474_) );
OAI21X1 OAI21X1_143 ( .A(_470_), .B(micro_hash_ucr_pipe22_bF_buf1), .C(_474_), .Y(_475_) );
INVX2 INVX2_28 ( .A(micro_hash_ucr_Wx_64_), .Y(_476_) );
OAI21X1 OAI21X1_144 ( .A(_423_), .B(_422_), .C(_476_), .Y(_477_) );
NOR2X1 NOR2X1_227 ( .A(_476_), .B(_426__bF_buf2), .Y(_478_) );
NOR2X1 NOR2X1_228 ( .A(_4233__bF_buf0), .B(_478_), .Y(_479_) );
AOI21X1 AOI21X1_69 ( .A(_477_), .B(_479_), .C(micro_hash_ucr_pipe26_bF_buf0), .Y(_480_) );
OAI21X1 OAI21X1_145 ( .A(_475_), .B(micro_hash_ucr_pipe24_bF_buf1), .C(_480_), .Y(_481_) );
NOR2X1 NOR2X1_229 ( .A(micro_hash_ucr_Wx_72_), .B(_425__bF_buf0), .Y(_482_) );
INVX2 INVX2_29 ( .A(micro_hash_ucr_Wx_72_), .Y(_483_) );
NOR2X1 NOR2X1_230 ( .A(_483_), .B(_426__bF_buf2), .Y(_484_) );
OAI21X1 OAI21X1_146 ( .A(_484_), .B(_482_), .C(micro_hash_ucr_pipe26_bF_buf2), .Y(_485_) );
NAND3X1 NAND3X1_70 ( .A(_220__bF_buf3), .B(_485_), .C(_481_), .Y(_486_) );
NAND2X1 NAND2X1_138 ( .A(micro_hash_ucr_Wx_80_), .B(_425__bF_buf0), .Y(_487_) );
INVX2 INVX2_30 ( .A(micro_hash_ucr_Wx_80_), .Y(_488_) );
OAI21X1 OAI21X1_147 ( .A(_423_), .B(_422_), .C(_488_), .Y(_489_) );
NAND2X1 NAND2X1_139 ( .A(_489_), .B(_487_), .Y(_490_) );
OAI21X1 OAI21X1_148 ( .A(_220__bF_buf0), .B(_490_), .C(_486_), .Y(_491_) );
NOR2X1 NOR2X1_231 ( .A(micro_hash_ucr_Wx_88_), .B(_425__bF_buf0), .Y(_492_) );
INVX2 INVX2_31 ( .A(micro_hash_ucr_Wx_88_), .Y(_493_) );
NOR2X1 NOR2X1_232 ( .A(_493_), .B(_426__bF_buf2), .Y(_494_) );
OAI21X1 OAI21X1_149 ( .A(_494_), .B(_492_), .C(micro_hash_ucr_pipe30_bF_buf1), .Y(_495_) );
OAI21X1 OAI21X1_150 ( .A(_491_), .B(micro_hash_ucr_pipe30_bF_buf1), .C(_495_), .Y(_496_) );
NAND2X1 NAND2X1_140 ( .A(micro_hash_ucr_Wx_96_), .B(_425__bF_buf0), .Y(_497_) );
INVX2 INVX2_32 ( .A(micro_hash_ucr_Wx_96_), .Y(_498_) );
AOI21X1 AOI21X1_70 ( .A(_498_), .B(_426__bF_buf2), .C(_4226__bF_buf0), .Y(_499_) );
AOI21X1 AOI21X1_71 ( .A(_497_), .B(_499_), .C(micro_hash_ucr_pipe34_bF_buf2), .Y(_500_) );
OAI21X1 OAI21X1_151 ( .A(_496_), .B(micro_hash_ucr_pipe32_bF_buf3), .C(_500_), .Y(_501_) );
NOR2X1 NOR2X1_233 ( .A(micro_hash_ucr_Wx_104_), .B(_425__bF_buf5), .Y(_502_) );
INVX2 INVX2_33 ( .A(micro_hash_ucr_Wx_104_), .Y(_503_) );
NOR2X1 NOR2X1_234 ( .A(_503_), .B(_426__bF_buf0), .Y(_504_) );
OAI21X1 OAI21X1_152 ( .A(_504_), .B(_502_), .C(micro_hash_ucr_pipe34_bF_buf2), .Y(_505_) );
NAND3X1 NAND3X1_71 ( .A(_4224__bF_buf3), .B(_505_), .C(_501_), .Y(_506_) );
INVX2 INVX2_34 ( .A(micro_hash_ucr_Wx_112_), .Y(_507_) );
NOR2X1 NOR2X1_235 ( .A(_507_), .B(_426__bF_buf0), .Y(_508_) );
OAI21X1 OAI21X1_153 ( .A(_425__bF_buf5), .B(micro_hash_ucr_Wx_112_), .C(micro_hash_ucr_pipe36_bF_buf1), .Y(_509_) );
OAI21X1 OAI21X1_154 ( .A(_508_), .B(_509_), .C(_506_), .Y(_510_) );
NOR2X1 NOR2X1_236 ( .A(micro_hash_ucr_Wx_120_), .B(_425__bF_buf5), .Y(_511_) );
INVX2 INVX2_35 ( .A(micro_hash_ucr_Wx_120_), .Y(_512_) );
NOR2X1 NOR2X1_237 ( .A(_512_), .B(_426__bF_buf0), .Y(_513_) );
OAI21X1 OAI21X1_155 ( .A(_513_), .B(_511_), .C(micro_hash_ucr_pipe38_bF_buf3), .Y(_514_) );
OAI21X1 OAI21X1_156 ( .A(_510_), .B(micro_hash_ucr_pipe38_bF_buf3), .C(_514_), .Y(_515_) );
INVX2 INVX2_36 ( .A(micro_hash_ucr_Wx_128_), .Y(_516_) );
NOR2X1 NOR2X1_238 ( .A(_516_), .B(_426__bF_buf0), .Y(_517_) );
NOR2X1 NOR2X1_239 ( .A(_296__bF_buf2), .B(_517_), .Y(_518_) );
OAI21X1 OAI21X1_157 ( .A(micro_hash_ucr_Wx_128_), .B(_425__bF_buf5), .C(_518_), .Y(_519_) );
AND2X2 AND2X2_24 ( .A(_519_), .B(_4220__bF_buf4), .Y(_520_) );
OAI21X1 OAI21X1_158 ( .A(_515_), .B(micro_hash_ucr_pipe40_bF_buf4), .C(_520_), .Y(_521_) );
NOR2X1 NOR2X1_240 ( .A(micro_hash_ucr_Wx_136_), .B(_425__bF_buf5), .Y(_522_) );
INVX2 INVX2_37 ( .A(micro_hash_ucr_Wx_136_), .Y(_523_) );
NOR2X1 NOR2X1_241 ( .A(_523_), .B(_426__bF_buf1), .Y(_524_) );
OAI21X1 OAI21X1_159 ( .A(_524_), .B(_522_), .C(micro_hash_ucr_pipe42_bF_buf1), .Y(_525_) );
NAND3X1 NAND3X1_72 ( .A(_4219__bF_buf1), .B(_525_), .C(_521_), .Y(_526_) );
AND2X2 AND2X2_25 ( .A(_425__bF_buf4), .B(micro_hash_ucr_Wx_144_), .Y(_527_) );
OAI21X1 OAI21X1_160 ( .A(_425__bF_buf4), .B(micro_hash_ucr_Wx_144_), .C(micro_hash_ucr_pipe44_bF_buf1), .Y(_528_) );
OAI21X1 OAI21X1_161 ( .A(_527_), .B(_528_), .C(_526_), .Y(_529_) );
NOR2X1 NOR2X1_242 ( .A(micro_hash_ucr_Wx_152_), .B(_425__bF_buf4), .Y(_530_) );
AND2X2 AND2X2_26 ( .A(_425__bF_buf4), .B(micro_hash_ucr_Wx_152_), .Y(_531_) );
OAI21X1 OAI21X1_162 ( .A(_531_), .B(_530_), .C(micro_hash_ucr_pipe46_bF_buf0), .Y(_532_) );
OAI21X1 OAI21X1_163 ( .A(_529_), .B(micro_hash_ucr_pipe46_bF_buf0), .C(_532_), .Y(_533_) );
OAI21X1 OAI21X1_164 ( .A(_425__bF_buf3), .B(micro_hash_ucr_Wx_160_), .C(micro_hash_ucr_pipe48_bF_buf3), .Y(_534_) );
AOI21X1 AOI21X1_72 ( .A(micro_hash_ucr_Wx_160_), .B(_425__bF_buf3), .C(_534_), .Y(_535_) );
NOR2X1 NOR2X1_243 ( .A(micro_hash_ucr_pipe50_bF_buf2), .B(_535_), .Y(_536_) );
OAI21X1 OAI21X1_165 ( .A(_533_), .B(micro_hash_ucr_pipe48_bF_buf1), .C(_536_), .Y(_537_) );
NOR2X1 NOR2X1_244 ( .A(micro_hash_ucr_Wx_168_), .B(_425__bF_buf2), .Y(_538_) );
AND2X2 AND2X2_27 ( .A(_425__bF_buf2), .B(micro_hash_ucr_Wx_168_), .Y(_539_) );
OAI21X1 OAI21X1_166 ( .A(_539_), .B(_538_), .C(micro_hash_ucr_pipe50_bF_buf0), .Y(_540_) );
NAND2X1 NAND2X1_141 ( .A(_540_), .B(_537_), .Y(_541_) );
AND2X2 AND2X2_28 ( .A(_425__bF_buf4), .B(micro_hash_ucr_Wx_176_), .Y(_542_) );
OAI21X1 OAI21X1_167 ( .A(_425__bF_buf3), .B(micro_hash_ucr_Wx_176_), .C(micro_hash_ucr_pipe52_bF_buf1), .Y(_543_) );
OAI22X1 OAI22X1_16 ( .A(_542_), .B(_543_), .C(_541_), .D(micro_hash_ucr_pipe52_bF_buf3), .Y(_544_) );
NOR2X1 NOR2X1_245 ( .A(micro_hash_ucr_Wx_184_), .B(_425__bF_buf4), .Y(_545_) );
AND2X2 AND2X2_29 ( .A(_425__bF_buf4), .B(micro_hash_ucr_Wx_184_), .Y(_546_) );
OAI21X1 OAI21X1_168 ( .A(_546_), .B(_545_), .C(micro_hash_ucr_pipe54_bF_buf0), .Y(_547_) );
OAI21X1 OAI21X1_169 ( .A(_544_), .B(micro_hash_ucr_pipe54_bF_buf0), .C(_547_), .Y(_548_) );
NOR2X1 NOR2X1_246 ( .A(micro_hash_ucr_pipe56_bF_buf1), .B(_548_), .Y(_549_) );
AND2X2 AND2X2_30 ( .A(_425__bF_buf5), .B(micro_hash_ucr_Wx_192_), .Y(_550_) );
OAI21X1 OAI21X1_170 ( .A(_425__bF_buf5), .B(micro_hash_ucr_Wx_192_), .C(micro_hash_ucr_pipe56_bF_buf1), .Y(_551_) );
NOR2X1 NOR2X1_247 ( .A(_551_), .B(_550_), .Y(_552_) );
OAI21X1 OAI21X1_171 ( .A(_549_), .B(_552_), .C(_4211__bF_buf2), .Y(_553_) );
OAI21X1 OAI21X1_172 ( .A(_4211__bF_buf2), .B(_429_), .C(_553_), .Y(_554_) );
AND2X2 AND2X2_31 ( .A(_425__bF_buf3), .B(micro_hash_ucr_Wx_208_), .Y(_555_) );
OAI21X1 OAI21X1_173 ( .A(_425__bF_buf3), .B(micro_hash_ucr_Wx_208_), .C(micro_hash_ucr_pipe60_bF_buf0), .Y(_556_) );
OAI21X1 OAI21X1_174 ( .A(_555_), .B(_556_), .C(_4207__bF_buf0), .Y(_557_) );
AOI21X1 AOI21X1_73 ( .A(_4210__bF_buf2), .B(_554_), .C(_557_), .Y(_558_) );
NOR2X1 NOR2X1_248 ( .A(micro_hash_ucr_Wx_216_), .B(_425__bF_buf3), .Y(_559_) );
NAND2X1 NAND2X1_142 ( .A(micro_hash_ucr_Wx_216_), .B(_425__bF_buf3), .Y(_560_) );
INVX2 INVX2_38 ( .A(_560_), .Y(_561_) );
OAI21X1 OAI21X1_175 ( .A(_561_), .B(_559_), .C(micro_hash_ucr_pipe62_bF_buf1), .Y(_562_) );
NAND2X1 NAND2X1_143 ( .A(_278__bF_buf3), .B(_562_), .Y(_563_) );
AND2X2 AND2X2_32 ( .A(_425__bF_buf2), .B(micro_hash_ucr_Wx_224_), .Y(_564_) );
OAI21X1 OAI21X1_176 ( .A(_425__bF_buf2), .B(micro_hash_ucr_Wx_224_), .C(micro_hash_ucr_pipe64_bF_buf3), .Y(_565_) );
NOR2X1 NOR2X1_249 ( .A(_565_), .B(_564_), .Y(_566_) );
NOR2X1 NOR2X1_250 ( .A(micro_hash_ucr_pipe66_bF_buf1), .B(_566_), .Y(_567_) );
OAI21X1 OAI21X1_177 ( .A(_558_), .B(_563_), .C(_567_), .Y(_568_) );
NOR2X1 NOR2X1_251 ( .A(micro_hash_ucr_Wx_232_), .B(_425__bF_buf2), .Y(_569_) );
NAND2X1 NAND2X1_144 ( .A(micro_hash_ucr_Wx_232_), .B(_425__bF_buf2), .Y(_570_) );
INVX1 INVX1_90 ( .A(_570_), .Y(_571_) );
OAI21X1 OAI21X1_178 ( .A(_571_), .B(_569_), .C(micro_hash_ucr_pipe66_bF_buf1), .Y(_572_) );
AND2X2 AND2X2_33 ( .A(_568_), .B(_572_), .Y(_573_) );
NOR2X1 NOR2X1_252 ( .A(micro_hash_ucr_Wx_240_), .B(_425__bF_buf3), .Y(_574_) );
INVX1 INVX1_91 ( .A(micro_hash_ucr_Wx_240_), .Y(_575_) );
NOR2X1 NOR2X1_253 ( .A(_575_), .B(_426__bF_buf1), .Y(_576_) );
OAI21X1 OAI21X1_179 ( .A(_576_), .B(_574_), .C(micro_hash_ucr_pipe68), .Y(_577_) );
OAI21X1 OAI21X1_180 ( .A(_573_), .B(micro_hash_ucr_pipe68), .C(_577_), .Y(_578_) );
INVX2 INVX2_39 ( .A(micro_hash_ucr_Wx_248_), .Y(_579_) );
AOI21X1 AOI21X1_74 ( .A(_579_), .B(_426__bF_buf1), .C(_292__bF_buf8), .Y(_580_) );
OAI21X1 OAI21X1_181 ( .A(_579_), .B(_426__bF_buf1), .C(_580_), .Y(_581_) );
AOI22X1 AOI22X1_11 ( .A(_345_), .B(_581_), .C(_578_), .D(_287_), .Y(_128__0_) );
NAND2X1 NAND2X1_145 ( .A(micro_hash_ucr_Wx_160_), .B(_425__bF_buf4), .Y(_582_) );
NOR2X1 NOR2X1_254 ( .A(micro_hash_ucr_k_1_), .B(micro_hash_ucr_x_1_), .Y(_583_) );
AND2X2 AND2X2_34 ( .A(micro_hash_ucr_k_1_), .B(micro_hash_ucr_x_1_), .Y(_584_) );
NOR2X1 NOR2X1_255 ( .A(_583_), .B(_584_), .Y(_585_) );
AND2X2 AND2X2_35 ( .A(_585_), .B(_423_), .Y(_586_) );
NOR2X1 NOR2X1_256 ( .A(_423_), .B(_585_), .Y(_587_) );
NOR2X1 NOR2X1_257 ( .A(_587_), .B(_586_), .Y(_588_) );
XNOR2X1 XNOR2X1_8 ( .A(_588__bF_buf2), .B(micro_hash_ucr_Wx_161_), .Y(_589_) );
XNOR2X1 XNOR2X1_9 ( .A(_589_), .B(_582_), .Y(_590_) );
INVX8 INVX8_54 ( .A(micro_hash_ucr_c_1_bF_buf3_), .Y(_591_) );
NOR2X1 NOR2X1_258 ( .A(micro_hash_ucr_pipe6), .B(_591__bF_buf3), .Y(_592_) );
INVX2 INVX2_40 ( .A(H_17_), .Y(_593_) );
OAI21X1 OAI21X1_182 ( .A(_4252_), .B(_593_), .C(_438_), .Y(_594_) );
INVX1 INVX1_92 ( .A(micro_hash_ucr_Wx_1_), .Y(_595_) );
OAI21X1 OAI21X1_183 ( .A(_586_), .B(_587_), .C(_595_), .Y(_596_) );
INVX8 INVX8_55 ( .A(_588__bF_buf2), .Y(_597_) );
NOR2X1 NOR2X1_259 ( .A(_595_), .B(_597__bF_buf4), .Y(_598_) );
INVX1 INVX1_93 ( .A(_598_), .Y(_599_) );
NAND2X1 NAND2X1_146 ( .A(_596_), .B(_599_), .Y(_600_) );
XNOR2X1 XNOR2X1_10 ( .A(_600_), .B(_440_), .Y(_601_) );
OAI22X1 OAI22X1_17 ( .A(_592_), .B(_594_), .C(_601_), .D(_438_), .Y(_602_) );
INVX1 INVX1_94 ( .A(micro_hash_ucr_Wx_9_), .Y(_603_) );
OAI21X1 OAI21X1_184 ( .A(_586_), .B(_587_), .C(_603_), .Y(_604_) );
INVX1 INVX1_95 ( .A(_604_), .Y(_605_) );
NOR2X1 NOR2X1_260 ( .A(_603_), .B(_597__bF_buf4), .Y(_606_) );
NOR2X1 NOR2X1_261 ( .A(_605_), .B(_606_), .Y(_607_) );
XNOR2X1 XNOR2X1_11 ( .A(_607_), .B(_436_), .Y(_608_) );
MUX2X1 MUX2X1_34 ( .A(_602_), .B(_608_), .S(_4243_), .Y(_609_) );
INVX2 INVX2_41 ( .A(micro_hash_ucr_Wx_17_), .Y(_610_) );
OAI21X1 OAI21X1_185 ( .A(_586_), .B(_587_), .C(_610_), .Y(_611_) );
NAND2X1 NAND2X1_147 ( .A(micro_hash_ucr_Wx_17_), .B(_588__bF_buf0), .Y(_612_) );
NAND2X1 NAND2X1_148 ( .A(_611_), .B(_612_), .Y(_613_) );
XOR2X1 XOR2X1_2 ( .A(_613_), .B(_448_), .Y(_614_) );
MUX2X1 MUX2X1_35 ( .A(_609_), .B(_614_), .S(_4258_), .Y(_615_) );
INVX2 INVX2_42 ( .A(micro_hash_ucr_Wx_25_), .Y(_616_) );
OAI21X1 OAI21X1_186 ( .A(_586_), .B(_587_), .C(_616_), .Y(_617_) );
INVX1 INVX1_96 ( .A(_617_), .Y(_618_) );
NOR2X1 NOR2X1_262 ( .A(_616_), .B(_597__bF_buf4), .Y(_619_) );
NOR2X1 NOR2X1_263 ( .A(_618_), .B(_619_), .Y(_620_) );
XNOR2X1 XNOR2X1_12 ( .A(_620_), .B(_432_), .Y(_621_) );
MUX2X1 MUX2X1_36 ( .A(_615_), .B(_621_), .S(_4241__bF_buf1), .Y(_622_) );
NOR2X1 NOR2X1_264 ( .A(micro_hash_ucr_pipe16), .B(_622_), .Y(_623_) );
INVX8 INVX8_56 ( .A(micro_hash_ucr_pipe18_bF_buf2), .Y(_624_) );
INVX2 INVX2_43 ( .A(micro_hash_ucr_Wx_33_), .Y(_625_) );
OAI21X1 OAI21X1_187 ( .A(_586_), .B(_587_), .C(_625_), .Y(_626_) );
NAND2X1 NAND2X1_149 ( .A(micro_hash_ucr_Wx_33_), .B(_588__bF_buf0), .Y(_627_) );
NAND2X1 NAND2X1_150 ( .A(_626_), .B(_627_), .Y(_628_) );
XNOR2X1 XNOR2X1_13 ( .A(_628_), .B(_456_), .Y(_629_) );
OAI21X1 OAI21X1_188 ( .A(_629_), .B(_4239__bF_buf2), .C(_624__bF_buf0), .Y(_630_) );
INVX4 INVX4_11 ( .A(micro_hash_ucr_Wx_41_), .Y(_631_) );
XNOR2X1 XNOR2X1_14 ( .A(_588__bF_buf0), .B(_631_), .Y(_632_) );
XOR2X1 XOR2X1_3 ( .A(_632_), .B(_462_), .Y(_633_) );
AOI21X1 AOI21X1_75 ( .A(micro_hash_ucr_pipe18_bF_buf3), .B(_633_), .C(micro_hash_ucr_pipe20_bF_buf1), .Y(_634_) );
OAI21X1 OAI21X1_189 ( .A(_623_), .B(_630_), .C(_634_), .Y(_635_) );
INVX1 INVX1_97 ( .A(_468_), .Y(_636_) );
INVX2 INVX2_44 ( .A(micro_hash_ucr_Wx_49_), .Y(_637_) );
OAI21X1 OAI21X1_190 ( .A(_586_), .B(_587_), .C(_637_), .Y(_638_) );
NOR2X1 NOR2X1_265 ( .A(_637_), .B(_597__bF_buf4), .Y(_639_) );
INVX2 INVX2_45 ( .A(_639_), .Y(_640_) );
NAND2X1 NAND2X1_151 ( .A(_638_), .B(_640_), .Y(_641_) );
NOR2X1 NOR2X1_266 ( .A(_636_), .B(_641_), .Y(_642_) );
AOI21X1 AOI21X1_76 ( .A(_638_), .B(_640_), .C(_468_), .Y(_643_) );
OAI21X1 OAI21X1_191 ( .A(_642_), .B(_643_), .C(micro_hash_ucr_pipe20_bF_buf1), .Y(_644_) );
NAND3X1 NAND3X1_73 ( .A(_4262__bF_buf3), .B(_644_), .C(_635_), .Y(_645_) );
XNOR2X1 XNOR2X1_15 ( .A(_588__bF_buf1), .B(micro_hash_ucr_Wx_57_), .Y(_646_) );
OAI21X1 OAI21X1_192 ( .A(_471_), .B(_426__bF_buf3), .C(_646_), .Y(_647_) );
INVX1 INVX1_98 ( .A(_646_), .Y(_648_) );
AOI21X1 AOI21X1_77 ( .A(_472_), .B(_648_), .C(_4262__bF_buf3), .Y(_649_) );
AOI21X1 AOI21X1_78 ( .A(_647_), .B(_649_), .C(micro_hash_ucr_pipe24_bF_buf1), .Y(_650_) );
INVX2 INVX2_46 ( .A(micro_hash_ucr_Wx_65_), .Y(_651_) );
OAI21X1 OAI21X1_193 ( .A(_586_), .B(_587_), .C(_651_), .Y(_652_) );
NAND2X1 NAND2X1_152 ( .A(micro_hash_ucr_Wx_65_), .B(_588__bF_buf0), .Y(_653_) );
NAND2X1 NAND2X1_153 ( .A(_652_), .B(_653_), .Y(_654_) );
XNOR2X1 XNOR2X1_16 ( .A(_654_), .B(_478_), .Y(_655_) );
OAI21X1 OAI21X1_194 ( .A(_655_), .B(_4233__bF_buf0), .C(_4230__bF_buf4), .Y(_656_) );
AOI21X1 AOI21X1_79 ( .A(_650_), .B(_645_), .C(_656_), .Y(_657_) );
INVX1 INVX1_99 ( .A(_484_), .Y(_658_) );
XNOR2X1 XNOR2X1_17 ( .A(_588__bF_buf1), .B(micro_hash_ucr_Wx_73_), .Y(_659_) );
NOR2X1 NOR2X1_267 ( .A(_658_), .B(_659_), .Y(_660_) );
INVX1 INVX1_100 ( .A(_660_), .Y(_661_) );
AOI21X1 AOI21X1_80 ( .A(_658_), .B(_659_), .C(_4230__bF_buf4), .Y(_662_) );
AOI21X1 AOI21X1_81 ( .A(_661_), .B(_662_), .C(_657_), .Y(_663_) );
INVX2 INVX2_47 ( .A(micro_hash_ucr_Wx_81_), .Y(_664_) );
OAI21X1 OAI21X1_195 ( .A(_586_), .B(_587_), .C(_664_), .Y(_665_) );
NAND2X1 NAND2X1_154 ( .A(micro_hash_ucr_Wx_81_), .B(_588__bF_buf0), .Y(_666_) );
NAND2X1 NAND2X1_155 ( .A(_665_), .B(_666_), .Y(_667_) );
XOR2X1 XOR2X1_4 ( .A(_667_), .B(_487_), .Y(_668_) );
NAND2X1 NAND2X1_156 ( .A(micro_hash_ucr_pipe28_bF_buf3), .B(_668_), .Y(_669_) );
OAI21X1 OAI21X1_196 ( .A(_663_), .B(micro_hash_ucr_pipe28_bF_buf3), .C(_669_), .Y(_670_) );
INVX4 INVX4_12 ( .A(micro_hash_ucr_Wx_89_), .Y(_671_) );
XNOR2X1 XNOR2X1_18 ( .A(_588__bF_buf1), .B(_671_), .Y(_672_) );
NAND2X1 NAND2X1_157 ( .A(_494_), .B(_672_), .Y(_673_) );
INVX1 INVX1_101 ( .A(_673_), .Y(_674_) );
NOR2X1 NOR2X1_268 ( .A(_494_), .B(_672_), .Y(_675_) );
OAI21X1 OAI21X1_197 ( .A(_674_), .B(_675_), .C(micro_hash_ucr_pipe30_bF_buf1), .Y(_676_) );
OAI21X1 OAI21X1_198 ( .A(_670_), .B(micro_hash_ucr_pipe30_bF_buf1), .C(_676_), .Y(_677_) );
XNOR2X1 XNOR2X1_19 ( .A(_588__bF_buf1), .B(micro_hash_ucr_Wx_97_), .Y(_678_) );
NOR2X1 NOR2X1_269 ( .A(_497_), .B(_678_), .Y(_679_) );
INVX1 INVX1_102 ( .A(_679_), .Y(_680_) );
AOI21X1 AOI21X1_82 ( .A(_497_), .B(_678_), .C(_4226__bF_buf0), .Y(_681_) );
AOI21X1 AOI21X1_83 ( .A(_681_), .B(_680_), .C(micro_hash_ucr_pipe34_bF_buf2), .Y(_682_) );
OAI21X1 OAI21X1_199 ( .A(_677_), .B(micro_hash_ucr_pipe32_bF_buf3), .C(_682_), .Y(_683_) );
INVX1 INVX1_103 ( .A(_504_), .Y(_684_) );
INVX2 INVX2_48 ( .A(micro_hash_ucr_Wx_105_), .Y(_685_) );
OAI21X1 OAI21X1_200 ( .A(_586_), .B(_587_), .C(_685_), .Y(_686_) );
NOR2X1 NOR2X1_270 ( .A(_685_), .B(_597__bF_buf3), .Y(_687_) );
INVX2 INVX2_49 ( .A(_687_), .Y(_688_) );
NAND2X1 NAND2X1_158 ( .A(_686_), .B(_688_), .Y(_689_) );
NOR2X1 NOR2X1_271 ( .A(_684_), .B(_689_), .Y(_690_) );
AOI21X1 AOI21X1_84 ( .A(_686_), .B(_688_), .C(_504_), .Y(_691_) );
OAI21X1 OAI21X1_201 ( .A(_690_), .B(_691_), .C(micro_hash_ucr_pipe34_bF_buf2), .Y(_692_) );
NAND3X1 NAND3X1_74 ( .A(_4224__bF_buf4), .B(_692_), .C(_683_), .Y(_693_) );
XNOR2X1 XNOR2X1_20 ( .A(_588__bF_buf1), .B(micro_hash_ucr_Wx_113_), .Y(_694_) );
OAI21X1 OAI21X1_202 ( .A(_507_), .B(_426__bF_buf2), .C(_694_), .Y(_695_) );
INVX1 INVX1_104 ( .A(_694_), .Y(_696_) );
NAND2X1 NAND2X1_159 ( .A(_508_), .B(_696_), .Y(_697_) );
NAND2X1 NAND2X1_160 ( .A(_695_), .B(_697_), .Y(_698_) );
OAI21X1 OAI21X1_203 ( .A(_4224__bF_buf4), .B(_698_), .C(_693_), .Y(_699_) );
NOR2X1 NOR2X1_272 ( .A(micro_hash_ucr_pipe38_bF_buf3), .B(_699_), .Y(_700_) );
INVX8 INVX8_57 ( .A(micro_hash_ucr_pipe38_bF_buf0), .Y(_701_) );
INVX2 INVX2_50 ( .A(micro_hash_ucr_Wx_121_), .Y(_702_) );
OAI21X1 OAI21X1_204 ( .A(_586_), .B(_587_), .C(_702_), .Y(_703_) );
INVX1 INVX1_105 ( .A(_703_), .Y(_704_) );
NOR2X1 NOR2X1_273 ( .A(_702_), .B(_597__bF_buf1), .Y(_705_) );
NOR2X1 NOR2X1_274 ( .A(_704_), .B(_705_), .Y(_706_) );
XOR2X1 XOR2X1_5 ( .A(_706_), .B(_513_), .Y(_707_) );
OAI21X1 OAI21X1_205 ( .A(_707_), .B(_701__bF_buf2), .C(_296__bF_buf2), .Y(_708_) );
INVX4 INVX4_13 ( .A(micro_hash_ucr_Wx_129_), .Y(_709_) );
XNOR2X1 XNOR2X1_21 ( .A(_588__bF_buf1), .B(_709_), .Y(_710_) );
NAND2X1 NAND2X1_161 ( .A(_517_), .B(_710_), .Y(_711_) );
INVX1 INVX1_106 ( .A(_711_), .Y(_712_) );
OAI21X1 OAI21X1_206 ( .A(_710_), .B(_517_), .C(micro_hash_ucr_pipe40_bF_buf4), .Y(_713_) );
OAI22X1 OAI22X1_18 ( .A(_712_), .B(_713_), .C(_700_), .D(_708_), .Y(_714_) );
INVX4 INVX4_14 ( .A(micro_hash_ucr_Wx_137_), .Y(_715_) );
XNOR2X1 XNOR2X1_22 ( .A(_588__bF_buf3), .B(_715_), .Y(_716_) );
NOR2X1 NOR2X1_275 ( .A(_524_), .B(_716_), .Y(_717_) );
NAND2X1 NAND2X1_162 ( .A(_524_), .B(_716_), .Y(_718_) );
NAND2X1 NAND2X1_163 ( .A(micro_hash_ucr_pipe42_bF_buf2), .B(_718_), .Y(_719_) );
OAI21X1 OAI21X1_207 ( .A(_719_), .B(_717_), .C(_4219__bF_buf2), .Y(_720_) );
AOI21X1 AOI21X1_85 ( .A(_4220__bF_buf0), .B(_714_), .C(_720_), .Y(_721_) );
INVX2 INVX2_51 ( .A(micro_hash_ucr_Wx_145_), .Y(_722_) );
XNOR2X1 XNOR2X1_23 ( .A(_588__bF_buf3), .B(_722_), .Y(_723_) );
AND2X2 AND2X2_36 ( .A(_723_), .B(_527_), .Y(_724_) );
NOR2X1 NOR2X1_276 ( .A(_527_), .B(_723_), .Y(_725_) );
OAI21X1 OAI21X1_208 ( .A(_724_), .B(_725_), .C(micro_hash_ucr_pipe44_bF_buf1), .Y(_726_) );
NAND2X1 NAND2X1_164 ( .A(_4218__bF_buf3), .B(_726_), .Y(_727_) );
NOR2X1 NOR2X1_277 ( .A(_727_), .B(_721_), .Y(_728_) );
INVX2 INVX2_52 ( .A(micro_hash_ucr_Wx_153_), .Y(_729_) );
XNOR2X1 XNOR2X1_24 ( .A(_588__bF_buf2), .B(_729_), .Y(_730_) );
OAI21X1 OAI21X1_209 ( .A(_730_), .B(_531_), .C(micro_hash_ucr_pipe46_bF_buf0), .Y(_731_) );
AOI21X1 AOI21X1_86 ( .A(_531_), .B(_730_), .C(_731_), .Y(_732_) );
OAI21X1 OAI21X1_210 ( .A(_728_), .B(_732_), .C(_4217__bF_buf1), .Y(_733_) );
OAI21X1 OAI21X1_211 ( .A(_4217__bF_buf1), .B(_590_), .C(_733_), .Y(_734_) );
INVX2 INVX2_53 ( .A(micro_hash_ucr_Wx_169_), .Y(_735_) );
XNOR2X1 XNOR2X1_25 ( .A(_588__bF_buf4), .B(_735_), .Y(_736_) );
NOR2X1 NOR2X1_278 ( .A(_539_), .B(_736_), .Y(_737_) );
NAND2X1 NAND2X1_165 ( .A(_539_), .B(_736_), .Y(_738_) );
NAND2X1 NAND2X1_166 ( .A(micro_hash_ucr_pipe50_bF_buf0), .B(_738_), .Y(_739_) );
OAI21X1 OAI21X1_212 ( .A(_739_), .B(_737_), .C(_4214__bF_buf1), .Y(_740_) );
AOI21X1 AOI21X1_87 ( .A(_4215__bF_buf4), .B(_734_), .C(_740_), .Y(_741_) );
INVX8 INVX8_58 ( .A(micro_hash_ucr_pipe54_bF_buf1), .Y(_742_) );
INVX2 INVX2_54 ( .A(micro_hash_ucr_Wx_177_), .Y(_743_) );
XNOR2X1 XNOR2X1_26 ( .A(_588__bF_buf2), .B(_743_), .Y(_744_) );
AND2X2 AND2X2_37 ( .A(_744_), .B(_542_), .Y(_745_) );
NOR2X1 NOR2X1_279 ( .A(_542_), .B(_744_), .Y(_746_) );
OAI21X1 OAI21X1_213 ( .A(_745_), .B(_746_), .C(micro_hash_ucr_pipe52_bF_buf3), .Y(_747_) );
NAND2X1 NAND2X1_167 ( .A(_742__bF_buf3), .B(_747_), .Y(_748_) );
INVX2 INVX2_55 ( .A(micro_hash_ucr_Wx_185_), .Y(_749_) );
XNOR2X1 XNOR2X1_27 ( .A(_588__bF_buf3), .B(_749_), .Y(_750_) );
NAND2X1 NAND2X1_168 ( .A(_546_), .B(_750_), .Y(_751_) );
INVX1 INVX1_107 ( .A(_751_), .Y(_752_) );
OAI21X1 OAI21X1_214 ( .A(_750_), .B(_546_), .C(micro_hash_ucr_pipe54_bF_buf0), .Y(_753_) );
OAI22X1 OAI22X1_19 ( .A(_752_), .B(_753_), .C(_741_), .D(_748_), .Y(_754_) );
INVX2 INVX2_56 ( .A(micro_hash_ucr_Wx_193_), .Y(_755_) );
XNOR2X1 XNOR2X1_28 ( .A(_588__bF_buf3), .B(_755_), .Y(_756_) );
NAND2X1 NAND2X1_169 ( .A(_550_), .B(_756_), .Y(_757_) );
INVX1 INVX1_108 ( .A(_757_), .Y(_758_) );
NOR2X1 NOR2X1_280 ( .A(_550_), .B(_756_), .Y(_759_) );
OAI21X1 OAI21X1_215 ( .A(_758_), .B(_759_), .C(micro_hash_ucr_pipe56_bF_buf1), .Y(_760_) );
OAI21X1 OAI21X1_216 ( .A(_754_), .B(micro_hash_ucr_pipe56_bF_buf1), .C(_760_), .Y(_761_) );
INVX2 INVX2_57 ( .A(micro_hash_ucr_Wx_201_), .Y(_762_) );
OAI21X1 OAI21X1_217 ( .A(_586_), .B(_587_), .C(_762_), .Y(_763_) );
INVX1 INVX1_109 ( .A(_763_), .Y(_764_) );
NOR2X1 NOR2X1_281 ( .A(_762_), .B(_597__bF_buf1), .Y(_765_) );
OAI21X1 OAI21X1_218 ( .A(_765_), .B(_764_), .C(_428_), .Y(_766_) );
NOR2X1 NOR2X1_282 ( .A(_764_), .B(_765_), .Y(_767_) );
NAND2X1 NAND2X1_170 ( .A(_427_), .B(_767_), .Y(_768_) );
INVX1 INVX1_110 ( .A(_768_), .Y(_769_) );
NOR2X1 NOR2X1_283 ( .A(_4211__bF_buf2), .B(_769_), .Y(_770_) );
AOI21X1 AOI21X1_88 ( .A(_766_), .B(_770_), .C(micro_hash_ucr_pipe60_bF_buf0), .Y(_771_) );
OAI21X1 OAI21X1_219 ( .A(_761_), .B(micro_hash_ucr_pipe58_bF_buf1), .C(_771_), .Y(_772_) );
NAND2X1 NAND2X1_171 ( .A(micro_hash_ucr_Wx_208_), .B(_425__bF_buf2), .Y(_773_) );
NOR2X1 NOR2X1_284 ( .A(micro_hash_ucr_Wx_209_), .B(_588__bF_buf3), .Y(_774_) );
INVX1 INVX1_111 ( .A(_774_), .Y(_775_) );
NAND2X1 NAND2X1_172 ( .A(micro_hash_ucr_Wx_209_), .B(_588__bF_buf3), .Y(_776_) );
NAND2X1 NAND2X1_173 ( .A(_776_), .B(_775_), .Y(_777_) );
XNOR2X1 XNOR2X1_29 ( .A(_777_), .B(_773_), .Y(_778_) );
AOI21X1 AOI21X1_89 ( .A(micro_hash_ucr_pipe60_bF_buf0), .B(_778_), .C(micro_hash_ucr_pipe62_bF_buf1), .Y(_779_) );
INVX2 INVX2_58 ( .A(micro_hash_ucr_Wx_217_), .Y(_780_) );
XNOR2X1 XNOR2X1_30 ( .A(_588__bF_buf4), .B(_780_), .Y(_781_) );
NAND2X1 NAND2X1_174 ( .A(_561_), .B(_781_), .Y(_782_) );
INVX1 INVX1_112 ( .A(_782_), .Y(_783_) );
NOR2X1 NOR2X1_285 ( .A(_561_), .B(_781_), .Y(_784_) );
NOR2X1 NOR2X1_286 ( .A(_784_), .B(_783_), .Y(_785_) );
AOI22X1 AOI22X1_12 ( .A(micro_hash_ucr_pipe62_bF_buf1), .B(_785_), .C(_772_), .D(_779_), .Y(_786_) );
INVX2 INVX2_59 ( .A(micro_hash_ucr_Wx_225_), .Y(_787_) );
XNOR2X1 XNOR2X1_31 ( .A(_588__bF_buf4), .B(_787_), .Y(_788_) );
XOR2X1 XOR2X1_6 ( .A(_788_), .B(_564_), .Y(_789_) );
AOI21X1 AOI21X1_90 ( .A(micro_hash_ucr_pipe64_bF_buf3), .B(_789_), .C(micro_hash_ucr_pipe66_bF_buf1), .Y(_790_) );
OAI21X1 OAI21X1_220 ( .A(_786_), .B(micro_hash_ucr_pipe64_bF_buf3), .C(_790_), .Y(_791_) );
INVX1 INVX1_113 ( .A(micro_hash_ucr_Wx_233_), .Y(_792_) );
OAI21X1 OAI21X1_221 ( .A(_586_), .B(_587_), .C(_792_), .Y(_793_) );
NOR2X1 NOR2X1_287 ( .A(_792_), .B(_597__bF_buf2), .Y(_794_) );
INVX2 INVX2_60 ( .A(_794_), .Y(_795_) );
NAND2X1 NAND2X1_175 ( .A(_793_), .B(_795_), .Y(_796_) );
NOR2X1 NOR2X1_288 ( .A(_570_), .B(_796_), .Y(_797_) );
AOI21X1 AOI21X1_91 ( .A(_793_), .B(_795_), .C(_571_), .Y(_798_) );
OAI21X1 OAI21X1_222 ( .A(_797_), .B(_798_), .C(micro_hash_ucr_pipe66_bF_buf1), .Y(_799_) );
AND2X2 AND2X2_38 ( .A(_791_), .B(_799_), .Y(_800_) );
INVX1 INVX1_114 ( .A(_576_), .Y(_801_) );
XNOR2X1 XNOR2X1_32 ( .A(_588__bF_buf4), .B(micro_hash_ucr_Wx_241_), .Y(_802_) );
NOR2X1 NOR2X1_289 ( .A(_801_), .B(_802_), .Y(_803_) );
AND2X2 AND2X2_39 ( .A(_802_), .B(_801_), .Y(_804_) );
OAI21X1 OAI21X1_223 ( .A(_804_), .B(_803_), .C(micro_hash_ucr_pipe68), .Y(_805_) );
OAI21X1 OAI21X1_224 ( .A(_800_), .B(micro_hash_ucr_pipe68), .C(_805_), .Y(_806_) );
NOR2X1 NOR2X1_290 ( .A(_579_), .B(_426__bF_buf1), .Y(_807_) );
INVX2 INVX2_61 ( .A(micro_hash_ucr_Wx_249_), .Y(_808_) );
XNOR2X1 XNOR2X1_33 ( .A(_588__bF_buf4), .B(_808_), .Y(_809_) );
AND2X2 AND2X2_40 ( .A(_809_), .B(_807_), .Y(_810_) );
NOR2X1 NOR2X1_291 ( .A(_807_), .B(_809_), .Y(_811_) );
OAI21X1 OAI21X1_225 ( .A(_810_), .B(_811_), .C(micro_hash_ucr_pipe69), .Y(_812_) );
NAND2X1 NAND2X1_176 ( .A(_131__bF_buf3), .B(_812_), .Y(_813_) );
AOI21X1 AOI21X1_92 ( .A(_287_), .B(_806_), .C(_813_), .Y(_128__1_) );
OAI21X1 OAI21X1_226 ( .A(_774_), .B(_773_), .C(_776_), .Y(_814_) );
INVX2 INVX2_62 ( .A(micro_hash_ucr_Wx_210_), .Y(_815_) );
NOR2X1 NOR2X1_292 ( .A(_584_), .B(_586_), .Y(_816_) );
INVX1 INVX1_115 ( .A(micro_hash_ucr_k_2_), .Y(_817_) );
INVX1 INVX1_116 ( .A(micro_hash_ucr_x_2_), .Y(_818_) );
NAND2X1 NAND2X1_177 ( .A(_817_), .B(_818_), .Y(_819_) );
NOR2X1 NOR2X1_293 ( .A(_817_), .B(_818_), .Y(_820_) );
INVX1 INVX1_117 ( .A(_820_), .Y(_821_) );
NAND2X1 NAND2X1_178 ( .A(_819_), .B(_821_), .Y(_822_) );
NOR2X1 NOR2X1_294 ( .A(_822_), .B(_816_), .Y(_823_) );
AND2X2 AND2X2_41 ( .A(_816_), .B(_822_), .Y(_824_) );
OAI21X1 OAI21X1_227 ( .A(_824__bF_buf1), .B(_823__bF_buf0), .C(_815_), .Y(_825_) );
NOR2X1 NOR2X1_295 ( .A(_823__bF_buf1), .B(_824__bF_buf3), .Y(_826_) );
INVX8 INVX8_59 ( .A(_826__bF_buf1), .Y(_827_) );
NOR2X1 NOR2X1_296 ( .A(_815_), .B(_827__bF_buf1), .Y(_828_) );
INVX1 INVX1_118 ( .A(_828_), .Y(_829_) );
NAND2X1 NAND2X1_179 ( .A(_825_), .B(_829_), .Y(_830_) );
XOR2X1 XOR2X1_7 ( .A(_830_), .B(_814_), .Y(_831_) );
INVX8 INVX8_60 ( .A(micro_hash_ucr_pipe56_bF_buf1), .Y(_832_) );
INVX1 INVX1_119 ( .A(_456_), .Y(_833_) );
OAI21X1 OAI21X1_228 ( .A(_628_), .B(_833_), .C(_627_), .Y(_834_) );
INVX2 INVX2_63 ( .A(micro_hash_ucr_Wx_34_), .Y(_835_) );
OAI21X1 OAI21X1_229 ( .A(_824__bF_buf2), .B(_823__bF_buf3), .C(_835_), .Y(_836_) );
NOR2X1 NOR2X1_297 ( .A(_835_), .B(_827__bF_buf3), .Y(_837_) );
INVX1 INVX1_120 ( .A(_837_), .Y(_838_) );
NAND2X1 NAND2X1_180 ( .A(_836_), .B(_838_), .Y(_839_) );
XNOR2X1 XNOR2X1_34 ( .A(_839_), .B(_834_), .Y(_840_) );
OAI21X1 OAI21X1_230 ( .A(_613_), .B(_448_), .C(_612_), .Y(_841_) );
INVX4 INVX4_15 ( .A(micro_hash_ucr_Wx_18_), .Y(_842_) );
XNOR2X1 XNOR2X1_35 ( .A(_826__bF_buf0), .B(_842_), .Y(_843_) );
XOR2X1 XOR2X1_8 ( .A(_843_), .B(_841_), .Y(_844_) );
INVX8 INVX8_61 ( .A(micro_hash_ucr_c_2_bF_buf3_), .Y(_845_) );
NAND2X1 NAND2X1_181 ( .A(micro_hash_ucr_pipe6), .B(H_18_), .Y(_846_) );
OAI21X1 OAI21X1_231 ( .A(_845__bF_buf0), .B(micro_hash_ucr_pipe6), .C(_846_), .Y(_847_) );
OAI21X1 OAI21X1_232 ( .A(_600_), .B(_439_), .C(_599_), .Y(_848_) );
NOR2X1 NOR2X1_298 ( .A(micro_hash_ucr_Wx_2_), .B(_826__bF_buf0), .Y(_849_) );
NAND2X1 NAND2X1_182 ( .A(micro_hash_ucr_Wx_2_), .B(_826__bF_buf0), .Y(_850_) );
INVX1 INVX1_121 ( .A(_850_), .Y(_851_) );
NOR2X1 NOR2X1_299 ( .A(_849_), .B(_851_), .Y(_852_) );
AND2X2 AND2X2_42 ( .A(_852_), .B(_848_), .Y(_853_) );
NOR2X1 NOR2X1_300 ( .A(_848_), .B(_852_), .Y(_854_) );
OAI21X1 OAI21X1_233 ( .A(_853_), .B(_854_), .C(micro_hash_ucr_pipe8), .Y(_855_) );
OAI21X1 OAI21X1_234 ( .A(micro_hash_ucr_pipe8), .B(_847_), .C(_855_), .Y(_856_) );
AOI21X1 AOI21X1_93 ( .A(_436_), .B(_604_), .C(_606_), .Y(_857_) );
INVX1 INVX1_122 ( .A(_857_), .Y(_858_) );
INVX1 INVX1_123 ( .A(micro_hash_ucr_Wx_10_), .Y(_859_) );
OAI21X1 OAI21X1_235 ( .A(_824__bF_buf2), .B(_823__bF_buf3), .C(_859_), .Y(_860_) );
INVX1 INVX1_124 ( .A(_860_), .Y(_861_) );
NOR2X1 NOR2X1_301 ( .A(_859_), .B(_827__bF_buf3), .Y(_862_) );
NOR2X1 NOR2X1_302 ( .A(_861_), .B(_862_), .Y(_863_) );
NAND2X1 NAND2X1_183 ( .A(_858_), .B(_863_), .Y(_864_) );
OAI21X1 OAI21X1_236 ( .A(_862_), .B(_861_), .C(_857_), .Y(_865_) );
NAND3X1 NAND3X1_75 ( .A(micro_hash_ucr_pipe10), .B(_865_), .C(_864_), .Y(_866_) );
OAI21X1 OAI21X1_237 ( .A(micro_hash_ucr_pipe10), .B(_856_), .C(_866_), .Y(_867_) );
MUX2X1 MUX2X1_37 ( .A(_867_), .B(_844_), .S(_4258_), .Y(_868_) );
AOI21X1 AOI21X1_94 ( .A(_432_), .B(_617_), .C(_619_), .Y(_869_) );
INVX2 INVX2_64 ( .A(micro_hash_ucr_Wx_26_), .Y(_870_) );
OAI21X1 OAI21X1_238 ( .A(_824__bF_buf2), .B(_823__bF_buf3), .C(_870_), .Y(_871_) );
INVX1 INVX1_125 ( .A(_871_), .Y(_872_) );
NOR2X1 NOR2X1_303 ( .A(_870_), .B(_827__bF_buf3), .Y(_873_) );
NOR2X1 NOR2X1_304 ( .A(_872_), .B(_873_), .Y(_874_) );
INVX1 INVX1_126 ( .A(_874_), .Y(_875_) );
NOR2X1 NOR2X1_305 ( .A(_869_), .B(_875_), .Y(_876_) );
INVX1 INVX1_127 ( .A(_876_), .Y(_877_) );
OAI21X1 OAI21X1_239 ( .A(_873_), .B(_872_), .C(_869_), .Y(_878_) );
NAND3X1 NAND3X1_76 ( .A(micro_hash_ucr_pipe14), .B(_878_), .C(_877_), .Y(_879_) );
OAI21X1 OAI21X1_240 ( .A(_868_), .B(micro_hash_ucr_pipe14), .C(_879_), .Y(_880_) );
MUX2X1 MUX2X1_38 ( .A(_880_), .B(_840_), .S(_4239__bF_buf2), .Y(_881_) );
NAND2X1 NAND2X1_184 ( .A(_462_), .B(_632_), .Y(_882_) );
OAI21X1 OAI21X1_241 ( .A(_631_), .B(_597__bF_buf4), .C(_882_), .Y(_883_) );
INVX2 INVX2_65 ( .A(micro_hash_ucr_Wx_42_), .Y(_884_) );
OAI21X1 OAI21X1_242 ( .A(_824__bF_buf2), .B(_823__bF_buf3), .C(_884_), .Y(_885_) );
NOR2X1 NOR2X1_306 ( .A(_884_), .B(_827__bF_buf4), .Y(_886_) );
INVX1 INVX1_128 ( .A(_886_), .Y(_887_) );
NAND2X1 NAND2X1_185 ( .A(_885_), .B(_887_), .Y(_888_) );
XOR2X1 XOR2X1_9 ( .A(_888_), .B(_883_), .Y(_889_) );
MUX2X1 MUX2X1_39 ( .A(_881_), .B(_889_), .S(_624__bF_buf0), .Y(_890_) );
INVX4 INVX4_16 ( .A(micro_hash_ucr_Wx_50_), .Y(_891_) );
XNOR2X1 XNOR2X1_36 ( .A(_826__bF_buf0), .B(_891_), .Y(_892_) );
OAI21X1 OAI21X1_243 ( .A(_642_), .B(_639_), .C(_892_), .Y(_893_) );
INVX1 INVX1_129 ( .A(_893_), .Y(_894_) );
OAI21X1 OAI21X1_244 ( .A(_641_), .B(_636_), .C(_640_), .Y(_895_) );
NOR2X1 NOR2X1_307 ( .A(_892_), .B(_895_), .Y(_896_) );
OAI21X1 OAI21X1_245 ( .A(_894_), .B(_896_), .C(micro_hash_ucr_pipe20_bF_buf1), .Y(_897_) );
OAI21X1 OAI21X1_246 ( .A(_890_), .B(micro_hash_ucr_pipe20_bF_buf1), .C(_897_), .Y(_898_) );
NOR2X1 NOR2X1_308 ( .A(micro_hash_ucr_pipe22_bF_buf1), .B(_898_), .Y(_899_) );
INVX2 INVX2_66 ( .A(micro_hash_ucr_Wx_57_), .Y(_900_) );
NAND2X1 NAND2X1_186 ( .A(_472_), .B(_648_), .Y(_901_) );
OAI21X1 OAI21X1_247 ( .A(_900_), .B(_597__bF_buf4), .C(_901_), .Y(_902_) );
INVX4 INVX4_17 ( .A(micro_hash_ucr_Wx_58_), .Y(_903_) );
XNOR2X1 XNOR2X1_37 ( .A(_826__bF_buf2), .B(_903_), .Y(_904_) );
NOR2X1 NOR2X1_309 ( .A(_904_), .B(_902_), .Y(_905_) );
NAND2X1 NAND2X1_187 ( .A(_904_), .B(_902_), .Y(_906_) );
NAND2X1 NAND2X1_188 ( .A(micro_hash_ucr_pipe22_bF_buf1), .B(_906_), .Y(_907_) );
OAI21X1 OAI21X1_248 ( .A(_907_), .B(_905_), .C(_4233__bF_buf0), .Y(_908_) );
INVX1 INVX1_130 ( .A(_478_), .Y(_909_) );
OAI21X1 OAI21X1_249 ( .A(_654_), .B(_909_), .C(_653_), .Y(_910_) );
INVX2 INVX2_67 ( .A(micro_hash_ucr_Wx_66_), .Y(_911_) );
OAI21X1 OAI21X1_250 ( .A(_824__bF_buf2), .B(_823__bF_buf2), .C(_911_), .Y(_912_) );
NOR2X1 NOR2X1_310 ( .A(_911_), .B(_827__bF_buf4), .Y(_913_) );
INVX1 INVX1_131 ( .A(_913_), .Y(_914_) );
NAND2X1 NAND2X1_189 ( .A(_912_), .B(_914_), .Y(_915_) );
XOR2X1 XOR2X1_10 ( .A(_915_), .B(_910_), .Y(_916_) );
AOI21X1 AOI21X1_95 ( .A(micro_hash_ucr_pipe24_bF_buf1), .B(_916_), .C(micro_hash_ucr_pipe26_bF_buf0), .Y(_917_) );
OAI21X1 OAI21X1_251 ( .A(_899_), .B(_908_), .C(_917_), .Y(_918_) );
INVX2 INVX2_68 ( .A(micro_hash_ucr_Wx_73_), .Y(_919_) );
OAI21X1 OAI21X1_252 ( .A(_919_), .B(_597__bF_buf3), .C(_661_), .Y(_920_) );
INVX2 INVX2_69 ( .A(micro_hash_ucr_Wx_74_), .Y(_921_) );
OAI21X1 OAI21X1_253 ( .A(_824__bF_buf0), .B(_823__bF_buf2), .C(_921_), .Y(_922_) );
INVX1 INVX1_132 ( .A(_922_), .Y(_923_) );
NOR2X1 NOR2X1_311 ( .A(_921_), .B(_827__bF_buf4), .Y(_924_) );
NOR2X1 NOR2X1_312 ( .A(_923_), .B(_924_), .Y(_925_) );
AND2X2 AND2X2_43 ( .A(_925_), .B(_920_), .Y(_926_) );
OAI21X1 OAI21X1_254 ( .A(_925_), .B(_920_), .C(micro_hash_ucr_pipe26_bF_buf0), .Y(_927_) );
OAI21X1 OAI21X1_255 ( .A(_926_), .B(_927_), .C(_918_), .Y(_928_) );
NOR2X1 NOR2X1_313 ( .A(micro_hash_ucr_pipe28_bF_buf3), .B(_928_), .Y(_929_) );
OAI21X1 OAI21X1_256 ( .A(_667_), .B(_487_), .C(_666_), .Y(_930_) );
INVX2 INVX2_70 ( .A(micro_hash_ucr_Wx_82_), .Y(_931_) );
OAI21X1 OAI21X1_257 ( .A(_824__bF_buf0), .B(_823__bF_buf2), .C(_931_), .Y(_932_) );
NOR2X1 NOR2X1_314 ( .A(_931_), .B(_827__bF_buf0), .Y(_933_) );
INVX1 INVX1_133 ( .A(_933_), .Y(_934_) );
NAND2X1 NAND2X1_190 ( .A(_932_), .B(_934_), .Y(_935_) );
XNOR2X1 XNOR2X1_38 ( .A(_935_), .B(_930_), .Y(_936_) );
OAI21X1 OAI21X1_258 ( .A(_936_), .B(_220__bF_buf0), .C(_4228__bF_buf4), .Y(_937_) );
OAI21X1 OAI21X1_259 ( .A(_671_), .B(_597__bF_buf3), .C(_673_), .Y(_938_) );
INVX4 INVX4_18 ( .A(micro_hash_ucr_Wx_90_), .Y(_939_) );
XNOR2X1 XNOR2X1_39 ( .A(_826__bF_buf2), .B(_939_), .Y(_940_) );
XOR2X1 XOR2X1_11 ( .A(_940_), .B(_938_), .Y(_941_) );
AOI21X1 AOI21X1_96 ( .A(micro_hash_ucr_pipe30_bF_buf1), .B(_941_), .C(micro_hash_ucr_pipe32_bF_buf3), .Y(_942_) );
OAI21X1 OAI21X1_260 ( .A(_929_), .B(_937_), .C(_942_), .Y(_943_) );
INVX2 INVX2_71 ( .A(micro_hash_ucr_Wx_97_), .Y(_944_) );
OAI21X1 OAI21X1_261 ( .A(_944_), .B(_597__bF_buf3), .C(_680_), .Y(_945_) );
INVX4 INVX4_19 ( .A(micro_hash_ucr_Wx_98_), .Y(_946_) );
XNOR2X1 XNOR2X1_40 ( .A(_826__bF_buf2), .B(_946_), .Y(_947_) );
NAND2X1 NAND2X1_191 ( .A(_947_), .B(_945_), .Y(_948_) );
INVX1 INVX1_134 ( .A(_948_), .Y(_949_) );
NOR2X1 NOR2X1_315 ( .A(_947_), .B(_945_), .Y(_950_) );
OAI21X1 OAI21X1_262 ( .A(_949_), .B(_950_), .C(micro_hash_ucr_pipe32_bF_buf3), .Y(_951_) );
NAND3X1 NAND3X1_77 ( .A(_4225__bF_buf4), .B(_951_), .C(_943_), .Y(_952_) );
INVX4 INVX4_20 ( .A(micro_hash_ucr_Wx_106_), .Y(_953_) );
XNOR2X1 XNOR2X1_41 ( .A(_826__bF_buf2), .B(_953_), .Y(_954_) );
OAI21X1 OAI21X1_263 ( .A(_690_), .B(_687_), .C(_954_), .Y(_955_) );
INVX1 INVX1_135 ( .A(_955_), .Y(_956_) );
OAI21X1 OAI21X1_264 ( .A(_689_), .B(_684_), .C(_688_), .Y(_957_) );
OAI21X1 OAI21X1_265 ( .A(_957_), .B(_954_), .C(micro_hash_ucr_pipe34_bF_buf2), .Y(_958_) );
OAI21X1 OAI21X1_266 ( .A(_956_), .B(_958_), .C(_952_), .Y(_959_) );
NOR2X1 NOR2X1_316 ( .A(micro_hash_ucr_pipe36_bF_buf1), .B(_959_), .Y(_960_) );
INVX2 INVX2_72 ( .A(micro_hash_ucr_Wx_113_), .Y(_961_) );
OAI21X1 OAI21X1_267 ( .A(_961_), .B(_597__bF_buf3), .C(_697_), .Y(_962_) );
INVX4 INVX4_21 ( .A(micro_hash_ucr_Wx_114_), .Y(_963_) );
OAI21X1 OAI21X1_268 ( .A(_824__bF_buf0), .B(_823__bF_buf2), .C(_963_), .Y(_964_) );
NOR2X1 NOR2X1_317 ( .A(_963_), .B(_827__bF_buf0), .Y(_965_) );
INVX1 INVX1_136 ( .A(_965_), .Y(_966_) );
NAND2X1 NAND2X1_192 ( .A(_964_), .B(_966_), .Y(_967_) );
XNOR2X1 XNOR2X1_42 ( .A(_967_), .B(_962_), .Y(_968_) );
OAI21X1 OAI21X1_269 ( .A(_968_), .B(_4224__bF_buf4), .C(_701__bF_buf2), .Y(_969_) );
AOI21X1 AOI21X1_97 ( .A(_513_), .B(_703_), .C(_705_), .Y(_970_) );
INVX4 INVX4_22 ( .A(micro_hash_ucr_Wx_122_), .Y(_971_) );
OAI21X1 OAI21X1_270 ( .A(_824__bF_buf0), .B(_823__bF_buf2), .C(_971_), .Y(_972_) );
INVX1 INVX1_137 ( .A(_972_), .Y(_973_) );
NOR2X1 NOR2X1_318 ( .A(_971_), .B(_827__bF_buf0), .Y(_974_) );
NOR2X1 NOR2X1_319 ( .A(_973_), .B(_974_), .Y(_975_) );
INVX1 INVX1_138 ( .A(_975_), .Y(_976_) );
NOR2X1 NOR2X1_320 ( .A(_970_), .B(_976_), .Y(_977_) );
INVX1 INVX1_139 ( .A(_977_), .Y(_978_) );
OAI21X1 OAI21X1_271 ( .A(_974_), .B(_973_), .C(_970_), .Y(_979_) );
NAND3X1 NAND3X1_78 ( .A(micro_hash_ucr_pipe38_bF_buf3), .B(_979_), .C(_978_), .Y(_980_) );
OAI21X1 OAI21X1_272 ( .A(_960_), .B(_969_), .C(_980_), .Y(_981_) );
OAI21X1 OAI21X1_273 ( .A(_709_), .B(_597__bF_buf1), .C(_711_), .Y(_982_) );
INVX4 INVX4_23 ( .A(micro_hash_ucr_Wx_130_), .Y(_983_) );
XNOR2X1 XNOR2X1_43 ( .A(_826__bF_buf1), .B(_983_), .Y(_984_) );
NOR2X1 NOR2X1_321 ( .A(_982_), .B(_984_), .Y(_985_) );
NAND2X1 NAND2X1_193 ( .A(_982_), .B(_984_), .Y(_986_) );
NAND2X1 NAND2X1_194 ( .A(micro_hash_ucr_pipe40_bF_buf4), .B(_986_), .Y(_987_) );
OAI21X1 OAI21X1_274 ( .A(_987_), .B(_985_), .C(_4220__bF_buf0), .Y(_988_) );
AOI21X1 AOI21X1_98 ( .A(_296__bF_buf2), .B(_981_), .C(_988_), .Y(_989_) );
OAI21X1 OAI21X1_275 ( .A(_715_), .B(_597__bF_buf0), .C(_718_), .Y(_990_) );
INVX4 INVX4_24 ( .A(micro_hash_ucr_Wx_138_), .Y(_991_) );
OAI21X1 OAI21X1_276 ( .A(_824__bF_buf3), .B(_823__bF_buf1), .C(_991_), .Y(_992_) );
NOR2X1 NOR2X1_322 ( .A(_991_), .B(_827__bF_buf5), .Y(_993_) );
INVX1 INVX1_140 ( .A(_993_), .Y(_994_) );
NAND2X1 NAND2X1_195 ( .A(_992_), .B(_994_), .Y(_995_) );
XNOR2X1 XNOR2X1_44 ( .A(_995_), .B(_990_), .Y(_996_) );
OAI21X1 OAI21X1_277 ( .A(_996_), .B(_4220__bF_buf0), .C(_4219__bF_buf2), .Y(_997_) );
NOR2X1 NOR2X1_323 ( .A(_722_), .B(_597__bF_buf0), .Y(_998_) );
INVX2 INVX2_73 ( .A(micro_hash_ucr_Wx_146_), .Y(_999_) );
OAI21X1 OAI21X1_278 ( .A(_824__bF_buf3), .B(_823__bF_buf1), .C(_999_), .Y(_1000_) );
INVX1 INVX1_141 ( .A(_1000_), .Y(_1001_) );
NOR2X1 NOR2X1_324 ( .A(_999_), .B(_827__bF_buf5), .Y(_1002_) );
NOR2X1 NOR2X1_325 ( .A(_1001_), .B(_1002_), .Y(_1003_) );
OAI21X1 OAI21X1_279 ( .A(_724_), .B(_998_), .C(_1003_), .Y(_1004_) );
NOR2X1 NOR2X1_326 ( .A(_998_), .B(_724_), .Y(_1005_) );
OAI21X1 OAI21X1_280 ( .A(_1002_), .B(_1001_), .C(_1005_), .Y(_1006_) );
NAND2X1 NAND2X1_196 ( .A(_1006_), .B(_1004_), .Y(_1007_) );
OAI22X1 OAI22X1_20 ( .A(_4219__bF_buf2), .B(_1007_), .C(_989_), .D(_997_), .Y(_1008_) );
NAND2X1 NAND2X1_197 ( .A(_531_), .B(_730_), .Y(_1009_) );
OAI21X1 OAI21X1_281 ( .A(_729_), .B(_597__bF_buf0), .C(_1009_), .Y(_1010_) );
INVX2 INVX2_74 ( .A(micro_hash_ucr_Wx_154_), .Y(_1011_) );
XNOR2X1 XNOR2X1_45 ( .A(_826__bF_buf1), .B(_1011_), .Y(_1012_) );
NOR2X1 NOR2X1_327 ( .A(_1010_), .B(_1012_), .Y(_1013_) );
NAND2X1 NAND2X1_198 ( .A(_1010_), .B(_1012_), .Y(_1014_) );
INVX1 INVX1_142 ( .A(_1014_), .Y(_1015_) );
OAI21X1 OAI21X1_282 ( .A(_1015_), .B(_1013_), .C(micro_hash_ucr_pipe46_bF_buf0), .Y(_1016_) );
OAI21X1 OAI21X1_283 ( .A(_1008_), .B(micro_hash_ucr_pipe46_bF_buf0), .C(_1016_), .Y(_1017_) );
NAND2X1 NAND2X1_199 ( .A(micro_hash_ucr_Wx_161_), .B(_588__bF_buf2), .Y(_1018_) );
OAI21X1 OAI21X1_284 ( .A(_589_), .B(_582_), .C(_1018_), .Y(_1019_) );
INVX2 INVX2_75 ( .A(micro_hash_ucr_Wx_162_), .Y(_1020_) );
OAI21X1 OAI21X1_285 ( .A(_824__bF_buf3), .B(_823__bF_buf1), .C(_1020_), .Y(_1021_) );
NOR2X1 NOR2X1_328 ( .A(_1020_), .B(_827__bF_buf5), .Y(_1022_) );
INVX1 INVX1_143 ( .A(_1022_), .Y(_1023_) );
NAND2X1 NAND2X1_200 ( .A(_1021_), .B(_1023_), .Y(_1024_) );
XOR2X1 XOR2X1_12 ( .A(_1024_), .B(_1019_), .Y(_1025_) );
MUX2X1 MUX2X1_40 ( .A(_1017_), .B(_1025_), .S(_4217__bF_buf1), .Y(_1026_) );
OAI21X1 OAI21X1_286 ( .A(_735_), .B(_597__bF_buf0), .C(_738_), .Y(_1027_) );
INVX2 INVX2_76 ( .A(micro_hash_ucr_Wx_170_), .Y(_1028_) );
XNOR2X1 XNOR2X1_46 ( .A(_826__bF_buf3), .B(_1028_), .Y(_1029_) );
NAND2X1 NAND2X1_201 ( .A(_1027_), .B(_1029_), .Y(_1030_) );
INVX1 INVX1_144 ( .A(_1030_), .Y(_1031_) );
NOR2X1 NOR2X1_329 ( .A(_1027_), .B(_1029_), .Y(_1032_) );
OAI21X1 OAI21X1_287 ( .A(_1031_), .B(_1032_), .C(micro_hash_ucr_pipe50_bF_buf0), .Y(_1033_) );
OAI21X1 OAI21X1_288 ( .A(_1026_), .B(micro_hash_ucr_pipe50_bF_buf0), .C(_1033_), .Y(_1034_) );
NAND2X1 NAND2X1_202 ( .A(_542_), .B(_744_), .Y(_1035_) );
OAI21X1 OAI21X1_289 ( .A(_743_), .B(_597__bF_buf0), .C(_1035_), .Y(_1036_) );
INVX1 INVX1_145 ( .A(micro_hash_ucr_Wx_178_), .Y(_1037_) );
OAI21X1 OAI21X1_290 ( .A(_824__bF_buf3), .B(_823__bF_buf1), .C(_1037_), .Y(_1038_) );
NOR2X1 NOR2X1_330 ( .A(_1037_), .B(_827__bF_buf5), .Y(_1039_) );
INVX1 INVX1_146 ( .A(_1039_), .Y(_1040_) );
NAND2X1 NAND2X1_203 ( .A(_1038_), .B(_1040_), .Y(_1041_) );
XOR2X1 XOR2X1_13 ( .A(_1041_), .B(_1036_), .Y(_1042_) );
MUX2X1 MUX2X1_41 ( .A(_1034_), .B(_1042_), .S(_4214__bF_buf3), .Y(_1043_) );
OAI21X1 OAI21X1_291 ( .A(_749_), .B(_597__bF_buf2), .C(_751_), .Y(_1044_) );
INVX2 INVX2_77 ( .A(micro_hash_ucr_Wx_186_), .Y(_1045_) );
XNOR2X1 XNOR2X1_47 ( .A(_826__bF_buf3), .B(_1045_), .Y(_1046_) );
NOR2X1 NOR2X1_331 ( .A(_1044_), .B(_1046_), .Y(_1047_) );
NOR2X1 NOR2X1_332 ( .A(_749_), .B(_597__bF_buf2), .Y(_1048_) );
OAI21X1 OAI21X1_292 ( .A(_752_), .B(_1048_), .C(_1046_), .Y(_1049_) );
INVX1 INVX1_147 ( .A(_1049_), .Y(_1050_) );
OAI21X1 OAI21X1_293 ( .A(_1050_), .B(_1047_), .C(micro_hash_ucr_pipe54_bF_buf0), .Y(_1051_) );
OAI21X1 OAI21X1_294 ( .A(_1043_), .B(micro_hash_ucr_pipe54_bF_buf0), .C(_1051_), .Y(_1052_) );
NOR2X1 NOR2X1_333 ( .A(_755_), .B(_597__bF_buf1), .Y(_1053_) );
INVX2 INVX2_78 ( .A(micro_hash_ucr_Wx_194_), .Y(_1054_) );
XNOR2X1 XNOR2X1_48 ( .A(_826__bF_buf1), .B(_1054_), .Y(_1055_) );
OAI21X1 OAI21X1_295 ( .A(_758_), .B(_1053_), .C(_1055_), .Y(_1056_) );
INVX1 INVX1_148 ( .A(_1056_), .Y(_1057_) );
OAI21X1 OAI21X1_296 ( .A(_755_), .B(_597__bF_buf1), .C(_757_), .Y(_1058_) );
NOR2X1 NOR2X1_334 ( .A(_1058_), .B(_1055_), .Y(_1059_) );
OAI21X1 OAI21X1_297 ( .A(_1057_), .B(_1059_), .C(micro_hash_ucr_pipe56_bF_buf1), .Y(_1060_) );
NAND2X1 NAND2X1_204 ( .A(_4211__bF_buf2), .B(_1060_), .Y(_1061_) );
AOI21X1 AOI21X1_99 ( .A(_832__bF_buf3), .B(_1052_), .C(_1061_), .Y(_1062_) );
OAI21X1 OAI21X1_298 ( .A(_762_), .B(_597__bF_buf1), .C(_768_), .Y(_1063_) );
INVX2 INVX2_79 ( .A(micro_hash_ucr_Wx_202_), .Y(_1064_) );
XNOR2X1 XNOR2X1_49 ( .A(_826__bF_buf3), .B(_1064_), .Y(_1065_) );
OAI21X1 OAI21X1_299 ( .A(_1063_), .B(_1065_), .C(micro_hash_ucr_pipe58_bF_buf1), .Y(_1066_) );
AOI21X1 AOI21X1_100 ( .A(_1063_), .B(_1065_), .C(_1066_), .Y(_1067_) );
OAI21X1 OAI21X1_300 ( .A(_1062_), .B(_1067_), .C(_4210__bF_buf2), .Y(_1068_) );
OAI21X1 OAI21X1_301 ( .A(_4210__bF_buf2), .B(_831_), .C(_1068_), .Y(_1069_) );
OAI21X1 OAI21X1_302 ( .A(_780_), .B(_597__bF_buf2), .C(_782_), .Y(_1070_) );
INVX2 INVX2_80 ( .A(micro_hash_ucr_Wx_218_), .Y(_1071_) );
XNOR2X1 XNOR2X1_50 ( .A(_826__bF_buf3), .B(_1071_), .Y(_1072_) );
NOR2X1 NOR2X1_335 ( .A(_1070_), .B(_1072_), .Y(_1073_) );
NAND2X1 NAND2X1_205 ( .A(_1070_), .B(_1072_), .Y(_1074_) );
NAND2X1 NAND2X1_206 ( .A(micro_hash_ucr_pipe62_bF_buf1), .B(_1074_), .Y(_1075_) );
OAI21X1 OAI21X1_303 ( .A(_1075_), .B(_1073_), .C(_278__bF_buf3), .Y(_1076_) );
AOI21X1 AOI21X1_101 ( .A(_4207__bF_buf0), .B(_1069_), .C(_1076_), .Y(_1077_) );
INVX8 INVX8_62 ( .A(micro_hash_ucr_pipe66_bF_buf3), .Y(_1078_) );
NAND2X1 NAND2X1_207 ( .A(_564_), .B(_788_), .Y(_1079_) );
OAI21X1 OAI21X1_304 ( .A(_787_), .B(_597__bF_buf2), .C(_1079_), .Y(_1080_) );
INVX2 INVX2_81 ( .A(micro_hash_ucr_Wx_226_), .Y(_1081_) );
OAI21X1 OAI21X1_305 ( .A(_824__bF_buf1), .B(_823__bF_buf0), .C(_1081_), .Y(_1082_) );
NOR2X1 NOR2X1_336 ( .A(_1081_), .B(_827__bF_buf2), .Y(_1083_) );
INVX1 INVX1_149 ( .A(_1083_), .Y(_1084_) );
NAND2X1 NAND2X1_208 ( .A(_1082_), .B(_1084_), .Y(_1085_) );
XNOR2X1 XNOR2X1_51 ( .A(_1085_), .B(_1080_), .Y(_1086_) );
OAI21X1 OAI21X1_306 ( .A(_1086_), .B(_278__bF_buf3), .C(_1078__bF_buf0), .Y(_1087_) );
INVX2 INVX2_82 ( .A(micro_hash_ucr_Wx_234_), .Y(_1088_) );
XNOR2X1 XNOR2X1_52 ( .A(_826__bF_buf3), .B(_1088_), .Y(_1089_) );
OAI21X1 OAI21X1_307 ( .A(_797_), .B(_794_), .C(_1089_), .Y(_1090_) );
INVX1 INVX1_150 ( .A(_1090_), .Y(_1091_) );
OAI21X1 OAI21X1_308 ( .A(_796_), .B(_570_), .C(_795_), .Y(_1092_) );
OAI21X1 OAI21X1_309 ( .A(_1092_), .B(_1089_), .C(micro_hash_ucr_pipe66_bF_buf1), .Y(_1093_) );
OAI22X1 OAI22X1_21 ( .A(_1091_), .B(_1093_), .C(_1077_), .D(_1087_), .Y(_1094_) );
AOI21X1 AOI21X1_102 ( .A(micro_hash_ucr_Wx_241_), .B(_588__bF_buf4), .C(_803_), .Y(_1095_) );
INVX2 INVX2_83 ( .A(micro_hash_ucr_Wx_242_), .Y(_1096_) );
OAI21X1 OAI21X1_310 ( .A(_824__bF_buf1), .B(_823__bF_buf0), .C(_1096_), .Y(_1097_) );
INVX1 INVX1_151 ( .A(_1097_), .Y(_1098_) );
NOR2X1 NOR2X1_337 ( .A(_1096_), .B(_827__bF_buf1), .Y(_1099_) );
OAI21X1 OAI21X1_311 ( .A(_1099_), .B(_1098_), .C(_1095_), .Y(_1100_) );
NOR3X1 NOR3X1_18 ( .A(_1095_), .B(_1098_), .C(_1099_), .Y(_1101_) );
INVX1 INVX1_152 ( .A(_1101_), .Y(_1102_) );
NAND2X1 NAND2X1_209 ( .A(_1100_), .B(_1102_), .Y(_1103_) );
OAI21X1 OAI21X1_312 ( .A(_1103_), .B(_4199__bF_buf2), .C(_287_), .Y(_1104_) );
AOI21X1 AOI21X1_103 ( .A(_4199__bF_buf2), .B(_1094_), .C(_1104_), .Y(_1105_) );
NOR2X1 NOR2X1_338 ( .A(_808_), .B(_597__bF_buf2), .Y(_1106_) );
NOR2X1 NOR2X1_339 ( .A(_1106_), .B(_810_), .Y(_1107_) );
INVX2 INVX2_84 ( .A(micro_hash_ucr_Wx_250_), .Y(_1108_) );
OAI21X1 OAI21X1_313 ( .A(_824__bF_buf1), .B(_823__bF_buf0), .C(_1108_), .Y(_1109_) );
INVX1 INVX1_153 ( .A(_1109_), .Y(_1110_) );
NOR2X1 NOR2X1_340 ( .A(_1108_), .B(_827__bF_buf1), .Y(_1111_) );
OAI21X1 OAI21X1_314 ( .A(_1111_), .B(_1110_), .C(_1107_), .Y(_1112_) );
NOR2X1 NOR2X1_341 ( .A(_1110_), .B(_1111_), .Y(_1113_) );
OAI21X1 OAI21X1_315 ( .A(_810_), .B(_1106_), .C(_1113_), .Y(_1114_) );
NAND3X1 NAND3X1_79 ( .A(_131__bF_buf3), .B(_1112_), .C(_1114_), .Y(_1115_) );
AOI21X1 AOI21X1_104 ( .A(_345_), .B(_1115_), .C(_1105_), .Y(_128__2_) );
OAI21X1 OAI21X1_316 ( .A(_1096_), .B(_827__bF_buf1), .C(_1102_), .Y(_1116_) );
INVX1 INVX1_154 ( .A(micro_hash_ucr_Wx_243_), .Y(_1117_) );
XOR2X1 XOR2X1_14 ( .A(micro_hash_ucr_k_3_), .B(micro_hash_ucr_x_3_), .Y(_1118_) );
OAI21X1 OAI21X1_317 ( .A(_823__bF_buf3), .B(_820_), .C(_1118_), .Y(_1119_) );
INVX8 INVX8_63 ( .A(_1119_), .Y(_1120_) );
OAI21X1 OAI21X1_318 ( .A(_816_), .B(_822_), .C(_821_), .Y(_1121_) );
NOR2X1 NOR2X1_342 ( .A(_1118_), .B(_1121_), .Y(_1122_) );
OAI21X1 OAI21X1_319 ( .A(_1120__bF_buf1), .B(_1122__bF_buf2), .C(_1117_), .Y(_1123_) );
INVX1 INVX1_155 ( .A(_1123_), .Y(_1124_) );
OR2X2 OR2X2_12 ( .A(_1120__bF_buf0), .B(_1122__bF_buf1), .Y(_1125_) );
NOR2X1 NOR2X1_343 ( .A(_1117_), .B(_1125__bF_buf3), .Y(_1126_) );
OAI21X1 OAI21X1_320 ( .A(_1124_), .B(_1126_), .C(_1116_), .Y(_1127_) );
INVX1 INVX1_156 ( .A(_1116_), .Y(_1128_) );
INVX1 INVX1_157 ( .A(_1126_), .Y(_1129_) );
NAND3X1 NAND3X1_80 ( .A(_1123_), .B(_1129_), .C(_1128_), .Y(_1130_) );
NAND3X1 NAND3X1_81 ( .A(micro_hash_ucr_pipe68), .B(_1127_), .C(_1130_), .Y(_1131_) );
OAI21X1 OAI21X1_321 ( .A(_1071_), .B(_827__bF_buf2), .C(_1074_), .Y(_1132_) );
INVX1 INVX1_158 ( .A(micro_hash_ucr_Wx_219_), .Y(_1133_) );
OAI21X1 OAI21X1_322 ( .A(_1120__bF_buf1), .B(_1122__bF_buf2), .C(_1133_), .Y(_1134_) );
NOR2X1 NOR2X1_344 ( .A(_1133_), .B(_1125__bF_buf3), .Y(_1135_) );
INVX1 INVX1_159 ( .A(_1135_), .Y(_1136_) );
NAND2X1 NAND2X1_210 ( .A(_1134_), .B(_1136_), .Y(_1137_) );
XNOR2X1 XNOR2X1_53 ( .A(_1137_), .B(_1132_), .Y(_1138_) );
OAI21X1 OAI21X1_323 ( .A(_1045_), .B(_827__bF_buf2), .C(_1049_), .Y(_1139_) );
INVX1 INVX1_160 ( .A(micro_hash_ucr_Wx_187_), .Y(_1140_) );
OAI21X1 OAI21X1_324 ( .A(_1120__bF_buf2), .B(_1122__bF_buf0), .C(_1140_), .Y(_1141_) );
NOR2X1 NOR2X1_345 ( .A(_1140_), .B(_1125__bF_buf0), .Y(_1142_) );
INVX1 INVX1_161 ( .A(_1142_), .Y(_1143_) );
NAND2X1 NAND2X1_211 ( .A(_1141_), .B(_1143_), .Y(_1144_) );
XNOR2X1 XNOR2X1_54 ( .A(_1144_), .B(_1139_), .Y(_1145_) );
OAI21X1 OAI21X1_325 ( .A(_1011_), .B(_827__bF_buf5), .C(_1014_), .Y(_1146_) );
INVX1 INVX1_162 ( .A(micro_hash_ucr_Wx_155_), .Y(_1147_) );
OAI21X1 OAI21X1_326 ( .A(_1120__bF_buf3), .B(_1122__bF_buf3), .C(_1147_), .Y(_1148_) );
INVX1 INVX1_163 ( .A(_1148_), .Y(_1149_) );
NOR2X1 NOR2X1_346 ( .A(_1147_), .B(_1125__bF_buf1), .Y(_1150_) );
NOR2X1 NOR2X1_347 ( .A(_1149_), .B(_1150_), .Y(_1151_) );
XOR2X1 XOR2X1_15 ( .A(_1151_), .B(_1146_), .Y(_1152_) );
OAI21X1 OAI21X1_327 ( .A(_971_), .B(_827__bF_buf0), .C(_978_), .Y(_1153_) );
INVX2 INVX2_85 ( .A(micro_hash_ucr_Wx_123_), .Y(_1154_) );
OAI21X1 OAI21X1_328 ( .A(_1120__bF_buf3), .B(_1122__bF_buf3), .C(_1154_), .Y(_1155_) );
NOR2X1 NOR2X1_348 ( .A(_1154_), .B(_1125__bF_buf1), .Y(_1156_) );
INVX1 INVX1_164 ( .A(_1156_), .Y(_1157_) );
NAND2X1 NAND2X1_212 ( .A(_1155_), .B(_1157_), .Y(_1158_) );
XNOR2X1 XNOR2X1_55 ( .A(_1153_), .B(_1158_), .Y(_1159_) );
NOR2X1 NOR2X1_349 ( .A(_671_), .B(_597__bF_buf3), .Y(_1160_) );
OAI21X1 OAI21X1_329 ( .A(_674_), .B(_1160_), .C(_940_), .Y(_1161_) );
OAI21X1 OAI21X1_330 ( .A(_939_), .B(_827__bF_buf4), .C(_1161_), .Y(_1162_) );
INVX2 INVX2_86 ( .A(micro_hash_ucr_Wx_91_), .Y(_1163_) );
OAI21X1 OAI21X1_331 ( .A(_1120__bF_buf2), .B(_1122__bF_buf0), .C(_1163_), .Y(_1164_) );
NOR2X1 NOR2X1_350 ( .A(_1163_), .B(_1125__bF_buf2), .Y(_1165_) );
INVX1 INVX1_165 ( .A(_1165_), .Y(_1166_) );
NAND2X1 NAND2X1_213 ( .A(_1164_), .B(_1166_), .Y(_1167_) );
XNOR2X1 XNOR2X1_56 ( .A(_1167_), .B(_1162_), .Y(_1168_) );
OAI21X1 OAI21X1_332 ( .A(_903_), .B(_827__bF_buf4), .C(_906_), .Y(_1169_) );
INVX2 INVX2_87 ( .A(micro_hash_ucr_Wx_59_), .Y(_1170_) );
OAI21X1 OAI21X1_333 ( .A(_1120__bF_buf0), .B(_1122__bF_buf1), .C(_1170_), .Y(_1171_) );
NOR2X1 NOR2X1_351 ( .A(_1170_), .B(_1125__bF_buf2), .Y(_1172_) );
INVX1 INVX1_166 ( .A(_1172_), .Y(_1173_) );
NAND2X1 NAND2X1_214 ( .A(_1171_), .B(_1173_), .Y(_1174_) );
XNOR2X1 XNOR2X1_57 ( .A(_1174_), .B(_1169_), .Y(_1175_) );
NOR2X1 NOR2X1_352 ( .A(_851_), .B(_853_), .Y(_1176_) );
INVX1 INVX1_167 ( .A(micro_hash_ucr_Wx_3_), .Y(_1177_) );
OAI21X1 OAI21X1_334 ( .A(_1120__bF_buf4), .B(_1122__bF_buf4), .C(_1177_), .Y(_1178_) );
INVX1 INVX1_168 ( .A(_1178_), .Y(_1179_) );
NOR2X1 NOR2X1_353 ( .A(_1177_), .B(_1125__bF_buf4), .Y(_1180_) );
NOR2X1 NOR2X1_354 ( .A(_1179_), .B(_1180_), .Y(_1181_) );
OAI21X1 OAI21X1_335 ( .A(_1176_), .B(_1181_), .C(micro_hash_ucr_pipe8), .Y(_1182_) );
AOI21X1 AOI21X1_105 ( .A(_1176_), .B(_1181_), .C(_1182_), .Y(_1183_) );
INVX1 INVX1_169 ( .A(H_19_), .Y(_1184_) );
NOR2X1 NOR2X1_355 ( .A(_4252_), .B(_1184_), .Y(_1185_) );
OAI21X1 OAI21X1_336 ( .A(_4200_), .B(micro_hash_ucr_pipe6), .C(_438_), .Y(_1186_) );
OAI21X1 OAI21X1_337 ( .A(_1186_), .B(_1185_), .C(_4243_), .Y(_1187_) );
NOR2X1 NOR2X1_356 ( .A(_1187_), .B(_1183_), .Y(_1188_) );
AOI21X1 AOI21X1_106 ( .A(_860_), .B(_858_), .C(_862_), .Y(_1189_) );
INVX1 INVX1_170 ( .A(micro_hash_ucr_Wx_11_), .Y(_1190_) );
OAI21X1 OAI21X1_338 ( .A(_1120__bF_buf4), .B(_1122__bF_buf4), .C(_1190_), .Y(_1191_) );
INVX1 INVX1_171 ( .A(_1191_), .Y(_1192_) );
NOR2X1 NOR2X1_357 ( .A(_1190_), .B(_1125__bF_buf4), .Y(_1193_) );
NOR2X1 NOR2X1_358 ( .A(_1192_), .B(_1193_), .Y(_1194_) );
XOR2X1 XOR2X1_16 ( .A(_1194_), .B(_1189_), .Y(_1195_) );
OAI21X1 OAI21X1_339 ( .A(_1195_), .B(_4243_), .C(_4258_), .Y(_1196_) );
NAND2X1 NAND2X1_215 ( .A(_841_), .B(_843_), .Y(_1197_) );
OAI21X1 OAI21X1_340 ( .A(_842_), .B(_827__bF_buf3), .C(_1197_), .Y(_1198_) );
INVX2 INVX2_88 ( .A(micro_hash_ucr_Wx_19_), .Y(_1199_) );
OAI21X1 OAI21X1_341 ( .A(_1120__bF_buf4), .B(_1122__bF_buf4), .C(_1199_), .Y(_1200_) );
NOR2X1 NOR2X1_359 ( .A(_1199_), .B(_1125__bF_buf4), .Y(_1201_) );
INVX1 INVX1_172 ( .A(_1201_), .Y(_1202_) );
NAND2X1 NAND2X1_216 ( .A(_1200_), .B(_1202_), .Y(_1203_) );
AOI21X1 AOI21X1_107 ( .A(_1198_), .B(_1203_), .C(_4258_), .Y(_1204_) );
OAI21X1 OAI21X1_342 ( .A(_1198_), .B(_1203_), .C(_1204_), .Y(_1205_) );
OAI21X1 OAI21X1_343 ( .A(_1188_), .B(_1196_), .C(_1205_), .Y(_1206_) );
NAND2X1 NAND2X1_217 ( .A(_4241__bF_buf1), .B(_1206_), .Y(_1207_) );
OAI21X1 OAI21X1_344 ( .A(_870_), .B(_827__bF_buf3), .C(_877_), .Y(_1208_) );
INVX2 INVX2_89 ( .A(micro_hash_ucr_Wx_27_), .Y(_1209_) );
OAI21X1 OAI21X1_345 ( .A(_1120__bF_buf4), .B(_1122__bF_buf4), .C(_1209_), .Y(_1210_) );
NOR2X1 NOR2X1_360 ( .A(_1209_), .B(_1125__bF_buf4), .Y(_1211_) );
INVX1 INVX1_173 ( .A(_1211_), .Y(_1212_) );
NAND2X1 NAND2X1_218 ( .A(_1210_), .B(_1212_), .Y(_1213_) );
XNOR2X1 XNOR2X1_58 ( .A(_1208_), .B(_1213_), .Y(_1214_) );
OAI21X1 OAI21X1_346 ( .A(_4241__bF_buf1), .B(_1214_), .C(_1207_), .Y(_1215_) );
NAND3X1 NAND3X1_82 ( .A(_834_), .B(_836_), .C(_838_), .Y(_1216_) );
OAI21X1 OAI21X1_347 ( .A(_835_), .B(_827__bF_buf3), .C(_1216_), .Y(_1217_) );
INVX2 INVX2_90 ( .A(micro_hash_ucr_Wx_35_), .Y(_1218_) );
OAI21X1 OAI21X1_348 ( .A(_1120__bF_buf4), .B(_1122__bF_buf4), .C(_1218_), .Y(_1219_) );
NOR2X1 NOR2X1_361 ( .A(_1218_), .B(_1125__bF_buf4), .Y(_1220_) );
INVX1 INVX1_174 ( .A(_1220_), .Y(_1221_) );
NAND2X1 NAND2X1_219 ( .A(_1219_), .B(_1221_), .Y(_1222_) );
AOI21X1 AOI21X1_108 ( .A(_1217_), .B(_1222_), .C(_4239__bF_buf2), .Y(_1223_) );
OAI21X1 OAI21X1_349 ( .A(_1217_), .B(_1222_), .C(_1223_), .Y(_1224_) );
NAND2X1 NAND2X1_220 ( .A(_624__bF_buf0), .B(_1224_), .Y(_1225_) );
AOI21X1 AOI21X1_109 ( .A(_4239__bF_buf2), .B(_1215_), .C(_1225_), .Y(_1226_) );
NAND3X1 NAND3X1_83 ( .A(_883_), .B(_885_), .C(_887_), .Y(_1227_) );
OAI21X1 OAI21X1_350 ( .A(_884_), .B(_827__bF_buf3), .C(_1227_), .Y(_1228_) );
INVX2 INVX2_91 ( .A(micro_hash_ucr_Wx_43_), .Y(_1229_) );
OAI21X1 OAI21X1_351 ( .A(_1120__bF_buf0), .B(_1122__bF_buf4), .C(_1229_), .Y(_1230_) );
NOR2X1 NOR2X1_362 ( .A(_1229_), .B(_1125__bF_buf4), .Y(_1231_) );
INVX1 INVX1_175 ( .A(_1231_), .Y(_1232_) );
NAND2X1 NAND2X1_221 ( .A(_1230_), .B(_1232_), .Y(_1233_) );
XOR2X1 XOR2X1_17 ( .A(_1233_), .B(_1228_), .Y(_1234_) );
OAI21X1 OAI21X1_352 ( .A(_1234_), .B(_624__bF_buf0), .C(_4237__bF_buf1), .Y(_1235_) );
OAI21X1 OAI21X1_353 ( .A(_891_), .B(_827__bF_buf3), .C(_893_), .Y(_1236_) );
INVX2 INVX2_92 ( .A(micro_hash_ucr_Wx_51_), .Y(_1237_) );
OAI21X1 OAI21X1_354 ( .A(_1120__bF_buf4), .B(_1122__bF_buf4), .C(_1237_), .Y(_1238_) );
NOR2X1 NOR2X1_363 ( .A(_1237_), .B(_1125__bF_buf4), .Y(_1239_) );
INVX1 INVX1_176 ( .A(_1239_), .Y(_1240_) );
NAND2X1 NAND2X1_222 ( .A(_1238_), .B(_1240_), .Y(_1241_) );
AOI21X1 AOI21X1_110 ( .A(_1236_), .B(_1241_), .C(_4237__bF_buf1), .Y(_1242_) );
OAI21X1 OAI21X1_355 ( .A(_1236_), .B(_1241_), .C(_1242_), .Y(_1243_) );
OAI21X1 OAI21X1_356 ( .A(_1226_), .B(_1235_), .C(_1243_), .Y(_1244_) );
NAND2X1 NAND2X1_223 ( .A(_4262__bF_buf3), .B(_1244_), .Y(_1245_) );
OAI21X1 OAI21X1_357 ( .A(_4262__bF_buf3), .B(_1175_), .C(_1245_), .Y(_1246_) );
NAND3X1 NAND3X1_84 ( .A(_910_), .B(_912_), .C(_914_), .Y(_1247_) );
OAI21X1 OAI21X1_358 ( .A(_911_), .B(_827__bF_buf4), .C(_1247_), .Y(_1248_) );
INVX2 INVX2_93 ( .A(micro_hash_ucr_Wx_67_), .Y(_1249_) );
OAI21X1 OAI21X1_359 ( .A(_1120__bF_buf0), .B(_1122__bF_buf1), .C(_1249_), .Y(_1250_) );
NOR2X1 NOR2X1_364 ( .A(_1249_), .B(_1125__bF_buf2), .Y(_1251_) );
INVX1 INVX1_177 ( .A(_1251_), .Y(_1252_) );
NAND2X1 NAND2X1_224 ( .A(_1250_), .B(_1252_), .Y(_1253_) );
AOI21X1 AOI21X1_111 ( .A(_1248_), .B(_1253_), .C(_4233__bF_buf0), .Y(_1254_) );
OAI21X1 OAI21X1_360 ( .A(_1248_), .B(_1253_), .C(_1254_), .Y(_1255_) );
NAND2X1 NAND2X1_225 ( .A(_4230__bF_buf4), .B(_1255_), .Y(_1256_) );
AOI21X1 AOI21X1_112 ( .A(_4233__bF_buf0), .B(_1246_), .C(_1256_), .Y(_1257_) );
NOR2X1 NOR2X1_365 ( .A(_924_), .B(_926_), .Y(_1258_) );
INVX2 INVX2_94 ( .A(micro_hash_ucr_Wx_75_), .Y(_1259_) );
OAI21X1 OAI21X1_361 ( .A(_1120__bF_buf0), .B(_1122__bF_buf1), .C(_1259_), .Y(_1260_) );
NOR2X1 NOR2X1_366 ( .A(_1259_), .B(_1125__bF_buf2), .Y(_1261_) );
INVX1 INVX1_178 ( .A(_1261_), .Y(_1262_) );
NAND2X1 NAND2X1_226 ( .A(_1260_), .B(_1262_), .Y(_1263_) );
AND2X2 AND2X2_44 ( .A(_1258_), .B(_1263_), .Y(_1264_) );
OAI21X1 OAI21X1_362 ( .A(_1258_), .B(_1263_), .C(micro_hash_ucr_pipe26_bF_buf0), .Y(_1265_) );
OAI21X1 OAI21X1_363 ( .A(_1264_), .B(_1265_), .C(_220__bF_buf0), .Y(_1266_) );
NAND3X1 NAND3X1_85 ( .A(_930_), .B(_932_), .C(_934_), .Y(_1267_) );
OAI21X1 OAI21X1_364 ( .A(_931_), .B(_827__bF_buf0), .C(_1267_), .Y(_1268_) );
INVX2 INVX2_95 ( .A(micro_hash_ucr_Wx_83_), .Y(_1269_) );
OAI21X1 OAI21X1_365 ( .A(_1120__bF_buf2), .B(_1122__bF_buf1), .C(_1269_), .Y(_1270_) );
NOR2X1 NOR2X1_367 ( .A(_1269_), .B(_1125__bF_buf2), .Y(_1271_) );
INVX1 INVX1_179 ( .A(_1271_), .Y(_1272_) );
NAND2X1 NAND2X1_227 ( .A(_1270_), .B(_1272_), .Y(_1273_) );
AOI21X1 AOI21X1_113 ( .A(_1268_), .B(_1273_), .C(_220__bF_buf0), .Y(_1274_) );
OAI21X1 OAI21X1_366 ( .A(_1268_), .B(_1273_), .C(_1274_), .Y(_1275_) );
OAI21X1 OAI21X1_367 ( .A(_1257_), .B(_1266_), .C(_1275_), .Y(_1276_) );
NAND2X1 NAND2X1_228 ( .A(_4228__bF_buf4), .B(_1276_), .Y(_1277_) );
OAI21X1 OAI21X1_368 ( .A(_4228__bF_buf4), .B(_1168_), .C(_1277_), .Y(_1278_) );
OAI21X1 OAI21X1_369 ( .A(_946_), .B(_827__bF_buf4), .C(_948_), .Y(_1279_) );
INVX2 INVX2_96 ( .A(micro_hash_ucr_Wx_99_), .Y(_1280_) );
OAI21X1 OAI21X1_370 ( .A(_1120__bF_buf2), .B(_1122__bF_buf0), .C(_1280_), .Y(_1281_) );
NOR2X1 NOR2X1_368 ( .A(_1280_), .B(_1125__bF_buf0), .Y(_1282_) );
INVX1 INVX1_180 ( .A(_1282_), .Y(_1283_) );
NAND2X1 NAND2X1_229 ( .A(_1281_), .B(_1283_), .Y(_1284_) );
XNOR2X1 XNOR2X1_59 ( .A(_1284_), .B(_1279_), .Y(_1285_) );
OAI21X1 OAI21X1_371 ( .A(_1285_), .B(_4226__bF_buf0), .C(_4225__bF_buf4), .Y(_1286_) );
AOI21X1 AOI21X1_114 ( .A(_4226__bF_buf0), .B(_1278_), .C(_1286_), .Y(_1287_) );
OAI21X1 OAI21X1_372 ( .A(_953_), .B(_827__bF_buf4), .C(_955_), .Y(_1288_) );
INVX2 INVX2_97 ( .A(micro_hash_ucr_Wx_107_), .Y(_1289_) );
OAI21X1 OAI21X1_373 ( .A(_1120__bF_buf0), .B(_1122__bF_buf1), .C(_1289_), .Y(_1290_) );
NOR2X1 NOR2X1_369 ( .A(_1289_), .B(_1125__bF_buf2), .Y(_1291_) );
INVX1 INVX1_181 ( .A(_1291_), .Y(_1292_) );
NAND2X1 NAND2X1_230 ( .A(_1290_), .B(_1292_), .Y(_1293_) );
XOR2X1 XOR2X1_18 ( .A(_1293_), .B(_1288_), .Y(_1294_) );
OAI21X1 OAI21X1_374 ( .A(_1294_), .B(_4225__bF_buf4), .C(_4224__bF_buf4), .Y(_1295_) );
NAND3X1 NAND3X1_86 ( .A(_962_), .B(_964_), .C(_966_), .Y(_1296_) );
OAI21X1 OAI21X1_375 ( .A(_963_), .B(_827__bF_buf0), .C(_1296_), .Y(_1297_) );
INVX2 INVX2_98 ( .A(micro_hash_ucr_Wx_115_), .Y(_1298_) );
OAI21X1 OAI21X1_376 ( .A(_1120__bF_buf3), .B(_1122__bF_buf3), .C(_1298_), .Y(_1299_) );
NOR2X1 NOR2X1_370 ( .A(_1298_), .B(_1125__bF_buf1), .Y(_1300_) );
INVX1 INVX1_182 ( .A(_1300_), .Y(_1301_) );
NAND2X1 NAND2X1_231 ( .A(_1299_), .B(_1301_), .Y(_1302_) );
AOI21X1 AOI21X1_115 ( .A(_1297_), .B(_1302_), .C(_4224__bF_buf4), .Y(_1303_) );
OAI21X1 OAI21X1_377 ( .A(_1297_), .B(_1302_), .C(_1303_), .Y(_1304_) );
OAI21X1 OAI21X1_378 ( .A(_1287_), .B(_1295_), .C(_1304_), .Y(_1305_) );
NAND2X1 NAND2X1_232 ( .A(_701__bF_buf2), .B(_1305_), .Y(_1306_) );
OAI21X1 OAI21X1_379 ( .A(_701__bF_buf2), .B(_1159_), .C(_1306_), .Y(_1307_) );
OAI21X1 OAI21X1_380 ( .A(_983_), .B(_827__bF_buf5), .C(_986_), .Y(_1308_) );
INVX2 INVX2_99 ( .A(micro_hash_ucr_Wx_131_), .Y(_1309_) );
OAI21X1 OAI21X1_381 ( .A(_1120__bF_buf3), .B(_1122__bF_buf3), .C(_1309_), .Y(_1310_) );
NOR2X1 NOR2X1_371 ( .A(_1309_), .B(_1125__bF_buf1), .Y(_1311_) );
INVX1 INVX1_183 ( .A(_1311_), .Y(_1312_) );
NAND2X1 NAND2X1_233 ( .A(_1310_), .B(_1312_), .Y(_1313_) );
XNOR2X1 XNOR2X1_60 ( .A(_1313_), .B(_1308_), .Y(_1314_) );
OAI21X1 OAI21X1_382 ( .A(_1314_), .B(_296__bF_buf2), .C(_4220__bF_buf0), .Y(_1315_) );
AOI21X1 AOI21X1_116 ( .A(_296__bF_buf2), .B(_1307_), .C(_1315_), .Y(_1316_) );
NAND3X1 NAND3X1_87 ( .A(_990_), .B(_992_), .C(_994_), .Y(_1317_) );
OAI21X1 OAI21X1_383 ( .A(_991_), .B(_827__bF_buf0), .C(_1317_), .Y(_1318_) );
INVX2 INVX2_100 ( .A(micro_hash_ucr_Wx_139_), .Y(_1319_) );
OAI21X1 OAI21X1_384 ( .A(_1120__bF_buf3), .B(_1122__bF_buf3), .C(_1319_), .Y(_1320_) );
NOR2X1 NOR2X1_372 ( .A(_1319_), .B(_1125__bF_buf1), .Y(_1321_) );
INVX1 INVX1_184 ( .A(_1321_), .Y(_1322_) );
NAND2X1 NAND2X1_234 ( .A(_1320_), .B(_1322_), .Y(_1323_) );
XOR2X1 XOR2X1_19 ( .A(_1323_), .B(_1318_), .Y(_1324_) );
OAI21X1 OAI21X1_385 ( .A(_1324_), .B(_4220__bF_buf0), .C(_4219__bF_buf2), .Y(_1325_) );
OAI21X1 OAI21X1_386 ( .A(_999_), .B(_827__bF_buf5), .C(_1004_), .Y(_1326_) );
INVX1 INVX1_185 ( .A(micro_hash_ucr_Wx_147_), .Y(_1327_) );
OAI21X1 OAI21X1_387 ( .A(_1120__bF_buf3), .B(_1122__bF_buf3), .C(_1327_), .Y(_1328_) );
NOR2X1 NOR2X1_373 ( .A(_1327_), .B(_1125__bF_buf1), .Y(_1329_) );
INVX1 INVX1_186 ( .A(_1329_), .Y(_1330_) );
NAND2X1 NAND2X1_235 ( .A(_1328_), .B(_1330_), .Y(_1331_) );
AOI21X1 AOI21X1_117 ( .A(_1331_), .B(_1326_), .C(_4219__bF_buf2), .Y(_1332_) );
OAI21X1 OAI21X1_388 ( .A(_1326_), .B(_1331_), .C(_1332_), .Y(_1333_) );
OAI21X1 OAI21X1_389 ( .A(_1316_), .B(_1325_), .C(_1333_), .Y(_1334_) );
NAND2X1 NAND2X1_236 ( .A(_4218__bF_buf1), .B(_1334_), .Y(_1335_) );
OAI21X1 OAI21X1_390 ( .A(_4218__bF_buf1), .B(_1152_), .C(_1335_), .Y(_1336_) );
NAND3X1 NAND3X1_88 ( .A(_1019_), .B(_1021_), .C(_1023_), .Y(_1337_) );
OAI21X1 OAI21X1_391 ( .A(_1020_), .B(_827__bF_buf5), .C(_1337_), .Y(_1338_) );
INVX1 INVX1_187 ( .A(micro_hash_ucr_Wx_163_), .Y(_1339_) );
OAI21X1 OAI21X1_392 ( .A(_1120__bF_buf2), .B(_1122__bF_buf0), .C(_1339_), .Y(_1340_) );
NOR2X1 NOR2X1_374 ( .A(_1339_), .B(_1125__bF_buf0), .Y(_1341_) );
INVX1 INVX1_188 ( .A(_1341_), .Y(_1342_) );
NAND2X1 NAND2X1_237 ( .A(_1340_), .B(_1342_), .Y(_1343_) );
AOI21X1 AOI21X1_118 ( .A(_1338_), .B(_1343_), .C(_4217__bF_buf1), .Y(_1344_) );
OAI21X1 OAI21X1_393 ( .A(_1338_), .B(_1343_), .C(_1344_), .Y(_1345_) );
NAND2X1 NAND2X1_238 ( .A(_4215__bF_buf4), .B(_1345_), .Y(_1346_) );
AOI21X1 AOI21X1_119 ( .A(_4217__bF_buf1), .B(_1336_), .C(_1346_), .Y(_1347_) );
OAI21X1 OAI21X1_394 ( .A(_1028_), .B(_827__bF_buf1), .C(_1030_), .Y(_1348_) );
INVX1 INVX1_189 ( .A(micro_hash_ucr_Wx_171_), .Y(_1349_) );
OAI21X1 OAI21X1_395 ( .A(_1120__bF_buf1), .B(_1122__bF_buf2), .C(_1349_), .Y(_1350_) );
NOR2X1 NOR2X1_375 ( .A(_1349_), .B(_1125__bF_buf3), .Y(_1351_) );
INVX1 INVX1_190 ( .A(_1351_), .Y(_1352_) );
AOI21X1 AOI21X1_120 ( .A(_1350_), .B(_1352_), .C(_1348_), .Y(_1353_) );
INVX1 INVX1_191 ( .A(_1348_), .Y(_1354_) );
NAND2X1 NAND2X1_239 ( .A(_1350_), .B(_1352_), .Y(_1355_) );
OAI21X1 OAI21X1_396 ( .A(_1355_), .B(_1354_), .C(micro_hash_ucr_pipe50_bF_buf2), .Y(_1356_) );
OAI21X1 OAI21X1_397 ( .A(_1356_), .B(_1353_), .C(_4214__bF_buf3), .Y(_1357_) );
AOI21X1 AOI21X1_121 ( .A(micro_hash_ucr_Wx_177_), .B(_588__bF_buf2), .C(_745_), .Y(_1358_) );
OAI21X1 OAI21X1_398 ( .A(_1358_), .B(_1041_), .C(_1040_), .Y(_1359_) );
INVX1 INVX1_192 ( .A(micro_hash_ucr_Wx_179_), .Y(_1360_) );
OAI21X1 OAI21X1_399 ( .A(_1120__bF_buf3), .B(_1122__bF_buf3), .C(_1360_), .Y(_1361_) );
NOR2X1 NOR2X1_376 ( .A(_1360_), .B(_1125__bF_buf0), .Y(_1362_) );
INVX1 INVX1_193 ( .A(_1362_), .Y(_1363_) );
NAND2X1 NAND2X1_240 ( .A(_1361_), .B(_1363_), .Y(_1364_) );
AOI21X1 AOI21X1_122 ( .A(_1359_), .B(_1364_), .C(_4214__bF_buf3), .Y(_1365_) );
OAI21X1 OAI21X1_400 ( .A(_1359_), .B(_1364_), .C(_1365_), .Y(_1366_) );
OAI21X1 OAI21X1_401 ( .A(_1347_), .B(_1357_), .C(_1366_), .Y(_1367_) );
NAND2X1 NAND2X1_241 ( .A(_742__bF_buf3), .B(_1367_), .Y(_1368_) );
OAI21X1 OAI21X1_402 ( .A(_742__bF_buf3), .B(_1145_), .C(_1368_), .Y(_1369_) );
OAI21X1 OAI21X1_403 ( .A(_1054_), .B(_827__bF_buf2), .C(_1056_), .Y(_1370_) );
INVX1 INVX1_194 ( .A(micro_hash_ucr_Wx_195_), .Y(_1371_) );
OAI21X1 OAI21X1_404 ( .A(_1120__bF_buf2), .B(_1122__bF_buf0), .C(_1371_), .Y(_1372_) );
NOR2X1 NOR2X1_377 ( .A(_1371_), .B(_1125__bF_buf0), .Y(_1373_) );
INVX1 INVX1_195 ( .A(_1373_), .Y(_1374_) );
NAND2X1 NAND2X1_242 ( .A(_1372_), .B(_1374_), .Y(_1375_) );
XNOR2X1 XNOR2X1_61 ( .A(_1375_), .B(_1370_), .Y(_1376_) );
OAI21X1 OAI21X1_405 ( .A(_1376_), .B(_832__bF_buf3), .C(_4211__bF_buf3), .Y(_1377_) );
AOI21X1 AOI21X1_123 ( .A(_832__bF_buf3), .B(_1369_), .C(_1377_), .Y(_1378_) );
OAI21X1 OAI21X1_406 ( .A(_769_), .B(_765_), .C(_1065_), .Y(_1379_) );
OAI21X1 OAI21X1_407 ( .A(_1064_), .B(_827__bF_buf2), .C(_1379_), .Y(_1380_) );
INVX1 INVX1_196 ( .A(micro_hash_ucr_Wx_203_), .Y(_1381_) );
OAI21X1 OAI21X1_408 ( .A(_1120__bF_buf1), .B(_1122__bF_buf2), .C(_1381_), .Y(_1382_) );
NOR2X1 NOR2X1_378 ( .A(_1381_), .B(_1125__bF_buf3), .Y(_1383_) );
INVX1 INVX1_197 ( .A(_1383_), .Y(_1384_) );
NAND2X1 NAND2X1_243 ( .A(_1382_), .B(_1384_), .Y(_1385_) );
XOR2X1 XOR2X1_20 ( .A(_1385_), .B(_1380_), .Y(_1386_) );
OAI21X1 OAI21X1_409 ( .A(_1386_), .B(_4211__bF_buf2), .C(_4210__bF_buf2), .Y(_1387_) );
NAND3X1 NAND3X1_89 ( .A(_814_), .B(_825_), .C(_829_), .Y(_1388_) );
OAI21X1 OAI21X1_410 ( .A(_815_), .B(_827__bF_buf2), .C(_1388_), .Y(_1389_) );
INVX1 INVX1_198 ( .A(micro_hash_ucr_Wx_211_), .Y(_1390_) );
OAI21X1 OAI21X1_411 ( .A(_1120__bF_buf1), .B(_1122__bF_buf2), .C(_1390_), .Y(_1391_) );
NOR2X1 NOR2X1_379 ( .A(_1390_), .B(_1125__bF_buf3), .Y(_1392_) );
INVX1 INVX1_199 ( .A(_1392_), .Y(_1393_) );
NAND2X1 NAND2X1_244 ( .A(_1391_), .B(_1393_), .Y(_1394_) );
AOI21X1 AOI21X1_124 ( .A(_1389_), .B(_1394_), .C(_4210__bF_buf2), .Y(_1395_) );
OAI21X1 OAI21X1_412 ( .A(_1389_), .B(_1394_), .C(_1395_), .Y(_1396_) );
OAI21X1 OAI21X1_413 ( .A(_1378_), .B(_1387_), .C(_1396_), .Y(_1397_) );
NAND2X1 NAND2X1_245 ( .A(_4207__bF_buf0), .B(_1397_), .Y(_1398_) );
OAI21X1 OAI21X1_414 ( .A(_4207__bF_buf0), .B(_1138_), .C(_1398_), .Y(_1399_) );
NAND3X1 NAND3X1_90 ( .A(_1080_), .B(_1082_), .C(_1084_), .Y(_1400_) );
OAI21X1 OAI21X1_415 ( .A(_1081_), .B(_827__bF_buf2), .C(_1400_), .Y(_1401_) );
INVX1 INVX1_200 ( .A(micro_hash_ucr_Wx_227_), .Y(_1402_) );
OAI21X1 OAI21X1_416 ( .A(_1120__bF_buf2), .B(_1122__bF_buf0), .C(_1402_), .Y(_1403_) );
NOR2X1 NOR2X1_380 ( .A(_1402_), .B(_1125__bF_buf0), .Y(_1404_) );
INVX1 INVX1_201 ( .A(_1404_), .Y(_1405_) );
NAND2X1 NAND2X1_246 ( .A(_1403_), .B(_1405_), .Y(_1406_) );
XNOR2X1 XNOR2X1_62 ( .A(_1406_), .B(_1401_), .Y(_1407_) );
OAI21X1 OAI21X1_417 ( .A(_1407_), .B(_278__bF_buf3), .C(_1078__bF_buf0), .Y(_1408_) );
AOI21X1 AOI21X1_125 ( .A(_278__bF_buf3), .B(_1399_), .C(_1408_), .Y(_1409_) );
OAI21X1 OAI21X1_418 ( .A(_1088_), .B(_827__bF_buf1), .C(_1090_), .Y(_1410_) );
INVX1 INVX1_202 ( .A(micro_hash_ucr_Wx_235_), .Y(_1411_) );
OAI21X1 OAI21X1_419 ( .A(_1120__bF_buf1), .B(_1122__bF_buf2), .C(_1411_), .Y(_1412_) );
NOR2X1 NOR2X1_381 ( .A(_1411_), .B(_1125__bF_buf3), .Y(_1413_) );
INVX1 INVX1_203 ( .A(_1413_), .Y(_1414_) );
NAND2X1 NAND2X1_247 ( .A(_1412_), .B(_1414_), .Y(_1415_) );
XOR2X1 XOR2X1_21 ( .A(_1415_), .B(_1410_), .Y(_1416_) );
OAI21X1 OAI21X1_420 ( .A(_1416_), .B(_1078__bF_buf0), .C(_4199__bF_buf2), .Y(_1417_) );
OAI21X1 OAI21X1_421 ( .A(_1409_), .B(_1417_), .C(_1131_), .Y(_1418_) );
OAI21X1 OAI21X1_422 ( .A(_1108_), .B(_827__bF_buf1), .C(_1114_), .Y(_1419_) );
INVX1 INVX1_204 ( .A(micro_hash_ucr_Wx_251_), .Y(_1420_) );
OAI21X1 OAI21X1_423 ( .A(_1120__bF_buf1), .B(_1122__bF_buf2), .C(_1420_), .Y(_1421_) );
NOR2X1 NOR2X1_382 ( .A(_1420_), .B(_1125__bF_buf3), .Y(_1422_) );
INVX1 INVX1_205 ( .A(_1422_), .Y(_1423_) );
NAND2X1 NAND2X1_248 ( .A(_1421_), .B(_1423_), .Y(_1424_) );
AOI21X1 AOI21X1_126 ( .A(_1424_), .B(_1419_), .C(_287_), .Y(_1425_) );
OAI21X1 OAI21X1_424 ( .A(_1419_), .B(_1424_), .C(_1425_), .Y(_1426_) );
NAND2X1 NAND2X1_249 ( .A(_131__bF_buf3), .B(_1426_), .Y(_1427_) );
AOI21X1 AOI21X1_127 ( .A(_287_), .B(_1418_), .C(_1427_), .Y(_128__3_) );
AOI21X1 AOI21X1_128 ( .A(micro_hash_ucr_k_3_), .B(micro_hash_ucr_x_3_), .C(_1120__bF_buf4), .Y(_1428_) );
NOR2X1 NOR2X1_383 ( .A(micro_hash_ucr_k_4_), .B(micro_hash_ucr_x_4_), .Y(_1429_) );
INVX1 INVX1_206 ( .A(micro_hash_ucr_k_4_), .Y(_1430_) );
INVX1 INVX1_207 ( .A(micro_hash_ucr_x_4_), .Y(_1431_) );
NOR2X1 NOR2X1_384 ( .A(_1430_), .B(_1431_), .Y(_1432_) );
NOR2X1 NOR2X1_385 ( .A(_1429_), .B(_1432_), .Y(_1433_) );
INVX1 INVX1_208 ( .A(_1433_), .Y(_1434_) );
NOR2X1 NOR2X1_386 ( .A(_1434_), .B(_1428_), .Y(_1435_) );
INVX1 INVX1_209 ( .A(_1435_), .Y(_1436_) );
OAI21X1 OAI21X1_425 ( .A(_1429_), .B(_1432_), .C(_1428_), .Y(_1437_) );
NAND2X1 NAND2X1_250 ( .A(_1437_), .B(_1436_), .Y(_1438_) );
XOR2X1 XOR2X1_22 ( .A(_1438__bF_buf3), .B(micro_hash_ucr_Wx_12_), .Y(_1439_) );
INVX1 INVX1_210 ( .A(_1193_), .Y(_1440_) );
OAI21X1 OAI21X1_426 ( .A(_1189_), .B(_1192_), .C(_1440_), .Y(_1441_) );
XNOR2X1 XNOR2X1_63 ( .A(_1439_), .B(_1441_), .Y(_1442_) );
XOR2X1 XOR2X1_23 ( .A(_1438__bF_buf3), .B(micro_hash_ucr_Wx_4_), .Y(_1443_) );
INVX1 INVX1_211 ( .A(_1176_), .Y(_1444_) );
AOI21X1 AOI21X1_129 ( .A(_1178_), .B(_1444_), .C(_1180_), .Y(_1445_) );
OAI21X1 OAI21X1_427 ( .A(_1445_), .B(_1443_), .C(micro_hash_ucr_pipe8), .Y(_1446_) );
AOI21X1 AOI21X1_130 ( .A(_1443_), .B(_1445_), .C(_1446_), .Y(_1447_) );
MUX2X1 MUX2X1_42 ( .A(H_20_), .B(micro_hash_ucr_c_4_), .S(micro_hash_ucr_pipe6), .Y(_1448_) );
OAI21X1 OAI21X1_428 ( .A(_1448_), .B(micro_hash_ucr_pipe8), .C(_4243_), .Y(_1449_) );
OAI22X1 OAI22X1_22 ( .A(_4243_), .B(_1442_), .C(_1447_), .D(_1449_), .Y(_1450_) );
INVX2 INVX2_101 ( .A(micro_hash_ucr_Wx_20_), .Y(_1451_) );
XNOR2X1 XNOR2X1_64 ( .A(_1438__bF_buf3), .B(_1451_), .Y(_1452_) );
AOI21X1 AOI21X1_131 ( .A(_1200_), .B(_1198_), .C(_1201_), .Y(_1453_) );
NOR2X1 NOR2X1_387 ( .A(_1453_), .B(_1452_), .Y(_1454_) );
INVX1 INVX1_212 ( .A(_1454_), .Y(_1455_) );
NAND2X1 NAND2X1_251 ( .A(_1453_), .B(_1452_), .Y(_1456_) );
NAND3X1 NAND3X1_91 ( .A(micro_hash_ucr_pipe12_bF_buf2), .B(_1456_), .C(_1455_), .Y(_1457_) );
OAI21X1 OAI21X1_429 ( .A(_1450_), .B(micro_hash_ucr_pipe12_bF_buf2), .C(_1457_), .Y(_1458_) );
XNOR2X1 XNOR2X1_65 ( .A(_1438__bF_buf3), .B(micro_hash_ucr_Wx_28_), .Y(_1459_) );
AOI21X1 AOI21X1_132 ( .A(_1210_), .B(_1208_), .C(_1211_), .Y(_1460_) );
XNOR2X1 XNOR2X1_66 ( .A(_1460_), .B(_1459_), .Y(_1461_) );
MUX2X1 MUX2X1_43 ( .A(_1458_), .B(_1461_), .S(_4241__bF_buf1), .Y(_1462_) );
XNOR2X1 XNOR2X1_67 ( .A(_1438__bF_buf5), .B(micro_hash_ucr_Wx_36_), .Y(_1463_) );
INVX1 INVX1_213 ( .A(_1463_), .Y(_1464_) );
AOI21X1 AOI21X1_133 ( .A(_1219_), .B(_1217_), .C(_1220_), .Y(_1465_) );
NOR2X1 NOR2X1_388 ( .A(_1465_), .B(_1464_), .Y(_1466_) );
INVX1 INVX1_214 ( .A(_1466_), .Y(_1467_) );
NAND2X1 NAND2X1_252 ( .A(_1465_), .B(_1464_), .Y(_1468_) );
AND2X2 AND2X2_45 ( .A(_1467_), .B(_1468_), .Y(_1469_) );
AOI21X1 AOI21X1_134 ( .A(micro_hash_ucr_pipe16), .B(_1469_), .C(micro_hash_ucr_pipe18_bF_buf3), .Y(_1470_) );
OAI21X1 OAI21X1_430 ( .A(_1462_), .B(micro_hash_ucr_pipe16), .C(_1470_), .Y(_1471_) );
XNOR2X1 XNOR2X1_68 ( .A(_1438__bF_buf3), .B(micro_hash_ucr_Wx_44_), .Y(_1472_) );
INVX1 INVX1_215 ( .A(_1472_), .Y(_1473_) );
AOI21X1 AOI21X1_135 ( .A(_1230_), .B(_1228_), .C(_1231_), .Y(_1474_) );
AND2X2 AND2X2_46 ( .A(_1473_), .B(_1474_), .Y(_1475_) );
NOR2X1 NOR2X1_389 ( .A(_1474_), .B(_1473_), .Y(_1476_) );
OAI21X1 OAI21X1_431 ( .A(_1475_), .B(_1476_), .C(micro_hash_ucr_pipe18_bF_buf3), .Y(_1477_) );
NAND3X1 NAND3X1_92 ( .A(_4237__bF_buf1), .B(_1477_), .C(_1471_), .Y(_1478_) );
XNOR2X1 XNOR2X1_69 ( .A(_1438__bF_buf5), .B(micro_hash_ucr_Wx_52_), .Y(_1479_) );
INVX1 INVX1_216 ( .A(_1479_), .Y(_1480_) );
AOI21X1 AOI21X1_136 ( .A(_1238_), .B(_1236_), .C(_1239_), .Y(_1481_) );
NOR2X1 NOR2X1_390 ( .A(_1481_), .B(_1480_), .Y(_1482_) );
INVX1 INVX1_217 ( .A(_1482_), .Y(_1483_) );
NAND2X1 NAND2X1_253 ( .A(_1481_), .B(_1480_), .Y(_1484_) );
NAND2X1 NAND2X1_254 ( .A(_1484_), .B(_1483_), .Y(_1485_) );
OAI21X1 OAI21X1_432 ( .A(_4237__bF_buf1), .B(_1485_), .C(_1478_), .Y(_1486_) );
NOR2X1 NOR2X1_391 ( .A(micro_hash_ucr_pipe22_bF_buf1), .B(_1486_), .Y(_1487_) );
XNOR2X1 XNOR2X1_70 ( .A(_1438__bF_buf5), .B(micro_hash_ucr_Wx_60_), .Y(_1488_) );
INVX1 INVX1_218 ( .A(_1488_), .Y(_1489_) );
AOI21X1 AOI21X1_137 ( .A(_1171_), .B(_1169_), .C(_1172_), .Y(_1490_) );
NAND2X1 NAND2X1_255 ( .A(_1490_), .B(_1489_), .Y(_1491_) );
NOR2X1 NOR2X1_392 ( .A(_1490_), .B(_1489_), .Y(_1492_) );
INVX1 INVX1_219 ( .A(_1492_), .Y(_1493_) );
AOI21X1 AOI21X1_138 ( .A(_1491_), .B(_1493_), .C(_4262__bF_buf3), .Y(_1494_) );
OAI21X1 OAI21X1_433 ( .A(_1487_), .B(_1494_), .C(_4233__bF_buf0), .Y(_1495_) );
XNOR2X1 XNOR2X1_71 ( .A(_1438__bF_buf0), .B(micro_hash_ucr_Wx_68_), .Y(_1496_) );
INVX1 INVX1_220 ( .A(_1496_), .Y(_1497_) );
AOI21X1 AOI21X1_139 ( .A(_1250_), .B(_1248_), .C(_1251_), .Y(_1498_) );
AND2X2 AND2X2_47 ( .A(_1497_), .B(_1498_), .Y(_1499_) );
NOR2X1 NOR2X1_393 ( .A(_1498_), .B(_1497_), .Y(_1500_) );
OAI21X1 OAI21X1_434 ( .A(_1499_), .B(_1500_), .C(micro_hash_ucr_pipe24_bF_buf1), .Y(_1501_) );
NAND3X1 NAND3X1_93 ( .A(_4230__bF_buf4), .B(_1501_), .C(_1495_), .Y(_1502_) );
XNOR2X1 XNOR2X1_72 ( .A(_1438__bF_buf2), .B(micro_hash_ucr_Wx_76_), .Y(_1503_) );
INVX1 INVX1_221 ( .A(_1260_), .Y(_1504_) );
OAI21X1 OAI21X1_435 ( .A(_1258_), .B(_1504_), .C(_1262_), .Y(_1505_) );
AND2X2 AND2X2_48 ( .A(_1503_), .B(_1505_), .Y(_1506_) );
OAI21X1 OAI21X1_436 ( .A(_1503_), .B(_1505_), .C(micro_hash_ucr_pipe26_bF_buf0), .Y(_1507_) );
OAI21X1 OAI21X1_437 ( .A(_1506_), .B(_1507_), .C(_1502_), .Y(_1508_) );
NOR2X1 NOR2X1_394 ( .A(micro_hash_ucr_pipe28_bF_buf3), .B(_1508_), .Y(_1509_) );
XNOR2X1 XNOR2X1_73 ( .A(_1438__bF_buf5), .B(micro_hash_ucr_Wx_84_), .Y(_1510_) );
INVX1 INVX1_222 ( .A(_1510_), .Y(_1511_) );
AOI21X1 AOI21X1_140 ( .A(_1270_), .B(_1268_), .C(_1271_), .Y(_1512_) );
NAND2X1 NAND2X1_256 ( .A(_1512_), .B(_1511_), .Y(_1513_) );
NOR2X1 NOR2X1_395 ( .A(_1512_), .B(_1511_), .Y(_1514_) );
INVX1 INVX1_223 ( .A(_1514_), .Y(_1515_) );
AOI21X1 AOI21X1_141 ( .A(_1513_), .B(_1515_), .C(_220__bF_buf0), .Y(_1516_) );
OAI21X1 OAI21X1_438 ( .A(_1509_), .B(_1516_), .C(_4228__bF_buf4), .Y(_1517_) );
XNOR2X1 XNOR2X1_74 ( .A(_1438__bF_buf2), .B(micro_hash_ucr_Wx_92_), .Y(_1518_) );
INVX1 INVX1_224 ( .A(_1518_), .Y(_1519_) );
AOI21X1 AOI21X1_142 ( .A(_1164_), .B(_1162_), .C(_1165_), .Y(_1520_) );
AND2X2 AND2X2_49 ( .A(_1519_), .B(_1520_), .Y(_1521_) );
NOR2X1 NOR2X1_396 ( .A(_1520_), .B(_1519_), .Y(_1522_) );
OAI21X1 OAI21X1_439 ( .A(_1521_), .B(_1522_), .C(micro_hash_ucr_pipe30_bF_buf2), .Y(_1523_) );
NAND3X1 NAND3X1_94 ( .A(_4226__bF_buf0), .B(_1523_), .C(_1517_), .Y(_1524_) );
INVX2 INVX2_102 ( .A(micro_hash_ucr_Wx_100_), .Y(_1525_) );
XNOR2X1 XNOR2X1_75 ( .A(_1438__bF_buf2), .B(_1525_), .Y(_1526_) );
AOI21X1 AOI21X1_143 ( .A(_1281_), .B(_1279_), .C(_1282_), .Y(_1527_) );
NOR2X1 NOR2X1_397 ( .A(_1527_), .B(_1526_), .Y(_1528_) );
NAND2X1 NAND2X1_257 ( .A(_1527_), .B(_1526_), .Y(_1529_) );
NAND2X1 NAND2X1_258 ( .A(micro_hash_ucr_pipe32_bF_buf3), .B(_1529_), .Y(_1530_) );
OAI21X1 OAI21X1_440 ( .A(_1528_), .B(_1530_), .C(_1524_), .Y(_1531_) );
INVX4 INVX4_25 ( .A(micro_hash_ucr_Wx_108_), .Y(_1532_) );
XNOR2X1 XNOR2X1_76 ( .A(_1438__bF_buf0), .B(_1532_), .Y(_1533_) );
AOI21X1 AOI21X1_144 ( .A(_1290_), .B(_1288_), .C(_1291_), .Y(_1534_) );
AND2X2 AND2X2_50 ( .A(_1533_), .B(_1534_), .Y(_1535_) );
NOR2X1 NOR2X1_398 ( .A(_1534_), .B(_1533_), .Y(_1536_) );
OAI21X1 OAI21X1_441 ( .A(_1535_), .B(_1536_), .C(micro_hash_ucr_pipe34_bF_buf0), .Y(_1537_) );
OAI21X1 OAI21X1_442 ( .A(_1531_), .B(micro_hash_ucr_pipe34_bF_buf0), .C(_1537_), .Y(_1538_) );
NOR2X1 NOR2X1_399 ( .A(micro_hash_ucr_pipe36_bF_buf1), .B(_1538_), .Y(_1539_) );
XNOR2X1 XNOR2X1_77 ( .A(_1438__bF_buf2), .B(micro_hash_ucr_Wx_116_), .Y(_1540_) );
INVX1 INVX1_225 ( .A(_1540_), .Y(_1541_) );
AOI21X1 AOI21X1_145 ( .A(_1299_), .B(_1297_), .C(_1300_), .Y(_1542_) );
NOR2X1 NOR2X1_400 ( .A(_1542_), .B(_1541_), .Y(_1543_) );
INVX1 INVX1_226 ( .A(_1543_), .Y(_1544_) );
AOI21X1 AOI21X1_146 ( .A(_1542_), .B(_1541_), .C(_4224__bF_buf4), .Y(_1545_) );
AOI21X1 AOI21X1_147 ( .A(_1544_), .B(_1545_), .C(_1539_), .Y(_1546_) );
XNOR2X1 XNOR2X1_78 ( .A(_1438__bF_buf2), .B(micro_hash_ucr_Wx_124_), .Y(_1547_) );
INVX1 INVX1_227 ( .A(_1547_), .Y(_1548_) );
AOI21X1 AOI21X1_148 ( .A(_1155_), .B(_1153_), .C(_1156_), .Y(_1549_) );
NAND2X1 NAND2X1_259 ( .A(_1548_), .B(_1549_), .Y(_1550_) );
NOR2X1 NOR2X1_401 ( .A(_1548_), .B(_1549_), .Y(_1551_) );
INVX1 INVX1_228 ( .A(_1551_), .Y(_1552_) );
NAND3X1 NAND3X1_95 ( .A(micro_hash_ucr_pipe38_bF_buf3), .B(_1550_), .C(_1552_), .Y(_1553_) );
OAI21X1 OAI21X1_443 ( .A(_1546_), .B(micro_hash_ucr_pipe38_bF_buf3), .C(_1553_), .Y(_1554_) );
INVX4 INVX4_26 ( .A(micro_hash_ucr_Wx_132_), .Y(_1555_) );
XNOR2X1 XNOR2X1_79 ( .A(_1438__bF_buf0), .B(_1555_), .Y(_1556_) );
AOI21X1 AOI21X1_149 ( .A(_1310_), .B(_1308_), .C(_1311_), .Y(_1557_) );
NOR2X1 NOR2X1_402 ( .A(_1557_), .B(_1556_), .Y(_1558_) );
AND2X2 AND2X2_51 ( .A(_1556_), .B(_1557_), .Y(_1559_) );
OAI21X1 OAI21X1_444 ( .A(_1559_), .B(_1558_), .C(micro_hash_ucr_pipe40_bF_buf4), .Y(_1560_) );
OAI21X1 OAI21X1_445 ( .A(_1554_), .B(micro_hash_ucr_pipe40_bF_buf4), .C(_1560_), .Y(_1561_) );
NAND2X1 NAND2X1_260 ( .A(_4220__bF_buf4), .B(_1561_), .Y(_1562_) );
INVX4 INVX4_27 ( .A(micro_hash_ucr_Wx_140_), .Y(_1563_) );
XNOR2X1 XNOR2X1_80 ( .A(_1438__bF_buf4), .B(_1563_), .Y(_1564_) );
AOI21X1 AOI21X1_150 ( .A(_1320_), .B(_1318_), .C(_1321_), .Y(_1565_) );
AND2X2 AND2X2_52 ( .A(_1564_), .B(_1565_), .Y(_1566_) );
NOR2X1 NOR2X1_403 ( .A(_1565_), .B(_1564_), .Y(_1567_) );
OAI21X1 OAI21X1_446 ( .A(_1566_), .B(_1567_), .C(micro_hash_ucr_pipe42_bF_buf2), .Y(_1568_) );
AOI21X1 AOI21X1_151 ( .A(_1568_), .B(_1562_), .C(micro_hash_ucr_pipe44_bF_buf1), .Y(_1569_) );
XNOR2X1 XNOR2X1_81 ( .A(_1438__bF_buf2), .B(micro_hash_ucr_Wx_148_), .Y(_1570_) );
INVX1 INVX1_229 ( .A(_1570_), .Y(_1571_) );
AOI21X1 AOI21X1_152 ( .A(_1328_), .B(_1326_), .C(_1329_), .Y(_1572_) );
NAND2X1 NAND2X1_261 ( .A(_1572_), .B(_1571_), .Y(_1573_) );
NOR2X1 NOR2X1_404 ( .A(_1572_), .B(_1571_), .Y(_1574_) );
INVX1 INVX1_230 ( .A(_1574_), .Y(_1575_) );
AOI21X1 AOI21X1_153 ( .A(_1573_), .B(_1575_), .C(_4219__bF_buf1), .Y(_1576_) );
OAI21X1 OAI21X1_447 ( .A(_1569_), .B(_1576_), .C(_4218__bF_buf3), .Y(_1577_) );
XNOR2X1 XNOR2X1_82 ( .A(_1438__bF_buf4), .B(micro_hash_ucr_Wx_156_), .Y(_1578_) );
INVX1 INVX1_231 ( .A(_1578_), .Y(_1579_) );
AOI21X1 AOI21X1_154 ( .A(_1148_), .B(_1146_), .C(_1150_), .Y(_1580_) );
AND2X2 AND2X2_53 ( .A(_1579_), .B(_1580_), .Y(_1581_) );
NOR2X1 NOR2X1_405 ( .A(_1580_), .B(_1579_), .Y(_1582_) );
OAI21X1 OAI21X1_448 ( .A(_1581_), .B(_1582_), .C(micro_hash_ucr_pipe46_bF_buf2), .Y(_1583_) );
AOI21X1 AOI21X1_155 ( .A(_1583_), .B(_1577_), .C(micro_hash_ucr_pipe48_bF_buf1), .Y(_1584_) );
XNOR2X1 XNOR2X1_83 ( .A(_1438__bF_buf4), .B(micro_hash_ucr_Wx_164_), .Y(_1585_) );
INVX1 INVX1_232 ( .A(_1585_), .Y(_1586_) );
AOI21X1 AOI21X1_156 ( .A(_1340_), .B(_1338_), .C(_1341_), .Y(_1587_) );
NOR2X1 NOR2X1_406 ( .A(_1587_), .B(_1586_), .Y(_1588_) );
INVX1 INVX1_233 ( .A(_1588_), .Y(_1589_) );
NAND2X1 NAND2X1_262 ( .A(_1587_), .B(_1586_), .Y(_1590_) );
AOI21X1 AOI21X1_157 ( .A(_1590_), .B(_1589_), .C(_4217__bF_buf1), .Y(_1591_) );
OAI21X1 OAI21X1_449 ( .A(_1584_), .B(_1591_), .C(_4215__bF_buf4), .Y(_1592_) );
XOR2X1 XOR2X1_24 ( .A(_1438__bF_buf4), .B(micro_hash_ucr_Wx_172_), .Y(_1593_) );
AOI21X1 AOI21X1_158 ( .A(_1350_), .B(_1348_), .C(_1351_), .Y(_1594_) );
AND2X2 AND2X2_54 ( .A(_1593_), .B(_1594_), .Y(_1595_) );
NOR2X1 NOR2X1_407 ( .A(_1594_), .B(_1593_), .Y(_1596_) );
OAI21X1 OAI21X1_450 ( .A(_1595_), .B(_1596_), .C(micro_hash_ucr_pipe50_bF_buf2), .Y(_1597_) );
NAND2X1 NAND2X1_263 ( .A(_1597_), .B(_1592_), .Y(_1598_) );
XNOR2X1 XNOR2X1_84 ( .A(_1438__bF_buf4), .B(micro_hash_ucr_Wx_180_), .Y(_1599_) );
AOI21X1 AOI21X1_159 ( .A(_1361_), .B(_1359_), .C(_1362_), .Y(_1600_) );
INVX1 INVX1_234 ( .A(_1600_), .Y(_1601_) );
AND2X2 AND2X2_55 ( .A(_1601_), .B(_1599_), .Y(_1602_) );
OAI21X1 OAI21X1_451 ( .A(_1601_), .B(_1599_), .C(micro_hash_ucr_pipe52_bF_buf3), .Y(_1603_) );
OAI22X1 OAI22X1_23 ( .A(_1602_), .B(_1603_), .C(_1598_), .D(micro_hash_ucr_pipe52_bF_buf3), .Y(_1604_) );
XNOR2X1 XNOR2X1_85 ( .A(_1438__bF_buf4), .B(micro_hash_ucr_Wx_188_), .Y(_1605_) );
INVX1 INVX1_235 ( .A(_1605_), .Y(_1606_) );
AOI21X1 AOI21X1_160 ( .A(_1141_), .B(_1139_), .C(_1142_), .Y(_1607_) );
AND2X2 AND2X2_56 ( .A(_1606_), .B(_1607_), .Y(_1608_) );
NOR2X1 NOR2X1_408 ( .A(_1607_), .B(_1606_), .Y(_1609_) );
OAI21X1 OAI21X1_452 ( .A(_1608_), .B(_1609_), .C(micro_hash_ucr_pipe54_bF_buf2), .Y(_1610_) );
OAI21X1 OAI21X1_453 ( .A(_1604_), .B(micro_hash_ucr_pipe54_bF_buf2), .C(_1610_), .Y(_1611_) );
XNOR2X1 XNOR2X1_86 ( .A(_1438__bF_buf1), .B(micro_hash_ucr_Wx_196_), .Y(_1612_) );
INVX1 INVX1_236 ( .A(_1612_), .Y(_1613_) );
AOI21X1 AOI21X1_161 ( .A(_1372_), .B(_1370_), .C(_1373_), .Y(_1614_) );
AND2X2 AND2X2_57 ( .A(_1613_), .B(_1614_), .Y(_1615_) );
NOR2X1 NOR2X1_409 ( .A(_1614_), .B(_1613_), .Y(_1616_) );
OAI21X1 OAI21X1_454 ( .A(_1615_), .B(_1616_), .C(micro_hash_ucr_pipe56_bF_buf3), .Y(_1617_) );
NAND2X1 NAND2X1_264 ( .A(_4211__bF_buf3), .B(_1617_), .Y(_1618_) );
AOI21X1 AOI21X1_162 ( .A(_832__bF_buf3), .B(_1611_), .C(_1618_), .Y(_1619_) );
XOR2X1 XOR2X1_25 ( .A(_1438__bF_buf1), .B(micro_hash_ucr_Wx_204_), .Y(_1620_) );
AOI21X1 AOI21X1_163 ( .A(_1382_), .B(_1380_), .C(_1383_), .Y(_1621_) );
NOR2X1 NOR2X1_410 ( .A(_1621_), .B(_1620_), .Y(_1622_) );
NAND2X1 NAND2X1_265 ( .A(_1621_), .B(_1620_), .Y(_1623_) );
NAND2X1 NAND2X1_266 ( .A(micro_hash_ucr_pipe58_bF_buf1), .B(_1623_), .Y(_1624_) );
OAI21X1 OAI21X1_455 ( .A(_1624_), .B(_1622_), .C(_4210__bF_buf4), .Y(_1625_) );
XNOR2X1 XNOR2X1_87 ( .A(_1438__bF_buf4), .B(micro_hash_ucr_Wx_212_), .Y(_1626_) );
INVX1 INVX1_237 ( .A(_1626_), .Y(_1627_) );
AOI21X1 AOI21X1_164 ( .A(_1391_), .B(_1389_), .C(_1392_), .Y(_1628_) );
AND2X2 AND2X2_58 ( .A(_1627_), .B(_1628_), .Y(_1629_) );
NOR2X1 NOR2X1_411 ( .A(_1628_), .B(_1627_), .Y(_1630_) );
OAI21X1 OAI21X1_456 ( .A(_1629_), .B(_1630_), .C(micro_hash_ucr_pipe60_bF_buf0), .Y(_1631_) );
AND2X2 AND2X2_59 ( .A(_1631_), .B(_4207__bF_buf1), .Y(_1632_) );
OAI21X1 OAI21X1_457 ( .A(_1619_), .B(_1625_), .C(_1632_), .Y(_1633_) );
XNOR2X1 XNOR2X1_88 ( .A(_1438__bF_buf1), .B(micro_hash_ucr_Wx_220_), .Y(_1634_) );
INVX1 INVX1_238 ( .A(_1634_), .Y(_1635_) );
AOI21X1 AOI21X1_165 ( .A(_1134_), .B(_1132_), .C(_1135_), .Y(_1636_) );
NOR2X1 NOR2X1_412 ( .A(_1636_), .B(_1635_), .Y(_1637_) );
INVX1 INVX1_239 ( .A(_1637_), .Y(_1638_) );
AOI21X1 AOI21X1_166 ( .A(_1636_), .B(_1635_), .C(_4207__bF_buf0), .Y(_1639_) );
AOI21X1 AOI21X1_167 ( .A(_1639_), .B(_1638_), .C(micro_hash_ucr_pipe64_bF_buf3), .Y(_1640_) );
XNOR2X1 XNOR2X1_89 ( .A(_1438__bF_buf1), .B(micro_hash_ucr_Wx_228_), .Y(_1641_) );
AOI21X1 AOI21X1_168 ( .A(_1403_), .B(_1401_), .C(_1404_), .Y(_1642_) );
XNOR2X1 XNOR2X1_90 ( .A(_1642_), .B(_1641_), .Y(_1643_) );
OAI21X1 OAI21X1_458 ( .A(_1643_), .B(_278__bF_buf3), .C(_1078__bF_buf0), .Y(_1644_) );
AOI21X1 AOI21X1_169 ( .A(_1640_), .B(_1633_), .C(_1644_), .Y(_1645_) );
XOR2X1 XOR2X1_26 ( .A(_1438__bF_buf1), .B(micro_hash_ucr_Wx_236_), .Y(_1646_) );
AOI21X1 AOI21X1_170 ( .A(_1412_), .B(_1410_), .C(_1413_), .Y(_1647_) );
NOR2X1 NOR2X1_413 ( .A(_1647_), .B(_1646_), .Y(_1648_) );
NAND2X1 NAND2X1_267 ( .A(_1647_), .B(_1646_), .Y(_1649_) );
NAND2X1 NAND2X1_268 ( .A(micro_hash_ucr_pipe66_bF_buf1), .B(_1649_), .Y(_1650_) );
NOR2X1 NOR2X1_414 ( .A(_1648_), .B(_1650_), .Y(_1651_) );
OAI21X1 OAI21X1_459 ( .A(_1645_), .B(_1651_), .C(_4199__bF_buf2), .Y(_1652_) );
XNOR2X1 XNOR2X1_91 ( .A(_1438__bF_buf1), .B(micro_hash_ucr_Wx_244_), .Y(_1653_) );
OAI21X1 OAI21X1_460 ( .A(_1128_), .B(_1124_), .C(_1129_), .Y(_1654_) );
NOR2X1 NOR2X1_415 ( .A(_1653_), .B(_1654_), .Y(_1655_) );
NAND2X1 NAND2X1_269 ( .A(_1653_), .B(_1654_), .Y(_1656_) );
INVX1 INVX1_240 ( .A(_1656_), .Y(_1657_) );
NOR2X1 NOR2X1_416 ( .A(_1655_), .B(_1657_), .Y(_1658_) );
AOI21X1 AOI21X1_171 ( .A(micro_hash_ucr_pipe68), .B(_1658_), .C(micro_hash_ucr_pipe69), .Y(_1659_) );
XNOR2X1 XNOR2X1_92 ( .A(_1438__bF_buf1), .B(micro_hash_ucr_Wx_252_), .Y(_1660_) );
INVX2 INVX2_103 ( .A(_1660_), .Y(_1661_) );
AOI21X1 AOI21X1_172 ( .A(_1421_), .B(_1419_), .C(_1422_), .Y(_1662_) );
AOI21X1 AOI21X1_173 ( .A(_1662_), .B(_1661_), .C(_292__bF_buf6), .Y(_1663_) );
OAI21X1 OAI21X1_461 ( .A(_1661_), .B(_1662_), .C(_1663_), .Y(_1664_) );
AOI22X1 AOI22X1_13 ( .A(_345_), .B(_1664_), .C(_1652_), .D(_1659_), .Y(_128__4_) );
INVX8 INVX8_64 ( .A(_1438__bF_buf3), .Y(_1665_) );
AOI21X1 AOI21X1_174 ( .A(micro_hash_ucr_Wx_244_), .B(_1665__bF_buf3), .C(_1657_), .Y(_1666_) );
INVX1 INVX1_241 ( .A(micro_hash_ucr_Wx_245_), .Y(_1667_) );
NAND2X1 NAND2X1_270 ( .A(_299_), .B(_392_), .Y(_1668_) );
NOR2X1 NOR2X1_417 ( .A(_299_), .B(_392_), .Y(_1669_) );
INVX1 INVX1_242 ( .A(_1669_), .Y(_1670_) );
AND2X2 AND2X2_60 ( .A(_1670_), .B(_1668_), .Y(_1671_) );
OAI21X1 OAI21X1_462 ( .A(_1435_), .B(_1432_), .C(_1671_), .Y(_1672_) );
INVX8 INVX8_65 ( .A(_1672_), .Y(_1673_) );
OAI21X1 OAI21X1_463 ( .A(_1430_), .B(_1431_), .C(_1436_), .Y(_1674_) );
NOR2X1 NOR2X1_418 ( .A(_1671_), .B(_1674_), .Y(_1675_) );
OAI21X1 OAI21X1_464 ( .A(_1675_), .B(_1673__bF_buf3), .C(_1667_), .Y(_1676_) );
INVX1 INVX1_243 ( .A(_1676_), .Y(_1677_) );
NOR2X1 NOR2X1_419 ( .A(_1673__bF_buf3), .B(_1675_), .Y(_1678_) );
INVX8 INVX8_66 ( .A(_1678__bF_buf3), .Y(_1679_) );
NOR2X1 NOR2X1_420 ( .A(_1667_), .B(_1679__bF_buf0), .Y(_1680_) );
NOR2X1 NOR2X1_421 ( .A(_1677_), .B(_1680_), .Y(_1681_) );
AOI21X1 AOI21X1_175 ( .A(_1666_), .B(_1681_), .C(_4199__bF_buf5), .Y(_1682_) );
OAI21X1 OAI21X1_465 ( .A(_1666_), .B(_1681_), .C(_1682_), .Y(_1683_) );
AOI21X1 AOI21X1_176 ( .A(micro_hash_ucr_Wx_220_), .B(_1665__bF_buf2), .C(_1637_), .Y(_1684_) );
NOR2X1 NOR2X1_422 ( .A(micro_hash_ucr_Wx_221_), .B(_1678__bF_buf5), .Y(_1685_) );
INVX1 INVX1_244 ( .A(_1685_), .Y(_1686_) );
NAND2X1 NAND2X1_271 ( .A(micro_hash_ucr_Wx_221_), .B(_1678__bF_buf5), .Y(_1687_) );
NAND2X1 NAND2X1_272 ( .A(_1687_), .B(_1686_), .Y(_1688_) );
XOR2X1 XOR2X1_27 ( .A(_1688_), .B(_1684_), .Y(_1689_) );
AOI21X1 AOI21X1_177 ( .A(micro_hash_ucr_Wx_188_), .B(_1665__bF_buf3), .C(_1609_), .Y(_1690_) );
INVX1 INVX1_245 ( .A(micro_hash_ucr_Wx_189_), .Y(_1691_) );
OAI21X1 OAI21X1_466 ( .A(_1675_), .B(_1673__bF_buf2), .C(_1691_), .Y(_1692_) );
INVX1 INVX1_246 ( .A(_1692_), .Y(_1693_) );
NOR2X1 NOR2X1_423 ( .A(_1691_), .B(_1679__bF_buf1), .Y(_1694_) );
NOR2X1 NOR2X1_424 ( .A(_1693_), .B(_1694_), .Y(_1695_) );
XNOR2X1 XNOR2X1_93 ( .A(_1695_), .B(_1690_), .Y(_1696_) );
AOI21X1 AOI21X1_178 ( .A(micro_hash_ucr_Wx_156_), .B(_1665__bF_buf3), .C(_1582_), .Y(_1697_) );
INVX1 INVX1_247 ( .A(micro_hash_ucr_Wx_157_), .Y(_1698_) );
OAI21X1 OAI21X1_467 ( .A(_1675_), .B(_1673__bF_buf0), .C(_1698_), .Y(_1699_) );
NAND2X1 NAND2X1_273 ( .A(micro_hash_ucr_Wx_157_), .B(_1678__bF_buf1), .Y(_1700_) );
NAND2X1 NAND2X1_274 ( .A(_1699_), .B(_1700_), .Y(_1701_) );
XOR2X1 XOR2X1_28 ( .A(_1697_), .B(_1701_), .Y(_1702_) );
INVX2 INVX2_104 ( .A(micro_hash_ucr_Wx_124_), .Y(_1703_) );
OAI21X1 OAI21X1_468 ( .A(_1703_), .B(_1438__bF_buf0), .C(_1552_), .Y(_1704_) );
INVX2 INVX2_105 ( .A(micro_hash_ucr_Wx_125_), .Y(_1705_) );
OAI21X1 OAI21X1_469 ( .A(_1675_), .B(_1673__bF_buf2), .C(_1705_), .Y(_1706_) );
NOR2X1 NOR2X1_425 ( .A(_1705_), .B(_1679__bF_buf2), .Y(_1707_) );
INVX1 INVX1_248 ( .A(_1707_), .Y(_1708_) );
NAND2X1 NAND2X1_275 ( .A(_1706_), .B(_1708_), .Y(_1709_) );
XNOR2X1 XNOR2X1_94 ( .A(_1704_), .B(_1709_), .Y(_1710_) );
AOI21X1 AOI21X1_179 ( .A(micro_hash_ucr_Wx_92_), .B(_1665__bF_buf0), .C(_1522_), .Y(_1711_) );
INVX2 INVX2_106 ( .A(micro_hash_ucr_Wx_93_), .Y(_1712_) );
OAI21X1 OAI21X1_470 ( .A(_1675_), .B(_1673__bF_buf0), .C(_1712_), .Y(_1713_) );
INVX1 INVX1_249 ( .A(_1713_), .Y(_1714_) );
NOR2X1 NOR2X1_426 ( .A(_1712_), .B(_1679__bF_buf2), .Y(_1715_) );
NOR2X1 NOR2X1_427 ( .A(_1714_), .B(_1715_), .Y(_1716_) );
XNOR2X1 XNOR2X1_95 ( .A(_1716_), .B(_1711_), .Y(_1717_) );
INVX2 INVX2_107 ( .A(micro_hash_ucr_Wx_60_), .Y(_1718_) );
OAI21X1 OAI21X1_471 ( .A(_1718_), .B(_1438__bF_buf5), .C(_1493_), .Y(_1719_) );
XNOR2X1 XNOR2X1_96 ( .A(_1678__bF_buf4), .B(micro_hash_ucr_Wx_61_), .Y(_1720_) );
XNOR2X1 XNOR2X1_97 ( .A(_1719_), .B(_1720_), .Y(_1721_) );
NAND2X1 NAND2X1_276 ( .A(micro_hash_ucr_Wx_4_), .B(_1665__bF_buf1), .Y(_1722_) );
OAI21X1 OAI21X1_472 ( .A(_1445_), .B(_1443_), .C(_1722_), .Y(_1723_) );
INVX2 INVX2_108 ( .A(micro_hash_ucr_Wx_5_), .Y(_1724_) );
XNOR2X1 XNOR2X1_98 ( .A(_1678__bF_buf2), .B(_1724_), .Y(_1725_) );
XNOR2X1 XNOR2X1_99 ( .A(_1725_), .B(_1723_), .Y(_1726_) );
INVX1 INVX1_250 ( .A(H_21_), .Y(_1727_) );
NOR2X1 NOR2X1_428 ( .A(_4252_), .B(_1727_), .Y(_1728_) );
INVX1 INVX1_251 ( .A(micro_hash_ucr_c_5_), .Y(_1729_) );
OAI21X1 OAI21X1_473 ( .A(_1729_), .B(micro_hash_ucr_pipe6), .C(_438_), .Y(_1730_) );
OAI21X1 OAI21X1_474 ( .A(_1730_), .B(_1728_), .C(_4243_), .Y(_1731_) );
AOI21X1 AOI21X1_180 ( .A(micro_hash_ucr_pipe8), .B(_1726_), .C(_1731_), .Y(_1732_) );
INVX1 INVX1_252 ( .A(_1441_), .Y(_1733_) );
NOR2X1 NOR2X1_429 ( .A(_1733_), .B(_1439_), .Y(_1734_) );
AOI21X1 AOI21X1_181 ( .A(micro_hash_ucr_Wx_12_), .B(_1665__bF_buf1), .C(_1734_), .Y(_1735_) );
NOR2X1 NOR2X1_430 ( .A(micro_hash_ucr_Wx_13_), .B(_1678__bF_buf2), .Y(_1736_) );
INVX1 INVX1_253 ( .A(_1736_), .Y(_1737_) );
NAND2X1 NAND2X1_277 ( .A(micro_hash_ucr_Wx_13_), .B(_1678__bF_buf2), .Y(_1738_) );
NAND2X1 NAND2X1_278 ( .A(_1738_), .B(_1737_), .Y(_1739_) );
XNOR2X1 XNOR2X1_100 ( .A(_1739_), .B(_1735_), .Y(_1740_) );
OAI21X1 OAI21X1_475 ( .A(_1740_), .B(_4243_), .C(_4258_), .Y(_1741_) );
AOI21X1 AOI21X1_182 ( .A(micro_hash_ucr_Wx_20_), .B(_1665__bF_buf1), .C(_1454_), .Y(_1742_) );
INVX1 INVX1_254 ( .A(_1742_), .Y(_1743_) );
INVX2 INVX2_109 ( .A(micro_hash_ucr_Wx_21_), .Y(_1744_) );
OAI21X1 OAI21X1_476 ( .A(_1675_), .B(_1673__bF_buf1), .C(_1744_), .Y(_1745_) );
NAND2X1 NAND2X1_279 ( .A(micro_hash_ucr_Wx_21_), .B(_1678__bF_buf2), .Y(_1746_) );
NAND2X1 NAND2X1_280 ( .A(_1745_), .B(_1746_), .Y(_1747_) );
AOI21X1 AOI21X1_183 ( .A(_1747_), .B(_1743_), .C(_4258_), .Y(_1748_) );
OAI21X1 OAI21X1_477 ( .A(_1743_), .B(_1747_), .C(_1748_), .Y(_1749_) );
OAI21X1 OAI21X1_478 ( .A(_1741_), .B(_1732_), .C(_1749_), .Y(_1750_) );
NAND2X1 NAND2X1_281 ( .A(_4241__bF_buf2), .B(_1750_), .Y(_1751_) );
INVX1 INVX1_255 ( .A(_1459_), .Y(_1752_) );
NOR2X1 NOR2X1_431 ( .A(_1752_), .B(_1460_), .Y(_1753_) );
AOI21X1 AOI21X1_184 ( .A(micro_hash_ucr_Wx_28_), .B(_1665__bF_buf1), .C(_1753_), .Y(_1754_) );
INVX2 INVX2_110 ( .A(micro_hash_ucr_Wx_29_), .Y(_1755_) );
OAI21X1 OAI21X1_479 ( .A(_1675_), .B(_1673__bF_buf1), .C(_1755_), .Y(_1756_) );
INVX1 INVX1_256 ( .A(_1756_), .Y(_1757_) );
NOR2X1 NOR2X1_432 ( .A(_1755_), .B(_1679__bF_buf3), .Y(_1758_) );
NOR2X1 NOR2X1_433 ( .A(_1757_), .B(_1758_), .Y(_1759_) );
XNOR2X1 XNOR2X1_101 ( .A(_1754_), .B(_1759_), .Y(_1760_) );
OAI21X1 OAI21X1_480 ( .A(_4241__bF_buf2), .B(_1760_), .C(_1751_), .Y(_1761_) );
INVX2 INVX2_111 ( .A(micro_hash_ucr_Wx_36_), .Y(_1762_) );
OAI21X1 OAI21X1_481 ( .A(_1762_), .B(_1438__bF_buf5), .C(_1467_), .Y(_1763_) );
XNOR2X1 XNOR2X1_102 ( .A(_1678__bF_buf4), .B(micro_hash_ucr_Wx_37_), .Y(_1764_) );
XNOR2X1 XNOR2X1_103 ( .A(_1763_), .B(_1764_), .Y(_1765_) );
OAI21X1 OAI21X1_482 ( .A(_1765_), .B(_4239__bF_buf4), .C(_624__bF_buf0), .Y(_1766_) );
AOI21X1 AOI21X1_185 ( .A(_4239__bF_buf4), .B(_1761_), .C(_1766_), .Y(_1767_) );
AOI21X1 AOI21X1_186 ( .A(micro_hash_ucr_Wx_44_), .B(_1665__bF_buf1), .C(_1476_), .Y(_1768_) );
INVX2 INVX2_112 ( .A(micro_hash_ucr_Wx_45_), .Y(_1769_) );
OAI21X1 OAI21X1_483 ( .A(_1675_), .B(_1673__bF_buf1), .C(_1769_), .Y(_1770_) );
NAND2X1 NAND2X1_282 ( .A(micro_hash_ucr_Wx_45_), .B(_1678__bF_buf4), .Y(_1771_) );
NAND2X1 NAND2X1_283 ( .A(_1770_), .B(_1771_), .Y(_1772_) );
AND2X2 AND2X2_61 ( .A(_1768_), .B(_1772_), .Y(_1773_) );
OAI21X1 OAI21X1_484 ( .A(_1768_), .B(_1772_), .C(micro_hash_ucr_pipe18_bF_buf2), .Y(_1774_) );
OAI21X1 OAI21X1_485 ( .A(_1773_), .B(_1774_), .C(_4237__bF_buf4), .Y(_1775_) );
INVX2 INVX2_113 ( .A(micro_hash_ucr_Wx_52_), .Y(_1776_) );
OAI21X1 OAI21X1_486 ( .A(_1776_), .B(_1438__bF_buf3), .C(_1483_), .Y(_1777_) );
INVX2 INVX2_114 ( .A(micro_hash_ucr_Wx_53_), .Y(_1778_) );
OAI21X1 OAI21X1_487 ( .A(_1675_), .B(_1673__bF_buf1), .C(_1778_), .Y(_1779_) );
NOR2X1 NOR2X1_434 ( .A(_1778_), .B(_1679__bF_buf3), .Y(_1780_) );
INVX1 INVX1_257 ( .A(_1780_), .Y(_1781_) );
NAND2X1 NAND2X1_284 ( .A(_1779_), .B(_1781_), .Y(_1782_) );
AOI21X1 AOI21X1_187 ( .A(_1777_), .B(_1782_), .C(_4237__bF_buf4), .Y(_1783_) );
OAI21X1 OAI21X1_488 ( .A(_1777_), .B(_1782_), .C(_1783_), .Y(_1784_) );
OAI21X1 OAI21X1_489 ( .A(_1767_), .B(_1775_), .C(_1784_), .Y(_1785_) );
NAND2X1 NAND2X1_285 ( .A(_4262__bF_buf1), .B(_1785_), .Y(_1786_) );
OAI21X1 OAI21X1_490 ( .A(_4262__bF_buf1), .B(_1721_), .C(_1786_), .Y(_1787_) );
AOI21X1 AOI21X1_188 ( .A(micro_hash_ucr_Wx_68_), .B(_1665__bF_buf0), .C(_1500_), .Y(_1788_) );
INVX2 INVX2_115 ( .A(micro_hash_ucr_Wx_69_), .Y(_1789_) );
OAI21X1 OAI21X1_491 ( .A(_1675_), .B(_1673__bF_buf0), .C(_1789_), .Y(_1790_) );
NAND2X1 NAND2X1_286 ( .A(micro_hash_ucr_Wx_69_), .B(_1678__bF_buf4), .Y(_1791_) );
NAND2X1 NAND2X1_287 ( .A(_1790_), .B(_1791_), .Y(_1792_) );
XOR2X1 XOR2X1_29 ( .A(_1788_), .B(_1792_), .Y(_1793_) );
OAI21X1 OAI21X1_492 ( .A(_1793_), .B(_4233__bF_buf1), .C(_4230__bF_buf3), .Y(_1794_) );
AOI21X1 AOI21X1_189 ( .A(_4233__bF_buf1), .B(_1787_), .C(_1794_), .Y(_1795_) );
INVX2 INVX2_116 ( .A(micro_hash_ucr_Wx_76_), .Y(_1796_) );
NAND2X1 NAND2X1_288 ( .A(_1505_), .B(_1503_), .Y(_1797_) );
OAI21X1 OAI21X1_493 ( .A(_1796_), .B(_1438__bF_buf2), .C(_1797_), .Y(_1798_) );
INVX2 INVX2_117 ( .A(micro_hash_ucr_Wx_77_), .Y(_1799_) );
OAI21X1 OAI21X1_494 ( .A(_1675_), .B(_1673__bF_buf0), .C(_1799_), .Y(_1800_) );
NOR2X1 NOR2X1_435 ( .A(_1799_), .B(_1679__bF_buf3), .Y(_1801_) );
INVX1 INVX1_258 ( .A(_1801_), .Y(_1802_) );
NAND2X1 NAND2X1_289 ( .A(_1800_), .B(_1802_), .Y(_1803_) );
XOR2X1 XOR2X1_30 ( .A(_1803_), .B(_1798_), .Y(_1804_) );
OAI21X1 OAI21X1_495 ( .A(_1804_), .B(_4230__bF_buf3), .C(_220__bF_buf3), .Y(_1805_) );
INVX2 INVX2_118 ( .A(micro_hash_ucr_Wx_84_), .Y(_1806_) );
OAI21X1 OAI21X1_496 ( .A(_1806_), .B(_1438__bF_buf5), .C(_1515_), .Y(_1807_) );
XNOR2X1 XNOR2X1_104 ( .A(_1678__bF_buf3), .B(micro_hash_ucr_Wx_85_), .Y(_1808_) );
AOI21X1 AOI21X1_190 ( .A(_1808_), .B(_1807_), .C(_220__bF_buf3), .Y(_1809_) );
OAI21X1 OAI21X1_497 ( .A(_1807_), .B(_1808_), .C(_1809_), .Y(_1810_) );
OAI21X1 OAI21X1_498 ( .A(_1795_), .B(_1805_), .C(_1810_), .Y(_1811_) );
NAND2X1 NAND2X1_290 ( .A(_4228__bF_buf3), .B(_1811_), .Y(_1812_) );
OAI21X1 OAI21X1_499 ( .A(_4228__bF_buf3), .B(_1717_), .C(_1812_), .Y(_1813_) );
AOI21X1 AOI21X1_191 ( .A(micro_hash_ucr_Wx_100_), .B(_1665__bF_buf0), .C(_1528_), .Y(_1814_) );
NOR2X1 NOR2X1_436 ( .A(micro_hash_ucr_Wx_101_), .B(_1678__bF_buf3), .Y(_1815_) );
INVX2 INVX2_119 ( .A(micro_hash_ucr_Wx_101_), .Y(_1816_) );
NOR2X1 NOR2X1_437 ( .A(_1816_), .B(_1679__bF_buf0), .Y(_1817_) );
NOR2X1 NOR2X1_438 ( .A(_1815_), .B(_1817_), .Y(_1818_) );
AND2X2 AND2X2_62 ( .A(_1818_), .B(_1814_), .Y(_1819_) );
OAI21X1 OAI21X1_500 ( .A(_1818_), .B(_1814_), .C(micro_hash_ucr_pipe32_bF_buf4), .Y(_1820_) );
OAI21X1 OAI21X1_501 ( .A(_1819_), .B(_1820_), .C(_4225__bF_buf1), .Y(_1821_) );
AOI21X1 AOI21X1_192 ( .A(_4226__bF_buf2), .B(_1813_), .C(_1821_), .Y(_1822_) );
AOI21X1 AOI21X1_193 ( .A(micro_hash_ucr_Wx_108_), .B(_1665__bF_buf1), .C(_1536_), .Y(_1823_) );
XNOR2X1 XNOR2X1_105 ( .A(_1678__bF_buf3), .B(micro_hash_ucr_Wx_109_), .Y(_1824_) );
AND2X2 AND2X2_63 ( .A(_1824_), .B(_1823_), .Y(_1825_) );
OAI21X1 OAI21X1_502 ( .A(_1824_), .B(_1823_), .C(micro_hash_ucr_pipe34_bF_buf0), .Y(_1826_) );
OAI21X1 OAI21X1_503 ( .A(_1825_), .B(_1826_), .C(_4224__bF_buf1), .Y(_1827_) );
INVX2 INVX2_120 ( .A(micro_hash_ucr_Wx_116_), .Y(_1828_) );
OAI21X1 OAI21X1_504 ( .A(_1828_), .B(_1438__bF_buf0), .C(_1544_), .Y(_1829_) );
XNOR2X1 XNOR2X1_106 ( .A(_1678__bF_buf4), .B(micro_hash_ucr_Wx_117_), .Y(_1830_) );
AOI21X1 AOI21X1_194 ( .A(_1830_), .B(_1829_), .C(_4224__bF_buf1), .Y(_1831_) );
OAI21X1 OAI21X1_505 ( .A(_1829_), .B(_1830_), .C(_1831_), .Y(_1832_) );
OAI21X1 OAI21X1_506 ( .A(_1822_), .B(_1827_), .C(_1832_), .Y(_1833_) );
NAND2X1 NAND2X1_291 ( .A(_701__bF_buf4), .B(_1833_), .Y(_1834_) );
OAI21X1 OAI21X1_507 ( .A(_701__bF_buf4), .B(_1710_), .C(_1834_), .Y(_1835_) );
AOI21X1 AOI21X1_195 ( .A(micro_hash_ucr_Wx_132_), .B(_1665__bF_buf0), .C(_1558_), .Y(_1836_) );
NOR2X1 NOR2X1_439 ( .A(micro_hash_ucr_Wx_133_), .B(_1678__bF_buf0), .Y(_1837_) );
INVX2 INVX2_121 ( .A(micro_hash_ucr_Wx_133_), .Y(_1838_) );
NOR2X1 NOR2X1_440 ( .A(_1838_), .B(_1679__bF_buf1), .Y(_1839_) );
NOR2X1 NOR2X1_441 ( .A(_1837_), .B(_1839_), .Y(_1840_) );
AND2X2 AND2X2_64 ( .A(_1840_), .B(_1836_), .Y(_1841_) );
OAI21X1 OAI21X1_508 ( .A(_1840_), .B(_1836_), .C(micro_hash_ucr_pipe40_bF_buf3), .Y(_1842_) );
OAI21X1 OAI21X1_509 ( .A(_1841_), .B(_1842_), .C(_4220__bF_buf4), .Y(_1843_) );
AOI21X1 AOI21X1_196 ( .A(_296__bF_buf4), .B(_1835_), .C(_1843_), .Y(_1844_) );
AOI21X1 AOI21X1_197 ( .A(micro_hash_ucr_Wx_140_), .B(_1665__bF_buf0), .C(_1567_), .Y(_1845_) );
XNOR2X1 XNOR2X1_107 ( .A(_1678__bF_buf0), .B(micro_hash_ucr_Wx_141_), .Y(_1846_) );
AND2X2 AND2X2_65 ( .A(_1846_), .B(_1845_), .Y(_1847_) );
OAI21X1 OAI21X1_510 ( .A(_1846_), .B(_1845_), .C(micro_hash_ucr_pipe42_bF_buf2), .Y(_1848_) );
OAI21X1 OAI21X1_511 ( .A(_1847_), .B(_1848_), .C(_4219__bF_buf1), .Y(_1849_) );
INVX1 INVX1_259 ( .A(micro_hash_ucr_Wx_148_), .Y(_1850_) );
OAI21X1 OAI21X1_512 ( .A(_1850_), .B(_1438__bF_buf0), .C(_1575_), .Y(_1851_) );
XNOR2X1 XNOR2X1_108 ( .A(_1678__bF_buf1), .B(micro_hash_ucr_Wx_149_), .Y(_1852_) );
AOI21X1 AOI21X1_198 ( .A(_1852_), .B(_1851_), .C(_4219__bF_buf1), .Y(_1853_) );
OAI21X1 OAI21X1_513 ( .A(_1851_), .B(_1852_), .C(_1853_), .Y(_1854_) );
OAI21X1 OAI21X1_514 ( .A(_1844_), .B(_1849_), .C(_1854_), .Y(_1855_) );
NAND2X1 NAND2X1_292 ( .A(_4218__bF_buf3), .B(_1855_), .Y(_1856_) );
OAI21X1 OAI21X1_515 ( .A(_4218__bF_buf3), .B(_1702_), .C(_1856_), .Y(_1857_) );
INVX1 INVX1_260 ( .A(micro_hash_ucr_Wx_164_), .Y(_1858_) );
OAI21X1 OAI21X1_516 ( .A(_1858_), .B(_1438__bF_buf0), .C(_1589_), .Y(_1859_) );
XNOR2X1 XNOR2X1_109 ( .A(_1678__bF_buf1), .B(micro_hash_ucr_Wx_165_), .Y(_1860_) );
XNOR2X1 XNOR2X1_110 ( .A(_1859_), .B(_1860_), .Y(_1861_) );
OAI21X1 OAI21X1_517 ( .A(_1861_), .B(_4217__bF_buf2), .C(_4215__bF_buf4), .Y(_1862_) );
AOI21X1 AOI21X1_199 ( .A(_4217__bF_buf2), .B(_1857_), .C(_1862_), .Y(_1863_) );
AOI21X1 AOI21X1_200 ( .A(micro_hash_ucr_Wx_172_), .B(_1665__bF_buf3), .C(_1596_), .Y(_1864_) );
INVX1 INVX1_261 ( .A(micro_hash_ucr_Wx_173_), .Y(_1865_) );
OAI21X1 OAI21X1_518 ( .A(_1675_), .B(_1673__bF_buf2), .C(_1865_), .Y(_1866_) );
NAND2X1 NAND2X1_293 ( .A(micro_hash_ucr_Wx_173_), .B(_1678__bF_buf0), .Y(_1867_) );
NAND2X1 NAND2X1_294 ( .A(_1866_), .B(_1867_), .Y(_1868_) );
AND2X2 AND2X2_66 ( .A(_1868_), .B(_1864_), .Y(_1869_) );
OAI21X1 OAI21X1_519 ( .A(_1868_), .B(_1864_), .C(micro_hash_ucr_pipe50_bF_buf2), .Y(_1870_) );
OAI21X1 OAI21X1_520 ( .A(_1869_), .B(_1870_), .C(_4214__bF_buf3), .Y(_1871_) );
AOI21X1 AOI21X1_201 ( .A(micro_hash_ucr_Wx_180_), .B(_1665__bF_buf3), .C(_1602_), .Y(_1872_) );
INVX2 INVX2_122 ( .A(_1872_), .Y(_1873_) );
INVX1 INVX1_262 ( .A(micro_hash_ucr_Wx_181_), .Y(_1874_) );
OAI21X1 OAI21X1_521 ( .A(_1675_), .B(_1673__bF_buf2), .C(_1874_), .Y(_1875_) );
NOR2X1 NOR2X1_442 ( .A(_1874_), .B(_1679__bF_buf1), .Y(_1876_) );
INVX1 INVX1_263 ( .A(_1876_), .Y(_1877_) );
NAND2X1 NAND2X1_295 ( .A(_1875_), .B(_1877_), .Y(_1878_) );
AOI21X1 AOI21X1_202 ( .A(_1873_), .B(_1878_), .C(_4214__bF_buf3), .Y(_1879_) );
OAI21X1 OAI21X1_522 ( .A(_1873_), .B(_1878_), .C(_1879_), .Y(_1880_) );
OAI21X1 OAI21X1_523 ( .A(_1863_), .B(_1871_), .C(_1880_), .Y(_1881_) );
NAND2X1 NAND2X1_296 ( .A(_742__bF_buf3), .B(_1881_), .Y(_1882_) );
OAI21X1 OAI21X1_524 ( .A(_742__bF_buf3), .B(_1696_), .C(_1882_), .Y(_1883_) );
AOI21X1 AOI21X1_203 ( .A(micro_hash_ucr_Wx_196_), .B(_1665__bF_buf2), .C(_1616_), .Y(_1884_) );
INVX2 INVX2_123 ( .A(micro_hash_ucr_Wx_197_), .Y(_1885_) );
XNOR2X1 XNOR2X1_111 ( .A(_1678__bF_buf1), .B(_1885_), .Y(_1886_) );
AND2X2 AND2X2_67 ( .A(_1884_), .B(_1886_), .Y(_1887_) );
OAI21X1 OAI21X1_525 ( .A(_1884_), .B(_1886_), .C(micro_hash_ucr_pipe56_bF_buf3), .Y(_1888_) );
OAI21X1 OAI21X1_526 ( .A(_1887_), .B(_1888_), .C(_4211__bF_buf3), .Y(_1889_) );
AOI21X1 AOI21X1_204 ( .A(_832__bF_buf3), .B(_1883_), .C(_1889_), .Y(_1890_) );
AOI21X1 AOI21X1_205 ( .A(micro_hash_ucr_Wx_204_), .B(_1665__bF_buf2), .C(_1622_), .Y(_1891_) );
NOR2X1 NOR2X1_443 ( .A(micro_hash_ucr_Wx_205_), .B(_1678__bF_buf5), .Y(_1892_) );
INVX1 INVX1_264 ( .A(_1892_), .Y(_1893_) );
NAND2X1 NAND2X1_297 ( .A(micro_hash_ucr_Wx_205_), .B(_1678__bF_buf5), .Y(_1894_) );
NAND2X1 NAND2X1_298 ( .A(_1894_), .B(_1893_), .Y(_1895_) );
AND2X2 AND2X2_68 ( .A(_1895_), .B(_1891_), .Y(_1896_) );
OAI21X1 OAI21X1_527 ( .A(_1895_), .B(_1891_), .C(micro_hash_ucr_pipe58_bF_buf1), .Y(_1897_) );
OAI21X1 OAI21X1_528 ( .A(_1896_), .B(_1897_), .C(_4210__bF_buf4), .Y(_1898_) );
AOI21X1 AOI21X1_206 ( .A(micro_hash_ucr_Wx_212_), .B(_1665__bF_buf3), .C(_1630_), .Y(_1899_) );
INVX1 INVX1_265 ( .A(_1899_), .Y(_1900_) );
NOR2X1 NOR2X1_444 ( .A(micro_hash_ucr_Wx_213_), .B(_1678__bF_buf5), .Y(_1901_) );
INVX1 INVX1_266 ( .A(_1901_), .Y(_1902_) );
NAND2X1 NAND2X1_299 ( .A(micro_hash_ucr_Wx_213_), .B(_1678__bF_buf5), .Y(_1903_) );
NAND2X1 NAND2X1_300 ( .A(_1903_), .B(_1902_), .Y(_1904_) );
AOI21X1 AOI21X1_207 ( .A(_1904_), .B(_1900_), .C(_4210__bF_buf4), .Y(_1905_) );
OAI21X1 OAI21X1_529 ( .A(_1900_), .B(_1904_), .C(_1905_), .Y(_1906_) );
OAI21X1 OAI21X1_530 ( .A(_1890_), .B(_1898_), .C(_1906_), .Y(_1907_) );
NAND2X1 NAND2X1_301 ( .A(_4207__bF_buf1), .B(_1907_), .Y(_1908_) );
OAI21X1 OAI21X1_531 ( .A(_4207__bF_buf1), .B(_1689_), .C(_1908_), .Y(_1909_) );
INVX1 INVX1_267 ( .A(_1641_), .Y(_1910_) );
NOR2X1 NOR2X1_445 ( .A(_1642_), .B(_1910_), .Y(_1911_) );
AOI21X1 AOI21X1_208 ( .A(micro_hash_ucr_Wx_228_), .B(_1665__bF_buf2), .C(_1911_), .Y(_1912_) );
INVX1 INVX1_268 ( .A(micro_hash_ucr_Wx_229_), .Y(_1913_) );
OAI21X1 OAI21X1_532 ( .A(_1675_), .B(_1673__bF_buf3), .C(_1913_), .Y(_1914_) );
INVX1 INVX1_269 ( .A(_1914_), .Y(_1915_) );
NOR2X1 NOR2X1_446 ( .A(_1913_), .B(_1679__bF_buf0), .Y(_1916_) );
NOR2X1 NOR2X1_447 ( .A(_1915_), .B(_1916_), .Y(_1917_) );
AND2X2 AND2X2_69 ( .A(_1917_), .B(_1912_), .Y(_1918_) );
OAI21X1 OAI21X1_533 ( .A(_1917_), .B(_1912_), .C(micro_hash_ucr_pipe64_bF_buf3), .Y(_1919_) );
OAI21X1 OAI21X1_534 ( .A(_1918_), .B(_1919_), .C(_1078__bF_buf3), .Y(_1920_) );
AOI21X1 AOI21X1_209 ( .A(_278__bF_buf2), .B(_1909_), .C(_1920_), .Y(_1921_) );
AOI21X1 AOI21X1_210 ( .A(micro_hash_ucr_Wx_236_), .B(_1665__bF_buf2), .C(_1648_), .Y(_1922_) );
XNOR2X1 XNOR2X1_112 ( .A(_1678__bF_buf0), .B(micro_hash_ucr_Wx_237_), .Y(_1923_) );
AND2X2 AND2X2_70 ( .A(_1923_), .B(_1922_), .Y(_1924_) );
OAI21X1 OAI21X1_535 ( .A(_1923_), .B(_1922_), .C(micro_hash_ucr_pipe66_bF_buf3), .Y(_1925_) );
OAI21X1 OAI21X1_536 ( .A(_1924_), .B(_1925_), .C(_4199__bF_buf5), .Y(_1926_) );
OAI21X1 OAI21X1_537 ( .A(_1921_), .B(_1926_), .C(_1683_), .Y(_1927_) );
NAND2X1 NAND2X1_302 ( .A(micro_hash_ucr_Wx_252_), .B(_1665__bF_buf2), .Y(_1928_) );
OAI21X1 OAI21X1_538 ( .A(_1661_), .B(_1662_), .C(_1928_), .Y(_1929_) );
INVX1 INVX1_270 ( .A(micro_hash_ucr_Wx_253_), .Y(_1930_) );
OAI21X1 OAI21X1_539 ( .A(_1675_), .B(_1673__bF_buf3), .C(_1930_), .Y(_1931_) );
NOR2X1 NOR2X1_448 ( .A(_1930_), .B(_1679__bF_buf0), .Y(_1932_) );
INVX1 INVX1_271 ( .A(_1932_), .Y(_1933_) );
NAND2X1 NAND2X1_303 ( .A(_1931_), .B(_1933_), .Y(_1934_) );
XNOR2X1 XNOR2X1_113 ( .A(_1934_), .B(_1929_), .Y(_1935_) );
OAI21X1 OAI21X1_540 ( .A(_1935_), .B(_287_), .C(_131__bF_buf10), .Y(_1936_) );
AOI21X1 AOI21X1_211 ( .A(_287_), .B(_1927_), .C(_1936_), .Y(_128__5_) );
OAI21X1 OAI21X1_541 ( .A(_299_), .B(_392_), .C(_1672_), .Y(_1937_) );
XOR2X1 XOR2X1_31 ( .A(micro_hash_ucr_k_6_), .B(micro_hash_ucr_x_6_), .Y(_1938_) );
NOR2X1 NOR2X1_449 ( .A(_1938_), .B(_1937_), .Y(_1939_) );
OAI21X1 OAI21X1_542 ( .A(_1673__bF_buf3), .B(_1669_), .C(_1938_), .Y(_1940_) );
INVX1 INVX1_272 ( .A(_1940_), .Y(_1941_) );
NOR2X1 NOR2X1_450 ( .A(_1939_), .B(_1941_), .Y(_1942_) );
XNOR2X1 XNOR2X1_114 ( .A(_1942__bF_buf4), .B(micro_hash_ucr_Wx_14_), .Y(_1943_) );
OAI21X1 OAI21X1_543 ( .A(_1735_), .B(_1736_), .C(_1738_), .Y(_1944_) );
XNOR2X1 XNOR2X1_115 ( .A(_1944_), .B(_1943_), .Y(_1945_) );
INVX2 INVX2_124 ( .A(micro_hash_ucr_Wx_6_), .Y(_1946_) );
XNOR2X1 XNOR2X1_116 ( .A(_1942__bF_buf4), .B(_1946_), .Y(_1947_) );
OAI21X1 OAI21X1_544 ( .A(micro_hash_ucr_Wx_5_), .B(_1678__bF_buf2), .C(_1723_), .Y(_1948_) );
OAI21X1 OAI21X1_545 ( .A(_1724_), .B(_1679__bF_buf3), .C(_1948_), .Y(_1949_) );
AOI21X1 AOI21X1_212 ( .A(_1947_), .B(_1949_), .C(_438_), .Y(_1950_) );
OAI21X1 OAI21X1_546 ( .A(_1947_), .B(_1949_), .C(_1950_), .Y(_1951_) );
INVX1 INVX1_273 ( .A(H_22_), .Y(_1952_) );
NAND2X1 NAND2X1_304 ( .A(micro_hash_ucr_pipe6), .B(_1952_), .Y(_1953_) );
OAI21X1 OAI21X1_547 ( .A(micro_hash_ucr_pipe6), .B(micro_hash_ucr_c_6_), .C(_1953_), .Y(_1954_) );
OAI21X1 OAI21X1_548 ( .A(micro_hash_ucr_pipe8), .B(_1954_), .C(_1951_), .Y(_1955_) );
MUX2X1 MUX2X1_44 ( .A(_1955_), .B(_1945_), .S(_4243_), .Y(_1956_) );
INVX4 INVX4_28 ( .A(micro_hash_ucr_Wx_22_), .Y(_1957_) );
XNOR2X1 XNOR2X1_117 ( .A(_1942__bF_buf4), .B(_1957_), .Y(_1958_) );
INVX1 INVX1_274 ( .A(_1745_), .Y(_1959_) );
OAI21X1 OAI21X1_549 ( .A(_1742_), .B(_1959_), .C(_1746_), .Y(_1960_) );
XNOR2X1 XNOR2X1_118 ( .A(_1960_), .B(_1958_), .Y(_1961_) );
MUX2X1 MUX2X1_45 ( .A(_1956_), .B(_1961_), .S(_4258_), .Y(_1962_) );
INVX4 INVX4_29 ( .A(micro_hash_ucr_Wx_30_), .Y(_1963_) );
XNOR2X1 XNOR2X1_119 ( .A(_1942__bF_buf4), .B(_1963_), .Y(_1964_) );
INVX1 INVX1_275 ( .A(_1758_), .Y(_1965_) );
OAI21X1 OAI21X1_550 ( .A(_1754_), .B(_1757_), .C(_1965_), .Y(_1966_) );
XOR2X1 XOR2X1_32 ( .A(_1966_), .B(_1964_), .Y(_1967_) );
MUX2X1 MUX2X1_46 ( .A(_1962_), .B(_1967_), .S(_4241__bF_buf2), .Y(_1968_) );
NOR2X1 NOR2X1_451 ( .A(micro_hash_ucr_pipe16), .B(_1968_), .Y(_1969_) );
INVX4 INVX4_30 ( .A(micro_hash_ucr_Wx_38_), .Y(_1970_) );
XNOR2X1 XNOR2X1_120 ( .A(_1942__bF_buf2), .B(_1970_), .Y(_1971_) );
INVX2 INVX2_125 ( .A(micro_hash_ucr_Wx_37_), .Y(_1972_) );
OAI21X1 OAI21X1_551 ( .A(micro_hash_ucr_Wx_37_), .B(_1678__bF_buf4), .C(_1763_), .Y(_1973_) );
OAI21X1 OAI21X1_552 ( .A(_1972_), .B(_1679__bF_buf3), .C(_1973_), .Y(_1974_) );
XNOR2X1 XNOR2X1_121 ( .A(_1974_), .B(_1971_), .Y(_1975_) );
OAI21X1 OAI21X1_553 ( .A(_1975_), .B(_4239__bF_buf4), .C(_624__bF_buf3), .Y(_1976_) );
INVX2 INVX2_126 ( .A(micro_hash_ucr_Wx_46_), .Y(_1977_) );
XNOR2X1 XNOR2X1_122 ( .A(_1942__bF_buf2), .B(_1977_), .Y(_1978_) );
INVX1 INVX1_276 ( .A(_1770_), .Y(_1979_) );
OAI21X1 OAI21X1_554 ( .A(_1768_), .B(_1979_), .C(_1771_), .Y(_1980_) );
NOR2X1 NOR2X1_452 ( .A(_1978_), .B(_1980_), .Y(_1981_) );
AND2X2 AND2X2_71 ( .A(_1980_), .B(_1978_), .Y(_1982_) );
OAI21X1 OAI21X1_555 ( .A(_1982_), .B(_1981_), .C(micro_hash_ucr_pipe18_bF_buf2), .Y(_1983_) );
OAI21X1 OAI21X1_556 ( .A(_1969_), .B(_1976_), .C(_1983_), .Y(_1984_) );
INVX4 INVX4_31 ( .A(micro_hash_ucr_Wx_54_), .Y(_1985_) );
XNOR2X1 XNOR2X1_123 ( .A(_1942__bF_buf2), .B(_1985_), .Y(_1986_) );
INVX1 INVX1_277 ( .A(_1986_), .Y(_1987_) );
AOI21X1 AOI21X1_213 ( .A(_1779_), .B(_1777_), .C(_1780_), .Y(_1988_) );
OR2X2 OR2X2_13 ( .A(_1988_), .B(_1987_), .Y(_1989_) );
NAND2X1 NAND2X1_305 ( .A(_1987_), .B(_1988_), .Y(_1990_) );
AOI21X1 AOI21X1_214 ( .A(_1990_), .B(_1989_), .C(_4237__bF_buf4), .Y(_1991_) );
AOI21X1 AOI21X1_215 ( .A(_4237__bF_buf4), .B(_1984_), .C(_1991_), .Y(_1992_) );
NOR2X1 NOR2X1_453 ( .A(micro_hash_ucr_pipe22_bF_buf1), .B(_1992_), .Y(_1993_) );
INVX4 INVX4_32 ( .A(micro_hash_ucr_Wx_62_), .Y(_1994_) );
XNOR2X1 XNOR2X1_124 ( .A(_1942__bF_buf4), .B(_1994_), .Y(_1995_) );
INVX2 INVX2_127 ( .A(micro_hash_ucr_Wx_61_), .Y(_1996_) );
OAI21X1 OAI21X1_557 ( .A(micro_hash_ucr_Wx_61_), .B(_1678__bF_buf2), .C(_1719_), .Y(_1997_) );
OAI21X1 OAI21X1_558 ( .A(_1996_), .B(_1679__bF_buf3), .C(_1997_), .Y(_1998_) );
OR2X2 OR2X2_14 ( .A(_1998_), .B(_1995_), .Y(_1999_) );
NAND2X1 NAND2X1_306 ( .A(_1995_), .B(_1998_), .Y(_2000_) );
AOI21X1 AOI21X1_216 ( .A(_2000_), .B(_1999_), .C(_4262__bF_buf1), .Y(_2001_) );
OAI21X1 OAI21X1_559 ( .A(_1993_), .B(_2001_), .C(_4233__bF_buf1), .Y(_2002_) );
INVX4 INVX4_33 ( .A(micro_hash_ucr_Wx_70_), .Y(_2003_) );
XNOR2X1 XNOR2X1_125 ( .A(_1942__bF_buf5), .B(_2003_), .Y(_2004_) );
INVX1 INVX1_278 ( .A(_1790_), .Y(_2005_) );
OAI21X1 OAI21X1_560 ( .A(_1788_), .B(_2005_), .C(_1791_), .Y(_2006_) );
NOR2X1 NOR2X1_454 ( .A(_2004_), .B(_2006_), .Y(_2007_) );
NAND2X1 NAND2X1_307 ( .A(_2004_), .B(_2006_), .Y(_2008_) );
INVX1 INVX1_279 ( .A(_2008_), .Y(_2009_) );
OAI21X1 OAI21X1_561 ( .A(_2009_), .B(_2007_), .C(micro_hash_ucr_pipe24_bF_buf0), .Y(_2010_) );
NAND3X1 NAND3X1_96 ( .A(_4230__bF_buf3), .B(_2010_), .C(_2002_), .Y(_2011_) );
XNOR2X1 XNOR2X1_126 ( .A(_1942__bF_buf2), .B(micro_hash_ucr_Wx_78_), .Y(_2012_) );
AOI21X1 AOI21X1_217 ( .A(_1800_), .B(_1798_), .C(_1801_), .Y(_2013_) );
OR2X2 OR2X2_15 ( .A(_2012_), .B(_2013_), .Y(_2014_) );
NAND2X1 NAND2X1_308 ( .A(_2013_), .B(_2012_), .Y(_2015_) );
NAND2X1 NAND2X1_309 ( .A(_2015_), .B(_2014_), .Y(_2016_) );
OAI21X1 OAI21X1_562 ( .A(_4230__bF_buf3), .B(_2016_), .C(_2011_), .Y(_2017_) );
NOR2X1 NOR2X1_455 ( .A(micro_hash_ucr_pipe28_bF_buf3), .B(_2017_), .Y(_2018_) );
INVX4 INVX4_34 ( .A(micro_hash_ucr_Wx_86_), .Y(_2019_) );
XNOR2X1 XNOR2X1_127 ( .A(_1942__bF_buf5), .B(_2019_), .Y(_2020_) );
INVX2 INVX2_128 ( .A(micro_hash_ucr_Wx_85_), .Y(_2021_) );
OAI21X1 OAI21X1_563 ( .A(micro_hash_ucr_Wx_85_), .B(_1678__bF_buf3), .C(_1807_), .Y(_2022_) );
OAI21X1 OAI21X1_564 ( .A(_2021_), .B(_1679__bF_buf2), .C(_2022_), .Y(_2023_) );
OR2X2 OR2X2_16 ( .A(_2023_), .B(_2020_), .Y(_2024_) );
NAND2X1 NAND2X1_310 ( .A(_2020_), .B(_2023_), .Y(_2025_) );
AOI21X1 AOI21X1_218 ( .A(_2025_), .B(_2024_), .C(_220__bF_buf3), .Y(_2026_) );
OAI21X1 OAI21X1_565 ( .A(_2018_), .B(_2026_), .C(_4228__bF_buf3), .Y(_2027_) );
XNOR2X1 XNOR2X1_128 ( .A(_1942__bF_buf2), .B(micro_hash_ucr_Wx_94_), .Y(_2028_) );
INVX1 INVX1_280 ( .A(_1715_), .Y(_2029_) );
OAI21X1 OAI21X1_566 ( .A(_1711_), .B(_1714_), .C(_2029_), .Y(_2030_) );
INVX1 INVX1_281 ( .A(_2030_), .Y(_2031_) );
NOR2X1 NOR2X1_456 ( .A(_2028_), .B(_2031_), .Y(_2032_) );
AND2X2 AND2X2_72 ( .A(_2031_), .B(_2028_), .Y(_2033_) );
OAI21X1 OAI21X1_567 ( .A(_2033_), .B(_2032_), .C(micro_hash_ucr_pipe30_bF_buf2), .Y(_2034_) );
NAND2X1 NAND2X1_311 ( .A(_2034_), .B(_2027_), .Y(_2035_) );
INVX4 INVX4_35 ( .A(micro_hash_ucr_Wx_102_), .Y(_2036_) );
XNOR2X1 XNOR2X1_129 ( .A(_1942__bF_buf5), .B(_2036_), .Y(_2037_) );
INVX1 INVX1_282 ( .A(_1817_), .Y(_2038_) );
OAI21X1 OAI21X1_568 ( .A(_1814_), .B(_1815_), .C(_2038_), .Y(_2039_) );
OR2X2 OR2X2_17 ( .A(_2039_), .B(_2037_), .Y(_2040_) );
NAND2X1 NAND2X1_312 ( .A(_2037_), .B(_2039_), .Y(_2041_) );
NAND3X1 NAND3X1_97 ( .A(micro_hash_ucr_pipe32_bF_buf4), .B(_2041_), .C(_2040_), .Y(_2042_) );
OAI21X1 OAI21X1_569 ( .A(_2035_), .B(micro_hash_ucr_pipe32_bF_buf4), .C(_2042_), .Y(_2043_) );
XNOR2X1 XNOR2X1_130 ( .A(_1942__bF_buf5), .B(micro_hash_ucr_Wx_110_), .Y(_2044_) );
INVX2 INVX2_129 ( .A(micro_hash_ucr_Wx_109_), .Y(_2045_) );
OAI21X1 OAI21X1_570 ( .A(_2045_), .B(_1679__bF_buf2), .C(_1823_), .Y(_2046_) );
OAI21X1 OAI21X1_571 ( .A(micro_hash_ucr_Wx_109_), .B(_1678__bF_buf3), .C(_2046_), .Y(_2047_) );
NOR2X1 NOR2X1_457 ( .A(_2044_), .B(_2047_), .Y(_2048_) );
AND2X2 AND2X2_73 ( .A(_2047_), .B(_2044_), .Y(_2049_) );
OAI21X1 OAI21X1_572 ( .A(_2049_), .B(_2048_), .C(micro_hash_ucr_pipe34_bF_buf0), .Y(_2050_) );
OAI21X1 OAI21X1_573 ( .A(_2043_), .B(micro_hash_ucr_pipe34_bF_buf0), .C(_2050_), .Y(_2051_) );
INVX2 INVX2_130 ( .A(micro_hash_ucr_Wx_118_), .Y(_2052_) );
XNOR2X1 XNOR2X1_131 ( .A(_1942__bF_buf2), .B(_2052_), .Y(_2053_) );
INVX2 INVX2_131 ( .A(micro_hash_ucr_Wx_117_), .Y(_2054_) );
OAI21X1 OAI21X1_574 ( .A(micro_hash_ucr_Wx_117_), .B(_1678__bF_buf4), .C(_1829_), .Y(_2055_) );
OAI21X1 OAI21X1_575 ( .A(_2054_), .B(_1679__bF_buf2), .C(_2055_), .Y(_2056_) );
OR2X2 OR2X2_18 ( .A(_2056_), .B(_2053_), .Y(_2057_) );
NAND2X1 NAND2X1_313 ( .A(_2053_), .B(_2056_), .Y(_2058_) );
AND2X2 AND2X2_74 ( .A(_2057_), .B(_2058_), .Y(_2059_) );
OAI21X1 OAI21X1_576 ( .A(_2059_), .B(_4224__bF_buf1), .C(_701__bF_buf4), .Y(_2060_) );
AOI21X1 AOI21X1_219 ( .A(_4224__bF_buf1), .B(_2051_), .C(_2060_), .Y(_2061_) );
INVX2 INVX2_132 ( .A(micro_hash_ucr_Wx_126_), .Y(_2062_) );
XNOR2X1 XNOR2X1_132 ( .A(_1942__bF_buf5), .B(_2062_), .Y(_2063_) );
INVX1 INVX1_283 ( .A(_2063_), .Y(_2064_) );
AOI21X1 AOI21X1_220 ( .A(_1706_), .B(_1704_), .C(_1707_), .Y(_2065_) );
OR2X2 OR2X2_19 ( .A(_2065_), .B(_2064_), .Y(_2066_) );
AOI21X1 AOI21X1_221 ( .A(_2064_), .B(_2065_), .C(_701__bF_buf4), .Y(_2067_) );
AOI21X1 AOI21X1_222 ( .A(_2066_), .B(_2067_), .C(_2061_), .Y(_2068_) );
INVX4 INVX4_36 ( .A(micro_hash_ucr_Wx_134_), .Y(_2069_) );
XNOR2X1 XNOR2X1_133 ( .A(_1942__bF_buf0), .B(_2069_), .Y(_2070_) );
INVX1 INVX1_284 ( .A(_1839_), .Y(_2071_) );
OAI21X1 OAI21X1_577 ( .A(_1836_), .B(_1837_), .C(_2071_), .Y(_2072_) );
OR2X2 OR2X2_20 ( .A(_2072_), .B(_2070_), .Y(_2073_) );
NAND2X1 NAND2X1_314 ( .A(_2070_), .B(_2072_), .Y(_2074_) );
NAND3X1 NAND3X1_98 ( .A(micro_hash_ucr_pipe40_bF_buf3), .B(_2074_), .C(_2073_), .Y(_2075_) );
OAI21X1 OAI21X1_578 ( .A(_2068_), .B(micro_hash_ucr_pipe40_bF_buf3), .C(_2075_), .Y(_2076_) );
XNOR2X1 XNOR2X1_134 ( .A(_1942__bF_buf0), .B(micro_hash_ucr_Wx_142_), .Y(_2077_) );
INVX2 INVX2_133 ( .A(micro_hash_ucr_Wx_141_), .Y(_2078_) );
OAI21X1 OAI21X1_579 ( .A(_2078_), .B(_1679__bF_buf2), .C(_1845_), .Y(_2079_) );
OAI21X1 OAI21X1_580 ( .A(micro_hash_ucr_Wx_141_), .B(_1678__bF_buf0), .C(_2079_), .Y(_2080_) );
NOR2X1 NOR2X1_458 ( .A(_2077_), .B(_2080_), .Y(_2081_) );
AND2X2 AND2X2_75 ( .A(_2080_), .B(_2077_), .Y(_2082_) );
OAI21X1 OAI21X1_581 ( .A(_2082_), .B(_2081_), .C(micro_hash_ucr_pipe42_bF_buf2), .Y(_2083_) );
OAI21X1 OAI21X1_582 ( .A(_2076_), .B(micro_hash_ucr_pipe42_bF_buf2), .C(_2083_), .Y(_2084_) );
INVX4 INVX4_37 ( .A(micro_hash_ucr_Wx_150_), .Y(_2085_) );
XNOR2X1 XNOR2X1_135 ( .A(_1942__bF_buf1), .B(_2085_), .Y(_2086_) );
INVX1 INVX1_285 ( .A(micro_hash_ucr_Wx_149_), .Y(_2087_) );
OAI21X1 OAI21X1_583 ( .A(micro_hash_ucr_Wx_149_), .B(_1678__bF_buf1), .C(_1851_), .Y(_2088_) );
OAI21X1 OAI21X1_584 ( .A(_2087_), .B(_1679__bF_buf1), .C(_2088_), .Y(_2089_) );
OR2X2 OR2X2_21 ( .A(_2089_), .B(_2086_), .Y(_2090_) );
NAND2X1 NAND2X1_315 ( .A(_2086_), .B(_2089_), .Y(_2091_) );
NAND3X1 NAND3X1_99 ( .A(micro_hash_ucr_pipe44_bF_buf1), .B(_2091_), .C(_2090_), .Y(_2092_) );
OAI21X1 OAI21X1_585 ( .A(_2084_), .B(micro_hash_ucr_pipe44_bF_buf1), .C(_2092_), .Y(_2093_) );
INVX4 INVX4_38 ( .A(micro_hash_ucr_Wx_158_), .Y(_2094_) );
XNOR2X1 XNOR2X1_136 ( .A(_1942__bF_buf3), .B(_2094_), .Y(_2095_) );
INVX1 INVX1_286 ( .A(_1699_), .Y(_2096_) );
OAI21X1 OAI21X1_586 ( .A(_1697_), .B(_2096_), .C(_1700_), .Y(_2097_) );
AND2X2 AND2X2_76 ( .A(_2097_), .B(_2095_), .Y(_2098_) );
NOR2X1 NOR2X1_459 ( .A(_2095_), .B(_2097_), .Y(_2099_) );
OAI21X1 OAI21X1_587 ( .A(_2098_), .B(_2099_), .C(micro_hash_ucr_pipe46_bF_buf2), .Y(_2100_) );
OAI21X1 OAI21X1_588 ( .A(_2093_), .B(micro_hash_ucr_pipe46_bF_buf2), .C(_2100_), .Y(_2101_) );
INVX4 INVX4_39 ( .A(micro_hash_ucr_Wx_166_), .Y(_2102_) );
XNOR2X1 XNOR2X1_137 ( .A(_1942__bF_buf3), .B(_2102_), .Y(_2103_) );
INVX1 INVX1_287 ( .A(micro_hash_ucr_Wx_165_), .Y(_2104_) );
OAI21X1 OAI21X1_589 ( .A(micro_hash_ucr_Wx_165_), .B(_1678__bF_buf1), .C(_1859_), .Y(_2105_) );
OAI21X1 OAI21X1_590 ( .A(_2104_), .B(_1679__bF_buf1), .C(_2105_), .Y(_2106_) );
XOR2X1 XOR2X1_33 ( .A(_2106_), .B(_2103_), .Y(_2107_) );
AOI21X1 AOI21X1_223 ( .A(micro_hash_ucr_pipe48_bF_buf1), .B(_2107_), .C(micro_hash_ucr_pipe50_bF_buf2), .Y(_2108_) );
OAI21X1 OAI21X1_591 ( .A(_2101_), .B(micro_hash_ucr_pipe48_bF_buf1), .C(_2108_), .Y(_2109_) );
INVX4 INVX4_40 ( .A(micro_hash_ucr_Wx_174_), .Y(_2110_) );
XNOR2X1 XNOR2X1_138 ( .A(_1942__bF_buf1), .B(_2110_), .Y(_2111_) );
INVX1 INVX1_288 ( .A(_1866_), .Y(_2112_) );
OAI21X1 OAI21X1_592 ( .A(_1864_), .B(_2112_), .C(_1867_), .Y(_2113_) );
XNOR2X1 XNOR2X1_139 ( .A(_2113_), .B(_2111_), .Y(_2114_) );
AOI21X1 AOI21X1_224 ( .A(micro_hash_ucr_pipe50_bF_buf2), .B(_2114_), .C(micro_hash_ucr_pipe52_bF_buf3), .Y(_2115_) );
INVX4 INVX4_41 ( .A(micro_hash_ucr_Wx_182_), .Y(_2116_) );
XNOR2X1 XNOR2X1_140 ( .A(_1942__bF_buf1), .B(_2116_), .Y(_2117_) );
AOI21X1 AOI21X1_225 ( .A(_1875_), .B(_1873_), .C(_1876_), .Y(_2118_) );
INVX1 INVX1_289 ( .A(_2118_), .Y(_2119_) );
NAND2X1 NAND2X1_316 ( .A(_2117_), .B(_2119_), .Y(_2120_) );
INVX1 INVX1_290 ( .A(_2120_), .Y(_2121_) );
OAI21X1 OAI21X1_593 ( .A(_2119_), .B(_2117_), .C(micro_hash_ucr_pipe52_bF_buf3), .Y(_2122_) );
OAI21X1 OAI21X1_594 ( .A(_2121_), .B(_2122_), .C(_742__bF_buf2), .Y(_2123_) );
AOI21X1 AOI21X1_226 ( .A(_2115_), .B(_2109_), .C(_2123_), .Y(_2124_) );
XNOR2X1 XNOR2X1_141 ( .A(_1942__bF_buf3), .B(micro_hash_ucr_Wx_190_), .Y(_2125_) );
INVX1 INVX1_291 ( .A(_1694_), .Y(_2126_) );
OAI21X1 OAI21X1_595 ( .A(_1690_), .B(_1693_), .C(_2126_), .Y(_2127_) );
XNOR2X1 XNOR2X1_142 ( .A(_2127_), .B(_2125_), .Y(_2128_) );
OAI21X1 OAI21X1_596 ( .A(_2128_), .B(_742__bF_buf3), .C(_832__bF_buf3), .Y(_2129_) );
XNOR2X1 XNOR2X1_143 ( .A(_1942__bF_buf1), .B(micro_hash_ucr_Wx_198_), .Y(_2130_) );
OAI21X1 OAI21X1_597 ( .A(_1885_), .B(_1679__bF_buf1), .C(_1884_), .Y(_2131_) );
OAI21X1 OAI21X1_598 ( .A(micro_hash_ucr_Wx_197_), .B(_1678__bF_buf5), .C(_2131_), .Y(_2132_) );
OR2X2 OR2X2_22 ( .A(_2132_), .B(_2130_), .Y(_2133_) );
AOI21X1 AOI21X1_227 ( .A(_2130_), .B(_2132_), .C(_832__bF_buf1), .Y(_2134_) );
AOI21X1 AOI21X1_228 ( .A(_2134_), .B(_2133_), .C(micro_hash_ucr_pipe58_bF_buf1), .Y(_2135_) );
OAI21X1 OAI21X1_599 ( .A(_2124_), .B(_2129_), .C(_2135_), .Y(_2136_) );
INVX2 INVX2_134 ( .A(micro_hash_ucr_Wx_206_), .Y(_2137_) );
XNOR2X1 XNOR2X1_144 ( .A(_1942__bF_buf3), .B(_2137_), .Y(_2138_) );
OAI21X1 OAI21X1_600 ( .A(_1891_), .B(_1892_), .C(_1894_), .Y(_2139_) );
XNOR2X1 XNOR2X1_145 ( .A(_2139_), .B(_2138_), .Y(_2140_) );
AOI21X1 AOI21X1_229 ( .A(micro_hash_ucr_pipe58_bF_buf1), .B(_2140_), .C(micro_hash_ucr_pipe60_bF_buf0), .Y(_2141_) );
INVX2 INVX2_135 ( .A(micro_hash_ucr_Wx_214_), .Y(_2142_) );
XNOR2X1 XNOR2X1_146 ( .A(_1942__bF_buf3), .B(_2142_), .Y(_2143_) );
OAI21X1 OAI21X1_601 ( .A(_1899_), .B(_1901_), .C(_1903_), .Y(_2144_) );
NAND2X1 NAND2X1_317 ( .A(_2143_), .B(_2144_), .Y(_2145_) );
INVX1 INVX1_292 ( .A(_2145_), .Y(_2146_) );
OAI21X1 OAI21X1_602 ( .A(_2144_), .B(_2143_), .C(micro_hash_ucr_pipe60_bF_buf2), .Y(_2147_) );
OAI21X1 OAI21X1_603 ( .A(_2146_), .B(_2147_), .C(_4207__bF_buf1), .Y(_2148_) );
AOI21X1 AOI21X1_230 ( .A(_2141_), .B(_2136_), .C(_2148_), .Y(_2149_) );
INVX2 INVX2_136 ( .A(micro_hash_ucr_Wx_222_), .Y(_2150_) );
XNOR2X1 XNOR2X1_147 ( .A(_1942__bF_buf1), .B(_2150_), .Y(_2151_) );
OAI21X1 OAI21X1_604 ( .A(_1684_), .B(_1685_), .C(_1687_), .Y(_2152_) );
XOR2X1 XOR2X1_34 ( .A(_2152_), .B(_2151_), .Y(_2153_) );
OAI21X1 OAI21X1_605 ( .A(_2153_), .B(_4207__bF_buf3), .C(_278__bF_buf2), .Y(_2154_) );
INVX2 INVX2_137 ( .A(micro_hash_ucr_Wx_230_), .Y(_2155_) );
XNOR2X1 XNOR2X1_148 ( .A(_1942__bF_buf1), .B(_2155_), .Y(_2156_) );
INVX1 INVX1_293 ( .A(_1916_), .Y(_2157_) );
OAI21X1 OAI21X1_606 ( .A(_1912_), .B(_1915_), .C(_2157_), .Y(_2158_) );
NAND2X1 NAND2X1_318 ( .A(_2156_), .B(_2158_), .Y(_2159_) );
OR2X2 OR2X2_23 ( .A(_2158_), .B(_2156_), .Y(_2160_) );
NAND3X1 NAND3X1_100 ( .A(micro_hash_ucr_pipe64_bF_buf3), .B(_2159_), .C(_2160_), .Y(_2161_) );
OAI21X1 OAI21X1_607 ( .A(_2149_), .B(_2154_), .C(_2161_), .Y(_2162_) );
XNOR2X1 XNOR2X1_149 ( .A(_1942__bF_buf0), .B(micro_hash_ucr_Wx_238_), .Y(_2163_) );
INVX1 INVX1_294 ( .A(micro_hash_ucr_Wx_237_), .Y(_2164_) );
OAI21X1 OAI21X1_608 ( .A(_2164_), .B(_1679__bF_buf0), .C(_1922_), .Y(_2165_) );
OAI21X1 OAI21X1_609 ( .A(micro_hash_ucr_Wx_237_), .B(_1678__bF_buf0), .C(_2165_), .Y(_2166_) );
AND2X2 AND2X2_77 ( .A(_2166_), .B(_2163_), .Y(_2167_) );
OAI21X1 OAI21X1_610 ( .A(_2166_), .B(_2163_), .C(micro_hash_ucr_pipe66_bF_buf3), .Y(_2168_) );
OAI21X1 OAI21X1_611 ( .A(_2167_), .B(_2168_), .C(_4199__bF_buf5), .Y(_2169_) );
AOI21X1 AOI21X1_231 ( .A(_1078__bF_buf3), .B(_2162_), .C(_2169_), .Y(_2170_) );
INVX2 INVX2_138 ( .A(micro_hash_ucr_Wx_246_), .Y(_2171_) );
XNOR2X1 XNOR2X1_150 ( .A(_1942__bF_buf5), .B(_2171_), .Y(_2172_) );
INVX1 INVX1_295 ( .A(_1680_), .Y(_2173_) );
OAI21X1 OAI21X1_612 ( .A(_1666_), .B(_1677_), .C(_2173_), .Y(_2174_) );
XOR2X1 XOR2X1_35 ( .A(_2174_), .B(_2172_), .Y(_2175_) );
OAI21X1 OAI21X1_613 ( .A(_2175_), .B(_4199__bF_buf5), .C(_344_), .Y(_2176_) );
INVX2 INVX2_139 ( .A(micro_hash_ucr_Wx_254_), .Y(_2177_) );
XNOR2X1 XNOR2X1_151 ( .A(_1942__bF_buf0), .B(_2177_), .Y(_2178_) );
AOI21X1 AOI21X1_232 ( .A(_1931_), .B(_1929_), .C(_1932_), .Y(_2179_) );
INVX2 INVX2_140 ( .A(_2179_), .Y(_2180_) );
NOR2X1 NOR2X1_460 ( .A(_287_), .B(_292__bF_buf10), .Y(_198_) );
INVX4 INVX4_42 ( .A(_198_), .Y(_2181_) );
AOI21X1 AOI21X1_233 ( .A(_2178_), .B(_2180_), .C(_2181_), .Y(_2182_) );
OAI21X1 OAI21X1_614 ( .A(_2178_), .B(_2180_), .C(_2182_), .Y(_2183_) );
OAI21X1 OAI21X1_615 ( .A(_2170_), .B(_2176_), .C(_2183_), .Y(_128__6_) );
INVX8 INVX8_67 ( .A(_1942__bF_buf1), .Y(_2184_) );
NAND2X1 NAND2X1_319 ( .A(_2172_), .B(_2174_), .Y(_2185_) );
OAI21X1 OAI21X1_616 ( .A(_2171_), .B(_2184__bF_buf1), .C(_2185_), .Y(_2186_) );
NAND2X1 NAND2X1_320 ( .A(micro_hash_ucr_k_6_), .B(micro_hash_ucr_x_6_), .Y(_2187_) );
NAND2X1 NAND2X1_321 ( .A(_2187_), .B(_1940_), .Y(_2188_) );
XOR2X1 XOR2X1_36 ( .A(micro_hash_ucr_k_7_), .B(micro_hash_ucr_x_7_), .Y(_2189_) );
XOR2X1 XOR2X1_37 ( .A(_2188_), .B(_2189_), .Y(_2190_) );
XNOR2X1 XNOR2X1_152 ( .A(_2190__bF_buf2), .B(micro_hash_ucr_Wx_247_), .Y(_2191_) );
AND2X2 AND2X2_78 ( .A(_2186_), .B(_2191_), .Y(_2192_) );
NAND2X1 NAND2X1_322 ( .A(_2151_), .B(_2152_), .Y(_2193_) );
OAI21X1 OAI21X1_617 ( .A(_2150_), .B(_2184__bF_buf2), .C(_2193_), .Y(_2194_) );
XNOR2X1 XNOR2X1_153 ( .A(_2190__bF_buf2), .B(micro_hash_ucr_Wx_223_), .Y(_2195_) );
XNOR2X1 XNOR2X1_154 ( .A(_2194_), .B(_2195_), .Y(_2196_) );
NAND2X1 NAND2X1_323 ( .A(_2111_), .B(_2113_), .Y(_2197_) );
OAI21X1 OAI21X1_618 ( .A(_2110_), .B(_2184__bF_buf2), .C(_2197_), .Y(_2198_) );
XNOR2X1 XNOR2X1_155 ( .A(_2190__bF_buf0), .B(micro_hash_ucr_Wx_175_), .Y(_2199_) );
XNOR2X1 XNOR2X1_156 ( .A(_2198_), .B(_2199_), .Y(_2200_) );
OAI21X1 OAI21X1_619 ( .A(_2052_), .B(_2184__bF_buf1), .C(_2058_), .Y(_2201_) );
XNOR2X1 XNOR2X1_157 ( .A(_2190__bF_buf0), .B(micro_hash_ucr_Wx_119_), .Y(_2202_) );
XNOR2X1 XNOR2X1_158 ( .A(_2201_), .B(_2202_), .Y(_2203_) );
INVX2 INVX2_141 ( .A(micro_hash_ucr_Wx_78_), .Y(_2204_) );
OAI21X1 OAI21X1_620 ( .A(_2204_), .B(_2184__bF_buf3), .C(_2014_), .Y(_2205_) );
XNOR2X1 XNOR2X1_159 ( .A(_2190__bF_buf4), .B(micro_hash_ucr_Wx_79_), .Y(_2206_) );
XNOR2X1 XNOR2X1_160 ( .A(_2205_), .B(_2206_), .Y(_2207_) );
INVX1 INVX1_296 ( .A(H_23_), .Y(_2208_) );
AOI21X1 AOI21X1_234 ( .A(micro_hash_ucr_c_7_), .B(_4252_), .C(micro_hash_ucr_pipe8), .Y(_2209_) );
OAI21X1 OAI21X1_621 ( .A(_4252_), .B(_2208_), .C(_2209_), .Y(_2210_) );
NAND2X1 NAND2X1_324 ( .A(_1947_), .B(_1949_), .Y(_2211_) );
OAI21X1 OAI21X1_622 ( .A(_1946_), .B(_2184__bF_buf3), .C(_2211_), .Y(_2212_) );
XNOR2X1 XNOR2X1_161 ( .A(_2190__bF_buf1), .B(micro_hash_ucr_Wx_7_), .Y(_2213_) );
AND2X2 AND2X2_79 ( .A(_2212_), .B(_2213_), .Y(_2214_) );
OAI21X1 OAI21X1_623 ( .A(_2212_), .B(_2213_), .C(micro_hash_ucr_pipe8), .Y(_2215_) );
OAI21X1 OAI21X1_624 ( .A(_2214_), .B(_2215_), .C(_2210_), .Y(_2216_) );
NAND2X1 NAND2X1_325 ( .A(micro_hash_ucr_Wx_14_), .B(_1942__bF_buf4), .Y(_2217_) );
INVX1 INVX1_297 ( .A(_1944_), .Y(_2218_) );
OAI21X1 OAI21X1_625 ( .A(_2218_), .B(_1943_), .C(_2217_), .Y(_2219_) );
XOR2X1 XOR2X1_38 ( .A(_2190__bF_buf3), .B(micro_hash_ucr_Wx_15_), .Y(_2220_) );
XNOR2X1 XNOR2X1_162 ( .A(_2219_), .B(_2220_), .Y(_2221_) );
MUX2X1 MUX2X1_47 ( .A(_2216_), .B(_2221_), .S(_4243_), .Y(_2222_) );
NAND2X1 NAND2X1_326 ( .A(_4258_), .B(_2222_), .Y(_2223_) );
NAND2X1 NAND2X1_327 ( .A(_1958_), .B(_1960_), .Y(_2224_) );
OAI21X1 OAI21X1_626 ( .A(_1957_), .B(_2184__bF_buf3), .C(_2224_), .Y(_2225_) );
XNOR2X1 XNOR2X1_163 ( .A(_2190__bF_buf3), .B(micro_hash_ucr_Wx_23_), .Y(_2226_) );
XNOR2X1 XNOR2X1_164 ( .A(_2225_), .B(_2226_), .Y(_2227_) );
AOI21X1 AOI21X1_235 ( .A(micro_hash_ucr_pipe12_bF_buf2), .B(_2227_), .C(micro_hash_ucr_pipe14), .Y(_2228_) );
NAND2X1 NAND2X1_328 ( .A(_1964_), .B(_1966_), .Y(_2229_) );
OAI21X1 OAI21X1_627 ( .A(_1963_), .B(_2184__bF_buf3), .C(_2229_), .Y(_2230_) );
INVX2 INVX2_142 ( .A(micro_hash_ucr_Wx_31_), .Y(_2231_) );
XNOR2X1 XNOR2X1_165 ( .A(_2190__bF_buf3), .B(_2231_), .Y(_2232_) );
XNOR2X1 XNOR2X1_166 ( .A(_2230_), .B(_2232_), .Y(_2233_) );
AOI22X1 AOI22X1_14 ( .A(micro_hash_ucr_pipe14), .B(_2233_), .C(_2223_), .D(_2228_), .Y(_2234_) );
NOR2X1 NOR2X1_461 ( .A(micro_hash_ucr_pipe16), .B(_2234_), .Y(_2235_) );
NAND2X1 NAND2X1_329 ( .A(_1971_), .B(_1974_), .Y(_2236_) );
OAI21X1 OAI21X1_628 ( .A(_1970_), .B(_2184__bF_buf3), .C(_2236_), .Y(_2237_) );
XNOR2X1 XNOR2X1_167 ( .A(_2190__bF_buf4), .B(micro_hash_ucr_Wx_39_), .Y(_2238_) );
OAI21X1 OAI21X1_629 ( .A(_2237_), .B(_2238_), .C(micro_hash_ucr_pipe16), .Y(_2239_) );
AOI21X1 AOI21X1_236 ( .A(_2237_), .B(_2238_), .C(_2239_), .Y(_2240_) );
NOR2X1 NOR2X1_462 ( .A(_2240_), .B(_2235_), .Y(_2241_) );
AOI21X1 AOI21X1_237 ( .A(micro_hash_ucr_Wx_46_), .B(_1942__bF_buf2), .C(_1982_), .Y(_2242_) );
XNOR2X1 XNOR2X1_168 ( .A(_2190__bF_buf4), .B(micro_hash_ucr_Wx_47_), .Y(_2243_) );
AND2X2 AND2X2_80 ( .A(_2242_), .B(_2243_), .Y(_2244_) );
OAI21X1 OAI21X1_630 ( .A(_2242_), .B(_2243_), .C(micro_hash_ucr_pipe18_bF_buf2), .Y(_2245_) );
OAI21X1 OAI21X1_631 ( .A(_2244_), .B(_2245_), .C(_4237__bF_buf4), .Y(_2246_) );
AOI21X1 AOI21X1_238 ( .A(_624__bF_buf3), .B(_2241_), .C(_2246_), .Y(_2247_) );
OAI21X1 OAI21X1_632 ( .A(_1985_), .B(_2184__bF_buf1), .C(_1989_), .Y(_2248_) );
XNOR2X1 XNOR2X1_169 ( .A(_2190__bF_buf4), .B(micro_hash_ucr_Wx_55_), .Y(_2249_) );
OAI21X1 OAI21X1_633 ( .A(_2248_), .B(_2249_), .C(micro_hash_ucr_pipe20_bF_buf1), .Y(_2250_) );
AOI21X1 AOI21X1_239 ( .A(_2248_), .B(_2249_), .C(_2250_), .Y(_2251_) );
NOR2X1 NOR2X1_463 ( .A(_2251_), .B(_2247_), .Y(_2252_) );
OAI21X1 OAI21X1_634 ( .A(_1994_), .B(_2184__bF_buf3), .C(_2000_), .Y(_2253_) );
INVX2 INVX2_143 ( .A(micro_hash_ucr_Wx_63_), .Y(_2254_) );
XNOR2X1 XNOR2X1_170 ( .A(_2190__bF_buf3), .B(_2254_), .Y(_2255_) );
XNOR2X1 XNOR2X1_171 ( .A(_2253_), .B(_2255_), .Y(_2256_) );
OAI21X1 OAI21X1_635 ( .A(_2256_), .B(_4262__bF_buf1), .C(_4233__bF_buf1), .Y(_2257_) );
AOI21X1 AOI21X1_240 ( .A(_4262__bF_buf1), .B(_2252_), .C(_2257_), .Y(_2258_) );
OAI21X1 OAI21X1_636 ( .A(_2003_), .B(_2184__bF_buf1), .C(_2008_), .Y(_2259_) );
XNOR2X1 XNOR2X1_172 ( .A(_2190__bF_buf2), .B(micro_hash_ucr_Wx_71_), .Y(_2260_) );
OAI21X1 OAI21X1_637 ( .A(_2259_), .B(_2260_), .C(micro_hash_ucr_pipe24_bF_buf0), .Y(_2261_) );
AOI21X1 AOI21X1_241 ( .A(_2259_), .B(_2260_), .C(_2261_), .Y(_2262_) );
OAI21X1 OAI21X1_638 ( .A(_2258_), .B(_2262_), .C(_4230__bF_buf3), .Y(_2263_) );
OAI21X1 OAI21X1_639 ( .A(_4230__bF_buf3), .B(_2207_), .C(_2263_), .Y(_2264_) );
OAI21X1 OAI21X1_640 ( .A(_2019_), .B(_2184__bF_buf1), .C(_2025_), .Y(_2265_) );
INVX2 INVX2_144 ( .A(micro_hash_ucr_Wx_87_), .Y(_2266_) );
XNOR2X1 XNOR2X1_173 ( .A(_2190__bF_buf4), .B(_2266_), .Y(_2267_) );
XNOR2X1 XNOR2X1_174 ( .A(_2265_), .B(_2267_), .Y(_2268_) );
MUX2X1 MUX2X1_48 ( .A(_2264_), .B(_2268_), .S(_220__bF_buf3), .Y(_2269_) );
AOI21X1 AOI21X1_242 ( .A(micro_hash_ucr_Wx_94_), .B(_1942__bF_buf4), .C(_2032_), .Y(_2270_) );
INVX2 INVX2_145 ( .A(micro_hash_ucr_Wx_95_), .Y(_2271_) );
XNOR2X1 XNOR2X1_175 ( .A(_2190__bF_buf0), .B(_2271_), .Y(_2272_) );
AOI21X1 AOI21X1_243 ( .A(_2272_), .B(_2270_), .C(_4228__bF_buf3), .Y(_2273_) );
OAI21X1 OAI21X1_641 ( .A(_2270_), .B(_2272_), .C(_2273_), .Y(_2274_) );
OAI21X1 OAI21X1_642 ( .A(_2269_), .B(micro_hash_ucr_pipe30_bF_buf2), .C(_2274_), .Y(_2275_) );
OAI21X1 OAI21X1_643 ( .A(_2036_), .B(_2184__bF_buf1), .C(_2041_), .Y(_2276_) );
INVX2 INVX2_146 ( .A(micro_hash_ucr_Wx_103_), .Y(_2277_) );
XNOR2X1 XNOR2X1_176 ( .A(_2190__bF_buf3), .B(_2277_), .Y(_2278_) );
XNOR2X1 XNOR2X1_177 ( .A(_2276_), .B(_2278_), .Y(_2279_) );
MUX2X1 MUX2X1_49 ( .A(_2275_), .B(_2279_), .S(_4226__bF_buf2), .Y(_2280_) );
AOI21X1 AOI21X1_244 ( .A(micro_hash_ucr_Wx_110_), .B(_1942__bF_buf5), .C(_2048_), .Y(_2281_) );
INVX4 INVX4_43 ( .A(micro_hash_ucr_Wx_111_), .Y(_2282_) );
XNOR2X1 XNOR2X1_178 ( .A(_2190__bF_buf4), .B(_2282_), .Y(_2283_) );
AOI21X1 AOI21X1_245 ( .A(_2283_), .B(_2281_), .C(_4225__bF_buf1), .Y(_2284_) );
OAI21X1 OAI21X1_644 ( .A(_2281_), .B(_2283_), .C(_2284_), .Y(_2285_) );
OAI21X1 OAI21X1_645 ( .A(_2280_), .B(micro_hash_ucr_pipe34_bF_buf0), .C(_2285_), .Y(_2286_) );
NAND2X1 NAND2X1_330 ( .A(_4224__bF_buf1), .B(_2286_), .Y(_2287_) );
OAI21X1 OAI21X1_646 ( .A(_4224__bF_buf1), .B(_2203_), .C(_2287_), .Y(_2288_) );
OAI21X1 OAI21X1_647 ( .A(_2062_), .B(_2184__bF_buf2), .C(_2066_), .Y(_2289_) );
XNOR2X1 XNOR2X1_179 ( .A(_2190__bF_buf4), .B(micro_hash_ucr_Wx_127_), .Y(_2290_) );
XNOR2X1 XNOR2X1_180 ( .A(_2289_), .B(_2290_), .Y(_2291_) );
OAI21X1 OAI21X1_648 ( .A(_2291_), .B(_701__bF_buf4), .C(_296__bF_buf4), .Y(_2292_) );
AOI21X1 AOI21X1_246 ( .A(_701__bF_buf4), .B(_2288_), .C(_2292_), .Y(_2293_) );
OAI21X1 OAI21X1_649 ( .A(_2069_), .B(_2184__bF_buf2), .C(_2074_), .Y(_2294_) );
INVX4 INVX4_44 ( .A(micro_hash_ucr_Wx_135_), .Y(_2295_) );
XNOR2X1 XNOR2X1_181 ( .A(_2190__bF_buf2), .B(_2295_), .Y(_2296_) );
XNOR2X1 XNOR2X1_182 ( .A(_2294_), .B(_2296_), .Y(_2297_) );
OAI21X1 OAI21X1_650 ( .A(_2297_), .B(_296__bF_buf4), .C(_4220__bF_buf4), .Y(_2298_) );
AOI21X1 AOI21X1_247 ( .A(micro_hash_ucr_Wx_142_), .B(_1942__bF_buf0), .C(_2081_), .Y(_2299_) );
INVX2 INVX2_147 ( .A(micro_hash_ucr_Wx_143_), .Y(_2300_) );
XNOR2X1 XNOR2X1_183 ( .A(_2190__bF_buf3), .B(_2300_), .Y(_2301_) );
AOI21X1 AOI21X1_248 ( .A(_2301_), .B(_2299_), .C(_4220__bF_buf4), .Y(_2302_) );
OAI21X1 OAI21X1_651 ( .A(_2299_), .B(_2301_), .C(_2302_), .Y(_2303_) );
OAI21X1 OAI21X1_652 ( .A(_2293_), .B(_2298_), .C(_2303_), .Y(_2304_) );
OAI21X1 OAI21X1_653 ( .A(_2085_), .B(_2184__bF_buf0), .C(_2091_), .Y(_2305_) );
XNOR2X1 XNOR2X1_184 ( .A(_2190__bF_buf3), .B(micro_hash_ucr_Wx_151_), .Y(_2306_) );
OAI21X1 OAI21X1_654 ( .A(_2305_), .B(_2306_), .C(micro_hash_ucr_pipe44_bF_buf1), .Y(_2307_) );
AOI21X1 AOI21X1_249 ( .A(_2305_), .B(_2306_), .C(_2307_), .Y(_2308_) );
AOI21X1 AOI21X1_250 ( .A(_4219__bF_buf1), .B(_2304_), .C(_2308_), .Y(_2309_) );
AOI21X1 AOI21X1_251 ( .A(micro_hash_ucr_Wx_158_), .B(_1942__bF_buf3), .C(_2098_), .Y(_2310_) );
XNOR2X1 XNOR2X1_185 ( .A(_2190__bF_buf1), .B(micro_hash_ucr_Wx_159_), .Y(_2311_) );
AND2X2 AND2X2_81 ( .A(_2310_), .B(_2311_), .Y(_2312_) );
OAI21X1 OAI21X1_655 ( .A(_2310_), .B(_2311_), .C(micro_hash_ucr_pipe46_bF_buf2), .Y(_2313_) );
OAI21X1 OAI21X1_656 ( .A(_2312_), .B(_2313_), .C(_4217__bF_buf2), .Y(_2314_) );
AOI21X1 AOI21X1_252 ( .A(_4218__bF_buf3), .B(_2309_), .C(_2314_), .Y(_2315_) );
NAND2X1 NAND2X1_331 ( .A(_2103_), .B(_2106_), .Y(_2316_) );
OAI21X1 OAI21X1_657 ( .A(_2102_), .B(_2184__bF_buf0), .C(_2316_), .Y(_2317_) );
XNOR2X1 XNOR2X1_186 ( .A(_2190__bF_buf0), .B(micro_hash_ucr_Wx_167_), .Y(_2318_) );
OAI21X1 OAI21X1_658 ( .A(_2317_), .B(_2318_), .C(micro_hash_ucr_pipe48_bF_buf1), .Y(_2319_) );
AOI21X1 AOI21X1_253 ( .A(_2317_), .B(_2318_), .C(_2319_), .Y(_2320_) );
OAI21X1 OAI21X1_659 ( .A(_2315_), .B(_2320_), .C(_4215__bF_buf4), .Y(_2321_) );
OAI21X1 OAI21X1_660 ( .A(_4215__bF_buf4), .B(_2200_), .C(_2321_), .Y(_2322_) );
OAI21X1 OAI21X1_661 ( .A(_2116_), .B(_2184__bF_buf0), .C(_2120_), .Y(_2323_) );
INVX4 INVX4_45 ( .A(micro_hash_ucr_Wx_183_), .Y(_2324_) );
XNOR2X1 XNOR2X1_187 ( .A(_2190__bF_buf1), .B(_2324_), .Y(_2325_) );
XNOR2X1 XNOR2X1_188 ( .A(_2323_), .B(_2325_), .Y(_2326_) );
MUX2X1 MUX2X1_50 ( .A(_2322_), .B(_2326_), .S(_4214__bF_buf3), .Y(_2327_) );
INVX1 INVX1_298 ( .A(_2127_), .Y(_2328_) );
NOR2X1 NOR2X1_464 ( .A(_2125_), .B(_2328_), .Y(_2329_) );
AOI21X1 AOI21X1_254 ( .A(micro_hash_ucr_Wx_190_), .B(_1942__bF_buf3), .C(_2329_), .Y(_2330_) );
XOR2X1 XOR2X1_39 ( .A(_2190__bF_buf0), .B(micro_hash_ucr_Wx_191_), .Y(_2331_) );
AOI21X1 AOI21X1_255 ( .A(_2331_), .B(_2330_), .C(_742__bF_buf2), .Y(_2332_) );
OAI21X1 OAI21X1_662 ( .A(_2330_), .B(_2331_), .C(_2332_), .Y(_2333_) );
OAI21X1 OAI21X1_663 ( .A(_2327_), .B(micro_hash_ucr_pipe54_bF_buf2), .C(_2333_), .Y(_2334_) );
INVX1 INVX1_299 ( .A(micro_hash_ucr_Wx_198_), .Y(_2335_) );
OAI21X1 OAI21X1_664 ( .A(_2335_), .B(_2184__bF_buf0), .C(_2133_), .Y(_2336_) );
XNOR2X1 XNOR2X1_189 ( .A(_2190__bF_buf2), .B(micro_hash_ucr_Wx_199_), .Y(_2337_) );
OAI21X1 OAI21X1_665 ( .A(_2336_), .B(_2337_), .C(micro_hash_ucr_pipe56_bF_buf3), .Y(_2338_) );
AOI21X1 AOI21X1_256 ( .A(_2336_), .B(_2337_), .C(_2338_), .Y(_2339_) );
AOI21X1 AOI21X1_257 ( .A(_832__bF_buf1), .B(_2334_), .C(_2339_), .Y(_2340_) );
NAND2X1 NAND2X1_332 ( .A(_2138_), .B(_2139_), .Y(_2341_) );
OAI21X1 OAI21X1_666 ( .A(_2137_), .B(_2184__bF_buf0), .C(_2341_), .Y(_2342_) );
XOR2X1 XOR2X1_40 ( .A(_2190__bF_buf1), .B(micro_hash_ucr_Wx_207_), .Y(_2343_) );
XNOR2X1 XNOR2X1_190 ( .A(_2342_), .B(_2343_), .Y(_2344_) );
OAI21X1 OAI21X1_667 ( .A(_2344_), .B(_4211__bF_buf3), .C(_4210__bF_buf4), .Y(_2345_) );
AOI21X1 AOI21X1_258 ( .A(_4211__bF_buf3), .B(_2340_), .C(_2345_), .Y(_2346_) );
OAI21X1 OAI21X1_668 ( .A(_2142_), .B(_2184__bF_buf0), .C(_2145_), .Y(_2347_) );
XNOR2X1 XNOR2X1_191 ( .A(_2190__bF_buf0), .B(micro_hash_ucr_Wx_215_), .Y(_2348_) );
OAI21X1 OAI21X1_669 ( .A(_2347_), .B(_2348_), .C(micro_hash_ucr_pipe60_bF_buf2), .Y(_2349_) );
AOI21X1 AOI21X1_259 ( .A(_2347_), .B(_2348_), .C(_2349_), .Y(_2350_) );
OAI21X1 OAI21X1_670 ( .A(_2346_), .B(_2350_), .C(_4207__bF_buf1), .Y(_2351_) );
OAI21X1 OAI21X1_671 ( .A(_4207__bF_buf3), .B(_2196_), .C(_2351_), .Y(_2352_) );
OAI21X1 OAI21X1_672 ( .A(_2155_), .B(_2184__bF_buf2), .C(_2159_), .Y(_2353_) );
XOR2X1 XOR2X1_41 ( .A(_2190__bF_buf1), .B(micro_hash_ucr_Wx_231_), .Y(_2354_) );
XNOR2X1 XNOR2X1_192 ( .A(_2353_), .B(_2354_), .Y(_2355_) );
MUX2X1 MUX2X1_51 ( .A(_2352_), .B(_2355_), .S(_278__bF_buf2), .Y(_2356_) );
NOR2X1 NOR2X1_465 ( .A(_2163_), .B(_2166_), .Y(_2357_) );
AOI21X1 AOI21X1_260 ( .A(micro_hash_ucr_Wx_238_), .B(_1942__bF_buf0), .C(_2357_), .Y(_2358_) );
XOR2X1 XOR2X1_42 ( .A(_2190__bF_buf2), .B(micro_hash_ucr_Wx_239_), .Y(_2359_) );
AOI21X1 AOI21X1_261 ( .A(_2359_), .B(_2358_), .C(_1078__bF_buf3), .Y(_2360_) );
OAI21X1 OAI21X1_673 ( .A(_2358_), .B(_2359_), .C(_2360_), .Y(_2361_) );
OAI21X1 OAI21X1_674 ( .A(_2356_), .B(micro_hash_ucr_pipe66_bF_buf3), .C(_2361_), .Y(_2362_) );
NAND2X1 NAND2X1_333 ( .A(_4199__bF_buf5), .B(_2362_), .Y(_2363_) );
OAI21X1 OAI21X1_675 ( .A(_2186_), .B(_2191_), .C(micro_hash_ucr_pipe68), .Y(_2364_) );
OAI21X1 OAI21X1_676 ( .A(_2192_), .B(_2364_), .C(_2363_), .Y(_2365_) );
NAND2X1 NAND2X1_334 ( .A(_2178_), .B(_2180_), .Y(_2366_) );
OAI21X1 OAI21X1_677 ( .A(_2177_), .B(_2184__bF_buf2), .C(_2366_), .Y(_2367_) );
XNOR2X1 XNOR2X1_193 ( .A(_2190__bF_buf1), .B(micro_hash_ucr_Wx_255_), .Y(_2368_) );
AND2X2 AND2X2_82 ( .A(_2367_), .B(_2368_), .Y(_2369_) );
OAI21X1 OAI21X1_678 ( .A(_2367_), .B(_2368_), .C(micro_hash_ucr_pipe69), .Y(_2370_) );
OAI21X1 OAI21X1_679 ( .A(_2369_), .B(_2370_), .C(_131__bF_buf13), .Y(_2371_) );
AOI21X1 AOI21X1_262 ( .A(_287_), .B(_2365_), .C(_2371_), .Y(_128__7_) );
OAI21X1 OAI21X1_680 ( .A(comparador_valid_hash), .B(micro_hash_ucr_pipe70_bF_buf1), .C(_131__bF_buf6), .Y(_2372_) );
NOR2X1 NOR2X1_466 ( .A(micro_hash_ucr_pipe71), .B(_2372_), .Y(_203_) );
AOI21X1 AOI21X1_263 ( .A(micro_hash_ucr_Wx_176_), .B(_523_), .C(micro_hash_ucr_Wx_224_), .Y(_2373_) );
OAI21X1 OAI21X1_681 ( .A(_523_), .B(micro_hash_ucr_Wx_176_), .C(_2373_), .Y(_2374_) );
AND2X2 AND2X2_83 ( .A(_2374_), .B(_131__bF_buf3), .Y(_125__248_) );
OAI21X1 OAI21X1_682 ( .A(_715_), .B(micro_hash_ucr_Wx_177_), .C(_787_), .Y(_2375_) );
AOI21X1 AOI21X1_264 ( .A(_715_), .B(micro_hash_ucr_Wx_177_), .C(_2375_), .Y(_2376_) );
NOR2X1 NOR2X1_467 ( .A(_2376_), .B(_292__bF_buf8), .Y(_125__249_) );
OAI21X1 OAI21X1_683 ( .A(_991_), .B(micro_hash_ucr_Wx_178_), .C(_1081_), .Y(_2377_) );
AOI21X1 AOI21X1_265 ( .A(_991_), .B(micro_hash_ucr_Wx_178_), .C(_2377_), .Y(_2378_) );
NOR2X1 NOR2X1_468 ( .A(_2378_), .B(_292__bF_buf3), .Y(_125__250_) );
OAI21X1 OAI21X1_684 ( .A(_1319_), .B(micro_hash_ucr_Wx_179_), .C(_1402_), .Y(_2379_) );
AOI21X1 AOI21X1_266 ( .A(_1319_), .B(micro_hash_ucr_Wx_179_), .C(_2379_), .Y(_2380_) );
NOR2X1 NOR2X1_469 ( .A(_2380_), .B(_292__bF_buf12), .Y(_125__251_) );
AOI21X1 AOI21X1_267 ( .A(micro_hash_ucr_Wx_180_), .B(_1563_), .C(micro_hash_ucr_Wx_228_), .Y(_2381_) );
OAI21X1 OAI21X1_685 ( .A(_1563_), .B(micro_hash_ucr_Wx_180_), .C(_2381_), .Y(_2382_) );
AND2X2 AND2X2_84 ( .A(_2382_), .B(_131__bF_buf10), .Y(_125__252_) );
OAI21X1 OAI21X1_686 ( .A(_2078_), .B(micro_hash_ucr_Wx_181_), .C(_1913_), .Y(_2383_) );
AOI21X1 AOI21X1_268 ( .A(_2078_), .B(micro_hash_ucr_Wx_181_), .C(_2383_), .Y(_2384_) );
NOR2X1 NOR2X1_470 ( .A(_2384_), .B(_292__bF_buf11), .Y(_125__253_) );
OAI21X1 OAI21X1_687 ( .A(_2116_), .B(micro_hash_ucr_Wx_142_), .C(_2155_), .Y(_2385_) );
AOI21X1 AOI21X1_269 ( .A(_2116_), .B(micro_hash_ucr_Wx_142_), .C(_2385_), .Y(_2386_) );
NOR2X1 NOR2X1_471 ( .A(_2386_), .B(_292__bF_buf5), .Y(_125__254_) );
AOI21X1 AOI21X1_270 ( .A(micro_hash_ucr_Wx_143_), .B(_2324_), .C(micro_hash_ucr_Wx_231_), .Y(_2387_) );
OAI21X1 OAI21X1_688 ( .A(_2324_), .B(micro_hash_ucr_Wx_143_), .C(_2387_), .Y(_2388_) );
AND2X2 AND2X2_85 ( .A(_2388_), .B(_131__bF_buf13), .Y(_125__255_) );
NOR2X1 NOR2X1_472 ( .A(micro_hash_ucr_pipe70_bF_buf3), .B(micro_hash_ucr_pipe5), .Y(_2389_) );
NAND2X1 NAND2X1_335 ( .A(H_16_), .B(_2389_), .Y(_2390_) );
INVX8 INVX8_68 ( .A(micro_hash_ucr_c_0_bF_buf2_), .Y(_2391_) );
OAI21X1 OAI21X1_689 ( .A(_443_), .B(_2391_), .C(micro_hash_ucr_pipe70_bF_buf3), .Y(_2392_) );
OAI21X1 OAI21X1_690 ( .A(H_16_), .B(micro_hash_ucr_c_0_bF_buf1_), .C(_131__bF_buf13), .Y(_2393_) );
AOI21X1 AOI21X1_271 ( .A(_2390_), .B(_2392_), .C(_2393_), .Y(_129__16_) );
NOR2X1 NOR2X1_473 ( .A(_443_), .B(_2391_), .Y(_2394_) );
NOR2X1 NOR2X1_474 ( .A(H_17_), .B(micro_hash_ucr_c_1_bF_buf2_), .Y(_2395_) );
NOR2X1 NOR2X1_475 ( .A(_593_), .B(_591__bF_buf3), .Y(_2396_) );
NOR2X1 NOR2X1_476 ( .A(_2395_), .B(_2396_), .Y(_2397_) );
XNOR2X1 XNOR2X1_194 ( .A(_2397_), .B(_2394_), .Y(_2398_) );
INVX8 INVX8_69 ( .A(_2389_), .Y(_2399_) );
OAI21X1 OAI21X1_691 ( .A(H_17_), .B(_2399_), .C(_131__bF_buf13), .Y(_2400_) );
AOI21X1 AOI21X1_272 ( .A(micro_hash_ucr_pipe70_bF_buf1), .B(_2398_), .C(_2400_), .Y(_129__17_) );
NAND2X1 NAND2X1_336 ( .A(_2394_), .B(_2397_), .Y(_2401_) );
OAI21X1 OAI21X1_692 ( .A(_593_), .B(_591__bF_buf3), .C(_2401_), .Y(_2402_) );
XOR2X1 XOR2X1_43 ( .A(H_18_), .B(micro_hash_ucr_c_2_bF_buf2_), .Y(_2403_) );
XNOR2X1 XNOR2X1_195 ( .A(_2402_), .B(_2403_), .Y(_2404_) );
OAI21X1 OAI21X1_693 ( .A(H_18_), .B(_2399_), .C(_131__bF_buf6), .Y(_2405_) );
AOI21X1 AOI21X1_273 ( .A(micro_hash_ucr_pipe70_bF_buf1), .B(_2404_), .C(_2405_), .Y(_129__18_) );
INVX1 INVX1_300 ( .A(_2402_), .Y(_2406_) );
INVX1 INVX1_301 ( .A(_2403_), .Y(_2407_) );
NOR2X1 NOR2X1_477 ( .A(_2407_), .B(_2406_), .Y(_2408_) );
AOI21X1 AOI21X1_274 ( .A(H_18_), .B(micro_hash_ucr_c_2_bF_buf1_), .C(_2408_), .Y(_2409_) );
NOR2X1 NOR2X1_478 ( .A(micro_hash_ucr_c_3_bF_buf3_), .B(H_19_), .Y(_2410_) );
NOR2X1 NOR2X1_479 ( .A(_4200_), .B(_1184_), .Y(_2411_) );
OR2X2 OR2X2_24 ( .A(_2411_), .B(_2410_), .Y(_2412_) );
XNOR2X1 XNOR2X1_196 ( .A(_2409_), .B(_2412_), .Y(_2413_) );
OAI21X1 OAI21X1_694 ( .A(H_19_), .B(_2399_), .C(_131__bF_buf13), .Y(_2414_) );
AOI21X1 AOI21X1_275 ( .A(micro_hash_ucr_pipe70_bF_buf2), .B(_2413_), .C(_2414_), .Y(_129__19_) );
NOR2X1 NOR2X1_480 ( .A(H_20_), .B(micro_hash_ucr_c_4_), .Y(_2415_) );
AND2X2 AND2X2_86 ( .A(H_20_), .B(micro_hash_ucr_c_4_), .Y(_2416_) );
NOR2X1 NOR2X1_481 ( .A(_2415_), .B(_2416_), .Y(_2417_) );
INVX1 INVX1_302 ( .A(_2411_), .Y(_2418_) );
OAI21X1 OAI21X1_695 ( .A(_2409_), .B(_2410_), .C(_2418_), .Y(_2419_) );
XNOR2X1 XNOR2X1_197 ( .A(_2419_), .B(_2417_), .Y(_2420_) );
OAI21X1 OAI21X1_696 ( .A(H_20_), .B(_2399_), .C(_131__bF_buf6), .Y(_2421_) );
AOI21X1 AOI21X1_276 ( .A(micro_hash_ucr_pipe70_bF_buf2), .B(_2420_), .C(_2421_), .Y(_129__20_) );
AOI21X1 AOI21X1_277 ( .A(_2417_), .B(_2419_), .C(_2416_), .Y(_2422_) );
NOR2X1 NOR2X1_482 ( .A(H_21_), .B(micro_hash_ucr_c_5_), .Y(_2423_) );
NOR2X1 NOR2X1_483 ( .A(_1727_), .B(_1729_), .Y(_2424_) );
NOR2X1 NOR2X1_484 ( .A(_2423_), .B(_2424_), .Y(_2425_) );
OAI21X1 OAI21X1_697 ( .A(_2422_), .B(_2425_), .C(micro_hash_ucr_pipe70_bF_buf2), .Y(_2426_) );
AOI21X1 AOI21X1_278 ( .A(_2422_), .B(_2425_), .C(_2426_), .Y(_2427_) );
OAI21X1 OAI21X1_698 ( .A(H_21_), .B(_2399_), .C(_131__bF_buf6), .Y(_2428_) );
NOR2X1 NOR2X1_485 ( .A(_2428_), .B(_2427_), .Y(_129__21_) );
XOR2X1 XOR2X1_44 ( .A(H_22_), .B(micro_hash_ucr_c_6_), .Y(_2429_) );
INVX1 INVX1_303 ( .A(_2424_), .Y(_2430_) );
OAI21X1 OAI21X1_699 ( .A(_2422_), .B(_2423_), .C(_2430_), .Y(_2431_) );
XNOR2X1 XNOR2X1_198 ( .A(_2431_), .B(_2429_), .Y(_2432_) );
OAI21X1 OAI21X1_700 ( .A(H_22_), .B(_2399_), .C(_131__bF_buf6), .Y(_2433_) );
AOI21X1 AOI21X1_279 ( .A(micro_hash_ucr_pipe70_bF_buf2), .B(_2432_), .C(_2433_), .Y(_129__22_) );
INVX1 INVX1_304 ( .A(micro_hash_ucr_c_6_), .Y(_2434_) );
NAND2X1 NAND2X1_337 ( .A(_2429_), .B(_2431_), .Y(_2435_) );
OAI21X1 OAI21X1_701 ( .A(_1952_), .B(_2434_), .C(_2435_), .Y(_2436_) );
XOR2X1 XOR2X1_45 ( .A(H_23_), .B(micro_hash_ucr_c_7_), .Y(_2437_) );
XNOR2X1 XNOR2X1_199 ( .A(_2436_), .B(_2437_), .Y(_2438_) );
OAI21X1 OAI21X1_702 ( .A(H_23_), .B(_2399_), .C(_131__bF_buf13), .Y(_2439_) );
AOI21X1 AOI21X1_280 ( .A(micro_hash_ucr_pipe70_bF_buf2), .B(_2438_), .C(_2439_), .Y(_129__23_) );
INVX1 INVX1_305 ( .A(H_8_), .Y(_2440_) );
INVX8 INVX8_70 ( .A(micro_hash_ucr_pipe70_bF_buf3), .Y(_2441_) );
OAI21X1 OAI21X1_703 ( .A(micro_hash_ucr_b_0_bF_buf0_), .B(_2441__bF_buf3), .C(_2399_), .Y(_2442_) );
NOR2X1 NOR2X1_486 ( .A(_330_), .B(_2440_), .Y(_2443_) );
INVX1 INVX1_306 ( .A(_2443_), .Y(_2444_) );
OAI21X1 OAI21X1_704 ( .A(_2444_), .B(_2441__bF_buf1), .C(_131__bF_buf13), .Y(_2445_) );
AOI21X1 AOI21X1_281 ( .A(_2440_), .B(_2442_), .C(_2445_), .Y(_129__8_) );
INVX1 INVX1_307 ( .A(H_9_), .Y(_2446_) );
NOR2X1 NOR2X1_487 ( .A(micro_hash_ucr_b_1_bF_buf1_), .B(H_9_), .Y(_2447_) );
INVX8 INVX8_71 ( .A(micro_hash_ucr_b_1_bF_buf0_), .Y(_2448_) );
NOR2X1 NOR2X1_488 ( .A(_2448_), .B(_2446_), .Y(_2449_) );
NOR2X1 NOR2X1_489 ( .A(_2447_), .B(_2449_), .Y(_2450_) );
AOI21X1 AOI21X1_282 ( .A(_2443_), .B(_2450_), .C(_2441__bF_buf1), .Y(_2451_) );
OAI21X1 OAI21X1_705 ( .A(_2443_), .B(_2450_), .C(_2451_), .Y(_2452_) );
OAI21X1 OAI21X1_706 ( .A(_2446_), .B(_2399_), .C(_2452_), .Y(_2453_) );
AND2X2 AND2X2_87 ( .A(_2453_), .B(_131__bF_buf13), .Y(_129__9_) );
INVX1 INVX1_308 ( .A(H_10_), .Y(_2454_) );
INVX1 INVX1_309 ( .A(_2449_), .Y(_2455_) );
OAI21X1 OAI21X1_707 ( .A(_2444_), .B(_2447_), .C(_2455_), .Y(_2456_) );
XOR2X1 XOR2X1_46 ( .A(micro_hash_ucr_b_2_bF_buf1_), .B(H_10_), .Y(_2457_) );
INVX1 INVX1_310 ( .A(_2456_), .Y(_2458_) );
INVX1 INVX1_311 ( .A(_2457_), .Y(_2459_) );
NOR2X1 NOR2X1_490 ( .A(_2459_), .B(_2458_), .Y(_2460_) );
NOR2X1 NOR2X1_491 ( .A(_2441__bF_buf1), .B(_2460_), .Y(_2461_) );
OAI21X1 OAI21X1_708 ( .A(_2456_), .B(_2457_), .C(_2461_), .Y(_2462_) );
OAI21X1 OAI21X1_709 ( .A(_2454_), .B(_2399_), .C(_2462_), .Y(_2463_) );
AND2X2 AND2X2_88 ( .A(_2463_), .B(_131__bF_buf13), .Y(_129__10_) );
INVX8 INVX8_72 ( .A(micro_hash_ucr_b_2_bF_buf0_), .Y(_2464_) );
INVX1 INVX1_312 ( .A(_2460_), .Y(_2465_) );
OAI21X1 OAI21X1_710 ( .A(_2464_), .B(_2454_), .C(_2465_), .Y(_2466_) );
NOR2X1 NOR2X1_492 ( .A(micro_hash_ucr_b_3_bF_buf1_), .B(H_11_), .Y(_2467_) );
INVX8 INVX8_73 ( .A(micro_hash_ucr_b_3_bF_buf0_), .Y(_2468_) );
INVX1 INVX1_313 ( .A(H_11_), .Y(_2469_) );
NOR2X1 NOR2X1_493 ( .A(_2468_), .B(_2469_), .Y(_2470_) );
OR2X2 OR2X2_25 ( .A(_2470_), .B(_2467_), .Y(_2471_) );
OAI21X1 OAI21X1_711 ( .A(_2466_), .B(_2471_), .C(micro_hash_ucr_pipe70_bF_buf0), .Y(_2472_) );
AOI21X1 AOI21X1_283 ( .A(_2466_), .B(_2471_), .C(_2472_), .Y(_2473_) );
OAI21X1 OAI21X1_712 ( .A(H_11_), .B(_2399_), .C(_131__bF_buf13), .Y(_2474_) );
NOR2X1 NOR2X1_494 ( .A(_2474_), .B(_2473_), .Y(_129__11_) );
XOR2X1 XOR2X1_47 ( .A(micro_hash_ucr_b_4_), .B(H_12_), .Y(_2475_) );
INVX1 INVX1_314 ( .A(_2467_), .Y(_2476_) );
AOI21X1 AOI21X1_284 ( .A(_2476_), .B(_2466_), .C(_2470_), .Y(_2477_) );
XNOR2X1 XNOR2X1_200 ( .A(_2477_), .B(_2475_), .Y(_2478_) );
INVX1 INVX1_315 ( .A(H_12_), .Y(_2479_) );
OAI21X1 OAI21X1_713 ( .A(_2479_), .B(micro_hash_ucr_pipe5), .C(_2441__bF_buf2), .Y(_2480_) );
OAI21X1 OAI21X1_714 ( .A(_2478_), .B(_2441__bF_buf2), .C(_2480_), .Y(_2481_) );
NOR2X1 NOR2X1_495 ( .A(_292__bF_buf2), .B(_2481_), .Y(_129__12_) );
NAND2X1 NAND2X1_338 ( .A(micro_hash_ucr_b_4_), .B(H_12_), .Y(_2482_) );
INVX1 INVX1_316 ( .A(_2475_), .Y(_2483_) );
OAI21X1 OAI21X1_715 ( .A(_2477_), .B(_2483_), .C(_2482_), .Y(_2484_) );
INVX2 INVX2_148 ( .A(_2484_), .Y(_2485_) );
NOR2X1 NOR2X1_496 ( .A(micro_hash_ucr_b_5_bF_buf1_), .B(H_13_), .Y(_2486_) );
INVX8 INVX8_74 ( .A(micro_hash_ucr_b_5_bF_buf0_), .Y(_2487_) );
INVX1 INVX1_317 ( .A(H_13_), .Y(_2488_) );
NOR2X1 NOR2X1_497 ( .A(_2487__bF_buf1), .B(_2488_), .Y(_2489_) );
NOR2X1 NOR2X1_498 ( .A(_2486_), .B(_2489_), .Y(_2490_) );
AND2X2 AND2X2_89 ( .A(_2485_), .B(_2490_), .Y(_2491_) );
OAI21X1 OAI21X1_716 ( .A(_2485_), .B(_2490_), .C(micro_hash_ucr_pipe70_bF_buf0), .Y(_2492_) );
OAI21X1 OAI21X1_717 ( .A(_2488_), .B(micro_hash_ucr_pipe5), .C(_2441__bF_buf2), .Y(_2493_) );
OAI21X1 OAI21X1_718 ( .A(_2491_), .B(_2492_), .C(_2493_), .Y(_2494_) );
NOR2X1 NOR2X1_499 ( .A(_292__bF_buf2), .B(_2494_), .Y(_129__13_) );
XOR2X1 XOR2X1_48 ( .A(micro_hash_ucr_b_6_bF_buf1_), .B(H_14_), .Y(_2495_) );
INVX1 INVX1_318 ( .A(_2489_), .Y(_2496_) );
OAI21X1 OAI21X1_719 ( .A(_2485_), .B(_2486_), .C(_2496_), .Y(_2497_) );
XNOR2X1 XNOR2X1_201 ( .A(_2497_), .B(_2495_), .Y(_2498_) );
INVX1 INVX1_319 ( .A(H_14_), .Y(_2499_) );
OAI21X1 OAI21X1_720 ( .A(_2499_), .B(micro_hash_ucr_pipe5), .C(_2441__bF_buf2), .Y(_2500_) );
NAND2X1 NAND2X1_339 ( .A(_2500_), .B(_131__bF_buf13), .Y(_2501_) );
AOI21X1 AOI21X1_285 ( .A(micro_hash_ucr_pipe70_bF_buf1), .B(_2498_), .C(_2501_), .Y(_129__14_) );
NAND2X1 NAND2X1_340 ( .A(_2495_), .B(_2497_), .Y(_2502_) );
OAI21X1 OAI21X1_721 ( .A(_399__bF_buf3), .B(_2499_), .C(_2502_), .Y(_2503_) );
XOR2X1 XOR2X1_49 ( .A(micro_hash_ucr_b_7_bF_buf3_), .B(H_15_), .Y(_2504_) );
XNOR2X1 XNOR2X1_202 ( .A(_2503_), .B(_2504_), .Y(_2505_) );
OAI21X1 OAI21X1_722 ( .A(H_15_), .B(_2399_), .C(_131__bF_buf6), .Y(_2506_) );
AOI21X1 AOI21X1_286 ( .A(micro_hash_ucr_pipe70_bF_buf1), .B(_2505_), .C(_2506_), .Y(_129__15_) );
INVX1 INVX1_320 ( .A(H_0_), .Y(_2507_) );
OAI21X1 OAI21X1_723 ( .A(micro_hash_ucr_a_0_bF_buf0_), .B(_2441__bF_buf3), .C(_2399_), .Y(_2508_) );
NOR2X1 NOR2X1_500 ( .A(_331_), .B(_2507_), .Y(_2509_) );
INVX1 INVX1_321 ( .A(_2509_), .Y(_2510_) );
OAI21X1 OAI21X1_724 ( .A(_2510_), .B(_2441__bF_buf3), .C(_131__bF_buf13), .Y(_2511_) );
AOI21X1 AOI21X1_287 ( .A(_2507_), .B(_2508_), .C(_2511_), .Y(_129__0_) );
INVX1 INVX1_322 ( .A(H_1_), .Y(_2512_) );
NOR2X1 NOR2X1_501 ( .A(micro_hash_ucr_a_1_), .B(H_1_), .Y(_2513_) );
INVX8 INVX8_75 ( .A(micro_hash_ucr_a_1_), .Y(_2514_) );
NOR2X1 NOR2X1_502 ( .A(_2514__bF_buf2), .B(_2512_), .Y(_2515_) );
NOR2X1 NOR2X1_503 ( .A(_2513_), .B(_2515_), .Y(_2516_) );
AOI21X1 AOI21X1_288 ( .A(_2509_), .B(_2516_), .C(_2441__bF_buf3), .Y(_2517_) );
OAI21X1 OAI21X1_725 ( .A(_2509_), .B(_2516_), .C(_2517_), .Y(_2518_) );
OAI21X1 OAI21X1_726 ( .A(_2512_), .B(_2399_), .C(_2518_), .Y(_2519_) );
AND2X2 AND2X2_90 ( .A(_2519_), .B(_131__bF_buf13), .Y(_129__1_) );
INVX1 INVX1_323 ( .A(_2515_), .Y(_2520_) );
OAI21X1 OAI21X1_727 ( .A(_2510_), .B(_2513_), .C(_2520_), .Y(_2521_) );
XOR2X1 XOR2X1_50 ( .A(micro_hash_ucr_a_2_bF_buf2_), .B(H_2_), .Y(_2522_) );
INVX1 INVX1_324 ( .A(_2521_), .Y(_2523_) );
INVX1 INVX1_325 ( .A(_2522_), .Y(_2524_) );
NOR2X1 NOR2X1_504 ( .A(_2524_), .B(_2523_), .Y(_2525_) );
NOR2X1 NOR2X1_505 ( .A(_2441__bF_buf3), .B(_2525_), .Y(_2526_) );
OAI21X1 OAI21X1_728 ( .A(_2521_), .B(_2522_), .C(_2526_), .Y(_2527_) );
NAND2X1 NAND2X1_341 ( .A(H_2_), .B(_2389_), .Y(_2528_) );
AOI21X1 AOI21X1_289 ( .A(_2528_), .B(_2527_), .C(_292__bF_buf2), .Y(_129__2_) );
AOI21X1 AOI21X1_290 ( .A(micro_hash_ucr_a_2_bF_buf1_), .B(H_2_), .C(_2525_), .Y(_2529_) );
NOR2X1 NOR2X1_506 ( .A(micro_hash_ucr_a_3_bF_buf1_), .B(H_3_), .Y(_2530_) );
INVX8 INVX8_76 ( .A(micro_hash_ucr_a_3_bF_buf0_), .Y(_2531_) );
INVX2 INVX2_149 ( .A(H_3_), .Y(_2532_) );
NOR2X1 NOR2X1_507 ( .A(_2531_), .B(_2532_), .Y(_2533_) );
NOR2X1 NOR2X1_508 ( .A(_2530_), .B(_2533_), .Y(_2534_) );
AND2X2 AND2X2_91 ( .A(_2529_), .B(_2534_), .Y(_2535_) );
OAI21X1 OAI21X1_729 ( .A(_2529_), .B(_2534_), .C(micro_hash_ucr_pipe70_bF_buf3), .Y(_2536_) );
OAI21X1 OAI21X1_730 ( .A(_2532_), .B(micro_hash_ucr_pipe5), .C(_2441__bF_buf1), .Y(_2537_) );
OAI21X1 OAI21X1_731 ( .A(_2535_), .B(_2536_), .C(_2537_), .Y(_2538_) );
NOR2X1 NOR2X1_509 ( .A(_292__bF_buf2), .B(_2538_), .Y(_129__3_) );
XOR2X1 XOR2X1_51 ( .A(micro_hash_ucr_a_4_bF_buf1_), .B(H_4_), .Y(_2539_) );
INVX1 INVX1_326 ( .A(_2533_), .Y(_2540_) );
OAI21X1 OAI21X1_732 ( .A(_2529_), .B(_2530_), .C(_2540_), .Y(_2541_) );
XNOR2X1 XNOR2X1_203 ( .A(_2541_), .B(_2539_), .Y(_2542_) );
INVX2 INVX2_150 ( .A(H_4_), .Y(_2543_) );
OAI21X1 OAI21X1_733 ( .A(_2543_), .B(micro_hash_ucr_pipe5), .C(_2441__bF_buf1), .Y(_2544_) );
NAND2X1 NAND2X1_342 ( .A(_2544_), .B(_131__bF_buf13), .Y(_2545_) );
AOI21X1 AOI21X1_291 ( .A(micro_hash_ucr_pipe70_bF_buf3), .B(_2542_), .C(_2545_), .Y(_129__4_) );
INVX8 INVX8_77 ( .A(micro_hash_ucr_a_4_bF_buf0_), .Y(_2546_) );
NAND2X1 NAND2X1_343 ( .A(_2539_), .B(_2541_), .Y(_2547_) );
OAI21X1 OAI21X1_734 ( .A(_2546_), .B(_2543_), .C(_2547_), .Y(_2548_) );
INVX2 INVX2_151 ( .A(_2548_), .Y(_2549_) );
NOR2X1 NOR2X1_510 ( .A(micro_hash_ucr_a_5_bF_buf1_), .B(H_5_), .Y(_2550_) );
INVX8 INVX8_78 ( .A(micro_hash_ucr_a_5_bF_buf0_), .Y(_2551_) );
INVX1 INVX1_327 ( .A(H_5_), .Y(_2552_) );
NOR2X1 NOR2X1_511 ( .A(_2551_), .B(_2552_), .Y(_2553_) );
NOR2X1 NOR2X1_512 ( .A(_2550_), .B(_2553_), .Y(_2554_) );
AND2X2 AND2X2_92 ( .A(_2549_), .B(_2554_), .Y(_2555_) );
OAI21X1 OAI21X1_735 ( .A(_2549_), .B(_2554_), .C(micro_hash_ucr_pipe70_bF_buf0), .Y(_2556_) );
OAI21X1 OAI21X1_736 ( .A(_2552_), .B(micro_hash_ucr_pipe5), .C(_2441__bF_buf0), .Y(_2557_) );
OAI21X1 OAI21X1_737 ( .A(_2555_), .B(_2556_), .C(_2557_), .Y(_2558_) );
NOR2X1 NOR2X1_513 ( .A(_292__bF_buf2), .B(_2558_), .Y(_129__5_) );
XOR2X1 XOR2X1_52 ( .A(micro_hash_ucr_a_6_bF_buf1_), .B(H_6_), .Y(_2559_) );
INVX1 INVX1_328 ( .A(_2553_), .Y(_2560_) );
OAI21X1 OAI21X1_738 ( .A(_2549_), .B(_2550_), .C(_2560_), .Y(_2561_) );
XOR2X1 XOR2X1_53 ( .A(_2561_), .B(_2559_), .Y(_2562_) );
INVX1 INVX1_329 ( .A(H_6_), .Y(_2563_) );
OAI21X1 OAI21X1_739 ( .A(_2563_), .B(micro_hash_ucr_pipe5), .C(_2441__bF_buf0), .Y(_2564_) );
OAI21X1 OAI21X1_740 ( .A(_2562_), .B(_2441__bF_buf0), .C(_2564_), .Y(_2565_) );
NOR2X1 NOR2X1_514 ( .A(_292__bF_buf2), .B(_2565_), .Y(_129__6_) );
NAND2X1 NAND2X1_344 ( .A(_2559_), .B(_2561_), .Y(_2566_) );
OAI21X1 OAI21X1_741 ( .A(_400_), .B(_2563_), .C(_2566_), .Y(_2567_) );
XNOR2X1 XNOR2X1_204 ( .A(micro_hash_ucr_a_7_bF_buf1_), .B(H_7_), .Y(_2568_) );
AND2X2 AND2X2_93 ( .A(_2567_), .B(_2568_), .Y(_2569_) );
OAI21X1 OAI21X1_742 ( .A(_2567_), .B(_2568_), .C(micro_hash_ucr_pipe70_bF_buf0), .Y(_2570_) );
INVX1 INVX1_330 ( .A(H_7_), .Y(_2571_) );
OAI21X1 OAI21X1_743 ( .A(_2571_), .B(micro_hash_ucr_pipe5), .C(_2441__bF_buf0), .Y(_2572_) );
OAI21X1 OAI21X1_744 ( .A(_2569_), .B(_2570_), .C(_2572_), .Y(_2573_) );
NOR2X1 NOR2X1_515 ( .A(_292__bF_buf2), .B(_2573_), .Y(_129__7_) );
OAI21X1 OAI21X1_745 ( .A(_507_), .B(micro_hash_ucr_Wx_152_), .C(_421_), .Y(_2574_) );
AOI21X1 AOI21X1_292 ( .A(_507_), .B(micro_hash_ucr_Wx_152_), .C(_2574_), .Y(_2575_) );
NOR2X1 NOR2X1_516 ( .A(_2575_), .B(_292__bF_buf1), .Y(_125__224_) );
OAI21X1 OAI21X1_746 ( .A(_961_), .B(micro_hash_ucr_Wx_153_), .C(_762_), .Y(_2576_) );
AOI21X1 AOI21X1_293 ( .A(_961_), .B(micro_hash_ucr_Wx_153_), .C(_2576_), .Y(_2577_) );
NOR2X1 NOR2X1_517 ( .A(_2577_), .B(_292__bF_buf8), .Y(_125__225_) );
OAI21X1 OAI21X1_747 ( .A(_963_), .B(micro_hash_ucr_Wx_154_), .C(_1064_), .Y(_2578_) );
AOI21X1 AOI21X1_294 ( .A(_963_), .B(micro_hash_ucr_Wx_154_), .C(_2578_), .Y(_2579_) );
NOR2X1 NOR2X1_518 ( .A(_2579_), .B(_292__bF_buf3), .Y(_125__226_) );
OAI21X1 OAI21X1_748 ( .A(_1298_), .B(micro_hash_ucr_Wx_155_), .C(_1381_), .Y(_2580_) );
AOI21X1 AOI21X1_295 ( .A(_1298_), .B(micro_hash_ucr_Wx_155_), .C(_2580_), .Y(_2581_) );
NOR2X1 NOR2X1_519 ( .A(_2581_), .B(_292__bF_buf12), .Y(_125__227_) );
AOI21X1 AOI21X1_296 ( .A(micro_hash_ucr_Wx_156_), .B(_1828_), .C(micro_hash_ucr_Wx_204_), .Y(_2582_) );
OAI21X1 OAI21X1_749 ( .A(_1828_), .B(micro_hash_ucr_Wx_156_), .C(_2582_), .Y(_2583_) );
AND2X2 AND2X2_94 ( .A(_2583_), .B(_131__bF_buf12), .Y(_125__228_) );
AOI21X1 AOI21X1_297 ( .A(micro_hash_ucr_Wx_157_), .B(_2054_), .C(micro_hash_ucr_Wx_205_), .Y(_2584_) );
OAI21X1 OAI21X1_750 ( .A(_2054_), .B(micro_hash_ucr_Wx_157_), .C(_2584_), .Y(_2585_) );
AND2X2 AND2X2_95 ( .A(_2585_), .B(_131__bF_buf10), .Y(_125__229_) );
OAI21X1 OAI21X1_751 ( .A(_2094_), .B(micro_hash_ucr_Wx_118_), .C(_2137_), .Y(_2586_) );
AOI21X1 AOI21X1_298 ( .A(_2094_), .B(micro_hash_ucr_Wx_118_), .C(_2586_), .Y(_2587_) );
NOR2X1 NOR2X1_520 ( .A(_2587_), .B(_292__bF_buf9), .Y(_125__230_) );
INVX2 INVX2_152 ( .A(micro_hash_ucr_Wx_159_), .Y(_2588_) );
AOI21X1 AOI21X1_299 ( .A(micro_hash_ucr_Wx_119_), .B(_2588_), .C(micro_hash_ucr_Wx_207_), .Y(_2589_) );
OAI21X1 OAI21X1_752 ( .A(_2588_), .B(micro_hash_ucr_Wx_119_), .C(_2589_), .Y(_2590_) );
AND2X2 AND2X2_96 ( .A(_2590_), .B(_131__bF_buf0), .Y(_125__231_) );
AOI21X1 AOI21X1_300 ( .A(micro_hash_ucr_Wx_168_), .B(_516_), .C(micro_hash_ucr_Wx_216_), .Y(_2591_) );
OAI21X1 OAI21X1_753 ( .A(_516_), .B(micro_hash_ucr_Wx_168_), .C(_2591_), .Y(_2592_) );
AND2X2 AND2X2_97 ( .A(_2592_), .B(_131__bF_buf3), .Y(_125__240_) );
OAI21X1 OAI21X1_754 ( .A(_709_), .B(micro_hash_ucr_Wx_169_), .C(_780_), .Y(_2593_) );
AOI21X1 AOI21X1_301 ( .A(_709_), .B(micro_hash_ucr_Wx_169_), .C(_2593_), .Y(_2594_) );
NOR2X1 NOR2X1_521 ( .A(_2594_), .B(_292__bF_buf8), .Y(_125__241_) );
OAI21X1 OAI21X1_755 ( .A(_983_), .B(micro_hash_ucr_Wx_170_), .C(_1071_), .Y(_2595_) );
AOI21X1 AOI21X1_302 ( .A(_983_), .B(micro_hash_ucr_Wx_170_), .C(_2595_), .Y(_2596_) );
NOR2X1 NOR2X1_522 ( .A(_2596_), .B(_292__bF_buf3), .Y(_125__242_) );
OAI21X1 OAI21X1_756 ( .A(_1309_), .B(micro_hash_ucr_Wx_171_), .C(_1133_), .Y(_2597_) );
AOI21X1 AOI21X1_303 ( .A(_1309_), .B(micro_hash_ucr_Wx_171_), .C(_2597_), .Y(_2598_) );
NOR2X1 NOR2X1_523 ( .A(_2598_), .B(_292__bF_buf0), .Y(_125__243_) );
AOI21X1 AOI21X1_304 ( .A(micro_hash_ucr_Wx_172_), .B(_1555_), .C(micro_hash_ucr_Wx_220_), .Y(_2599_) );
OAI21X1 OAI21X1_757 ( .A(_1555_), .B(micro_hash_ucr_Wx_172_), .C(_2599_), .Y(_2600_) );
AND2X2 AND2X2_98 ( .A(_2600_), .B(_131__bF_buf10), .Y(_125__244_) );
AOI21X1 AOI21X1_305 ( .A(micro_hash_ucr_Wx_173_), .B(_1838_), .C(micro_hash_ucr_Wx_221_), .Y(_2601_) );
OAI21X1 OAI21X1_758 ( .A(_1838_), .B(micro_hash_ucr_Wx_173_), .C(_2601_), .Y(_2602_) );
AND2X2 AND2X2_99 ( .A(_2602_), .B(_131__bF_buf10), .Y(_125__245_) );
OAI21X1 OAI21X1_759 ( .A(_2110_), .B(micro_hash_ucr_Wx_134_), .C(_2150_), .Y(_2603_) );
AOI21X1 AOI21X1_306 ( .A(_2110_), .B(micro_hash_ucr_Wx_134_), .C(_2603_), .Y(_2604_) );
NOR2X1 NOR2X1_524 ( .A(_2604_), .B(_292__bF_buf9), .Y(_125__246_) );
AOI21X1 AOI21X1_307 ( .A(micro_hash_ucr_Wx_175_), .B(_2295_), .C(micro_hash_ucr_Wx_223_), .Y(_2605_) );
OAI21X1 OAI21X1_760 ( .A(micro_hash_ucr_Wx_175_), .B(_2295_), .C(_2605_), .Y(_2606_) );
AND2X2 AND2X2_100 ( .A(_2606_), .B(_131__bF_buf0), .Y(_125__247_) );
AOI21X1 AOI21X1_308 ( .A(micro_hash_ucr_Wx_160_), .B(_512_), .C(micro_hash_ucr_Wx_208_), .Y(_2607_) );
OAI21X1 OAI21X1_761 ( .A(_512_), .B(micro_hash_ucr_Wx_160_), .C(_2607_), .Y(_2608_) );
AND2X2 AND2X2_101 ( .A(_2608_), .B(_131__bF_buf3), .Y(_125__232_) );
AOI21X1 AOI21X1_309 ( .A(micro_hash_ucr_Wx_161_), .B(_702_), .C(micro_hash_ucr_Wx_209_), .Y(_2609_) );
OAI21X1 OAI21X1_762 ( .A(_702_), .B(micro_hash_ucr_Wx_161_), .C(_2609_), .Y(_2610_) );
AND2X2 AND2X2_102 ( .A(_2610_), .B(_131__bF_buf8), .Y(_125__233_) );
OAI21X1 OAI21X1_763 ( .A(_971_), .B(micro_hash_ucr_Wx_162_), .C(_815_), .Y(_2611_) );
AOI21X1 AOI21X1_310 ( .A(_971_), .B(micro_hash_ucr_Wx_162_), .C(_2611_), .Y(_2612_) );
NOR2X1 NOR2X1_525 ( .A(_2612_), .B(_292__bF_buf3), .Y(_125__234_) );
OAI21X1 OAI21X1_764 ( .A(_1154_), .B(micro_hash_ucr_Wx_163_), .C(_1390_), .Y(_2613_) );
AOI21X1 AOI21X1_311 ( .A(_1154_), .B(micro_hash_ucr_Wx_163_), .C(_2613_), .Y(_2614_) );
NOR2X1 NOR2X1_526 ( .A(_2614_), .B(_292__bF_buf0), .Y(_125__235_) );
AOI21X1 AOI21X1_312 ( .A(micro_hash_ucr_Wx_164_), .B(_1703_), .C(micro_hash_ucr_Wx_212_), .Y(_2615_) );
OAI21X1 OAI21X1_765 ( .A(_1703_), .B(micro_hash_ucr_Wx_164_), .C(_2615_), .Y(_2616_) );
AND2X2 AND2X2_103 ( .A(_2616_), .B(_131__bF_buf10), .Y(_125__236_) );
AOI21X1 AOI21X1_313 ( .A(micro_hash_ucr_Wx_165_), .B(_1705_), .C(micro_hash_ucr_Wx_213_), .Y(_2617_) );
OAI21X1 OAI21X1_766 ( .A(_1705_), .B(micro_hash_ucr_Wx_165_), .C(_2617_), .Y(_2618_) );
AND2X2 AND2X2_104 ( .A(_2618_), .B(_131__bF_buf10), .Y(_125__237_) );
OAI21X1 OAI21X1_767 ( .A(_2102_), .B(micro_hash_ucr_Wx_126_), .C(_2142_), .Y(_2619_) );
AOI21X1 AOI21X1_314 ( .A(_2102_), .B(micro_hash_ucr_Wx_126_), .C(_2619_), .Y(_2620_) );
NOR2X1 NOR2X1_527 ( .A(_2620_), .B(_292__bF_buf6), .Y(_125__238_) );
INVX2 INVX2_153 ( .A(micro_hash_ucr_Wx_127_), .Y(_2621_) );
AOI21X1 AOI21X1_315 ( .A(micro_hash_ucr_Wx_167_), .B(_2621_), .C(micro_hash_ucr_Wx_215_), .Y(_2622_) );
OAI21X1 OAI21X1_768 ( .A(micro_hash_ucr_Wx_167_), .B(_2621_), .C(_2622_), .Y(_2623_) );
AND2X2 AND2X2_105 ( .A(_2623_), .B(_131__bF_buf0), .Y(_125__239_) );
AOI21X1 AOI21X1_316 ( .A(micro_hash_ucr_Wx_128_), .B(_493_), .C(micro_hash_ucr_Wx_176_), .Y(_2624_) );
OAI21X1 OAI21X1_769 ( .A(_493_), .B(micro_hash_ucr_Wx_128_), .C(_2624_), .Y(_2625_) );
AND2X2 AND2X2_106 ( .A(_2625_), .B(_131__bF_buf3), .Y(_125__200_) );
OAI21X1 OAI21X1_770 ( .A(_671_), .B(micro_hash_ucr_Wx_129_), .C(_743_), .Y(_2626_) );
AOI21X1 AOI21X1_317 ( .A(_671_), .B(micro_hash_ucr_Wx_129_), .C(_2626_), .Y(_2627_) );
NOR2X1 NOR2X1_528 ( .A(_2627_), .B(_292__bF_buf0), .Y(_125__201_) );
OAI21X1 OAI21X1_771 ( .A(_939_), .B(micro_hash_ucr_Wx_130_), .C(_1037_), .Y(_2628_) );
AOI21X1 AOI21X1_318 ( .A(_939_), .B(micro_hash_ucr_Wx_130_), .C(_2628_), .Y(_2629_) );
NOR2X1 NOR2X1_529 ( .A(_2629_), .B(_292__bF_buf3), .Y(_125__202_) );
OAI21X1 OAI21X1_772 ( .A(_1163_), .B(micro_hash_ucr_Wx_131_), .C(_1360_), .Y(_2630_) );
AOI21X1 AOI21X1_319 ( .A(_1163_), .B(micro_hash_ucr_Wx_131_), .C(_2630_), .Y(_2631_) );
NOR2X1 NOR2X1_530 ( .A(_2631_), .B(_292__bF_buf12), .Y(_125__203_) );
AOI21X1 AOI21X1_320 ( .A(micro_hash_ucr_Wx_92_), .B(_1555_), .C(micro_hash_ucr_Wx_180_), .Y(_2632_) );
OAI21X1 OAI21X1_773 ( .A(micro_hash_ucr_Wx_92_), .B(_1555_), .C(_2632_), .Y(_2633_) );
AND2X2 AND2X2_107 ( .A(_2633_), .B(_131__bF_buf10), .Y(_125__204_) );
OAI21X1 OAI21X1_774 ( .A(_1712_), .B(micro_hash_ucr_Wx_133_), .C(_1874_), .Y(_2634_) );
AOI21X1 AOI21X1_321 ( .A(_1712_), .B(micro_hash_ucr_Wx_133_), .C(_2634_), .Y(_2635_) );
NOR2X1 NOR2X1_531 ( .A(_2635_), .B(_292__bF_buf11), .Y(_125__205_) );
OAI21X1 OAI21X1_775 ( .A(_2069_), .B(micro_hash_ucr_Wx_94_), .C(_2116_), .Y(_2636_) );
AOI21X1 AOI21X1_322 ( .A(micro_hash_ucr_Wx_94_), .B(_2069_), .C(_2636_), .Y(_2637_) );
NOR2X1 NOR2X1_532 ( .A(_2637_), .B(_292__bF_buf9), .Y(_125__206_) );
OAI21X1 OAI21X1_776 ( .A(_2271_), .B(micro_hash_ucr_Wx_135_), .C(_2324_), .Y(_2638_) );
AOI21X1 AOI21X1_323 ( .A(_2271_), .B(micro_hash_ucr_Wx_135_), .C(_2638_), .Y(_2639_) );
NOR2X1 NOR2X1_533 ( .A(_2639_), .B(_292__bF_buf9), .Y(_125__207_) );
AOI21X1 AOI21X1_324 ( .A(micro_hash_ucr_Wx_144_), .B(_503_), .C(micro_hash_ucr_Wx_192_), .Y(_2640_) );
OAI21X1 OAI21X1_777 ( .A(_503_), .B(micro_hash_ucr_Wx_144_), .C(_2640_), .Y(_2641_) );
AND2X2 AND2X2_108 ( .A(_2641_), .B(_131__bF_buf3), .Y(_125__216_) );
OAI21X1 OAI21X1_778 ( .A(_685_), .B(micro_hash_ucr_Wx_145_), .C(_755_), .Y(_2642_) );
AOI21X1 AOI21X1_325 ( .A(_685_), .B(micro_hash_ucr_Wx_145_), .C(_2642_), .Y(_2643_) );
NOR2X1 NOR2X1_534 ( .A(_2643_), .B(_292__bF_buf3), .Y(_125__217_) );
OAI21X1 OAI21X1_779 ( .A(_953_), .B(micro_hash_ucr_Wx_146_), .C(_1054_), .Y(_2644_) );
AOI21X1 AOI21X1_326 ( .A(_953_), .B(micro_hash_ucr_Wx_146_), .C(_2644_), .Y(_2645_) );
NOR2X1 NOR2X1_535 ( .A(_2645_), .B(_292__bF_buf3), .Y(_125__218_) );
OAI21X1 OAI21X1_780 ( .A(_1289_), .B(micro_hash_ucr_Wx_147_), .C(_1371_), .Y(_2646_) );
AOI21X1 AOI21X1_327 ( .A(_1289_), .B(micro_hash_ucr_Wx_147_), .C(_2646_), .Y(_2647_) );
NOR2X1 NOR2X1_536 ( .A(_2647_), .B(_292__bF_buf12), .Y(_125__219_) );
AOI21X1 AOI21X1_328 ( .A(micro_hash_ucr_Wx_148_), .B(_1532_), .C(micro_hash_ucr_Wx_196_), .Y(_2648_) );
OAI21X1 OAI21X1_781 ( .A(_1532_), .B(micro_hash_ucr_Wx_148_), .C(_2648_), .Y(_2649_) );
AND2X2 AND2X2_109 ( .A(_2649_), .B(_131__bF_buf12), .Y(_125__220_) );
OAI21X1 OAI21X1_782 ( .A(_2045_), .B(micro_hash_ucr_Wx_149_), .C(_1885_), .Y(_2650_) );
AOI21X1 AOI21X1_329 ( .A(_2045_), .B(micro_hash_ucr_Wx_149_), .C(_2650_), .Y(_2651_) );
NOR2X1 NOR2X1_537 ( .A(_2651_), .B(_292__bF_buf6), .Y(_125__221_) );
OAI21X1 OAI21X1_783 ( .A(_2085_), .B(micro_hash_ucr_Wx_110_), .C(_2335_), .Y(_2652_) );
AOI21X1 AOI21X1_330 ( .A(_2085_), .B(micro_hash_ucr_Wx_110_), .C(_2652_), .Y(_2653_) );
NOR2X1 NOR2X1_538 ( .A(_2653_), .B(_292__bF_buf6), .Y(_125__222_) );
AOI21X1 AOI21X1_331 ( .A(micro_hash_ucr_Wx_151_), .B(_2282_), .C(micro_hash_ucr_Wx_199_), .Y(_2654_) );
OAI21X1 OAI21X1_784 ( .A(micro_hash_ucr_Wx_151_), .B(_2282_), .C(_2654_), .Y(_2655_) );
AND2X2 AND2X2_110 ( .A(_2655_), .B(_131__bF_buf0), .Y(_125__223_) );
AOI21X1 AOI21X1_332 ( .A(micro_hash_ucr_Wx_136_), .B(_498_), .C(micro_hash_ucr_Wx_184_), .Y(_2656_) );
OAI21X1 OAI21X1_785 ( .A(_498_), .B(micro_hash_ucr_Wx_136_), .C(_2656_), .Y(_2657_) );
AND2X2 AND2X2_111 ( .A(_2657_), .B(_131__bF_buf3), .Y(_125__208_) );
OAI21X1 OAI21X1_786 ( .A(_944_), .B(micro_hash_ucr_Wx_137_), .C(_749_), .Y(_2658_) );
AOI21X1 AOI21X1_333 ( .A(_944_), .B(micro_hash_ucr_Wx_137_), .C(_2658_), .Y(_2659_) );
NOR2X1 NOR2X1_539 ( .A(_2659_), .B(_292__bF_buf8), .Y(_125__209_) );
OAI21X1 OAI21X1_787 ( .A(_946_), .B(micro_hash_ucr_Wx_138_), .C(_1045_), .Y(_2660_) );
AOI21X1 AOI21X1_334 ( .A(_946_), .B(micro_hash_ucr_Wx_138_), .C(_2660_), .Y(_2661_) );
NOR2X1 NOR2X1_540 ( .A(_2661_), .B(_292__bF_buf3), .Y(_125__210_) );
OAI21X1 OAI21X1_788 ( .A(_1280_), .B(micro_hash_ucr_Wx_139_), .C(_1140_), .Y(_2662_) );
AOI21X1 AOI21X1_335 ( .A(_1280_), .B(micro_hash_ucr_Wx_139_), .C(_2662_), .Y(_2663_) );
NOR2X1 NOR2X1_541 ( .A(_2663_), .B(_292__bF_buf12), .Y(_125__211_) );
AOI21X1 AOI21X1_336 ( .A(micro_hash_ucr_Wx_140_), .B(_1525_), .C(micro_hash_ucr_Wx_188_), .Y(_2664_) );
OAI21X1 OAI21X1_789 ( .A(_1525_), .B(micro_hash_ucr_Wx_140_), .C(_2664_), .Y(_2665_) );
AND2X2 AND2X2_112 ( .A(_2665_), .B(_131__bF_buf12), .Y(_125__212_) );
OAI21X1 OAI21X1_790 ( .A(_1816_), .B(micro_hash_ucr_Wx_141_), .C(_1691_), .Y(_2666_) );
AOI21X1 AOI21X1_337 ( .A(_1816_), .B(micro_hash_ucr_Wx_141_), .C(_2666_), .Y(_2667_) );
NOR2X1 NOR2X1_542 ( .A(_2667_), .B(_292__bF_buf6), .Y(_125__213_) );
AOI21X1 AOI21X1_338 ( .A(micro_hash_ucr_Wx_142_), .B(_2036_), .C(micro_hash_ucr_Wx_190_), .Y(_2668_) );
OAI21X1 OAI21X1_791 ( .A(_2036_), .B(micro_hash_ucr_Wx_142_), .C(_2668_), .Y(_2669_) );
AND2X2 AND2X2_113 ( .A(_2669_), .B(_131__bF_buf10), .Y(_125__214_) );
AOI21X1 AOI21X1_339 ( .A(micro_hash_ucr_Wx_143_), .B(_2277_), .C(micro_hash_ucr_Wx_191_), .Y(_2670_) );
OAI21X1 OAI21X1_792 ( .A(_2277_), .B(micro_hash_ucr_Wx_143_), .C(_2670_), .Y(_2671_) );
AND2X2 AND2X2_114 ( .A(_2671_), .B(_131__bF_buf0), .Y(_125__215_) );
AOI21X1 AOI21X1_340 ( .A(micro_hash_ucr_Wx_104_), .B(_476_), .C(micro_hash_ucr_Wx_152_), .Y(_2672_) );
OAI21X1 OAI21X1_793 ( .A(_476_), .B(micro_hash_ucr_Wx_104_), .C(_2672_), .Y(_2673_) );
AND2X2 AND2X2_115 ( .A(_2673_), .B(_131__bF_buf3), .Y(_125__176_) );
OAI21X1 OAI21X1_794 ( .A(_651_), .B(micro_hash_ucr_Wx_105_), .C(_729_), .Y(_2674_) );
AOI21X1 AOI21X1_341 ( .A(_651_), .B(micro_hash_ucr_Wx_105_), .C(_2674_), .Y(_2675_) );
NOR2X1 NOR2X1_543 ( .A(_2675_), .B(_292__bF_buf0), .Y(_125__177_) );
OAI21X1 OAI21X1_795 ( .A(_911_), .B(micro_hash_ucr_Wx_106_), .C(_1011_), .Y(_2676_) );
AOI21X1 AOI21X1_342 ( .A(_911_), .B(micro_hash_ucr_Wx_106_), .C(_2676_), .Y(_2677_) );
NOR2X1 NOR2X1_544 ( .A(_2677_), .B(_292__bF_buf3), .Y(_125__178_) );
OAI21X1 OAI21X1_796 ( .A(_1249_), .B(micro_hash_ucr_Wx_107_), .C(_1147_), .Y(_2678_) );
AOI21X1 AOI21X1_343 ( .A(_1249_), .B(micro_hash_ucr_Wx_107_), .C(_2678_), .Y(_2679_) );
NOR2X1 NOR2X1_545 ( .A(_2679_), .B(_292__bF_buf12), .Y(_125__179_) );
AOI21X1 AOI21X1_344 ( .A(micro_hash_ucr_Wx_68_), .B(_1532_), .C(micro_hash_ucr_Wx_156_), .Y(_2680_) );
OAI21X1 OAI21X1_797 ( .A(micro_hash_ucr_Wx_68_), .B(_1532_), .C(_2680_), .Y(_2681_) );
AND2X2 AND2X2_116 ( .A(_2681_), .B(_131__bF_buf12), .Y(_125__180_) );
OAI21X1 OAI21X1_798 ( .A(_1789_), .B(micro_hash_ucr_Wx_109_), .C(_1698_), .Y(_2682_) );
AOI21X1 AOI21X1_345 ( .A(_1789_), .B(micro_hash_ucr_Wx_109_), .C(_2682_), .Y(_2683_) );
NOR2X1 NOR2X1_546 ( .A(_2683_), .B(_292__bF_buf11), .Y(_125__181_) );
OAI21X1 OAI21X1_799 ( .A(_2003_), .B(micro_hash_ucr_Wx_110_), .C(_2094_), .Y(_2684_) );
AOI21X1 AOI21X1_346 ( .A(_2003_), .B(micro_hash_ucr_Wx_110_), .C(_2684_), .Y(_2685_) );
NOR2X1 NOR2X1_547 ( .A(_2685_), .B(_292__bF_buf9), .Y(_125__182_) );
OAI21X1 OAI21X1_800 ( .A(_2282_), .B(micro_hash_ucr_Wx_71_), .C(_2588_), .Y(_2686_) );
AOI21X1 AOI21X1_347 ( .A(micro_hash_ucr_Wx_71_), .B(_2282_), .C(_2686_), .Y(_2687_) );
NOR2X1 NOR2X1_548 ( .A(_2687_), .B(_292__bF_buf9), .Y(_125__183_) );
AOI21X1 AOI21X1_348 ( .A(micro_hash_ucr_Wx_120_), .B(_488_), .C(micro_hash_ucr_Wx_168_), .Y(_2688_) );
OAI21X1 OAI21X1_801 ( .A(_488_), .B(micro_hash_ucr_Wx_120_), .C(_2688_), .Y(_2689_) );
AND2X2 AND2X2_117 ( .A(_2689_), .B(_131__bF_buf3), .Y(_125__192_) );
OAI21X1 OAI21X1_802 ( .A(_664_), .B(micro_hash_ucr_Wx_121_), .C(_735_), .Y(_2690_) );
AOI21X1 AOI21X1_349 ( .A(_664_), .B(micro_hash_ucr_Wx_121_), .C(_2690_), .Y(_2691_) );
NOR2X1 NOR2X1_549 ( .A(_2691_), .B(_292__bF_buf3), .Y(_125__193_) );
OAI21X1 OAI21X1_803 ( .A(_931_), .B(micro_hash_ucr_Wx_122_), .C(_1028_), .Y(_2692_) );
AOI21X1 AOI21X1_350 ( .A(_931_), .B(micro_hash_ucr_Wx_122_), .C(_2692_), .Y(_2693_) );
NOR2X1 NOR2X1_550 ( .A(_2693_), .B(_292__bF_buf3), .Y(_125__194_) );
OAI21X1 OAI21X1_804 ( .A(_1269_), .B(micro_hash_ucr_Wx_123_), .C(_1349_), .Y(_2694_) );
AOI21X1 AOI21X1_351 ( .A(_1269_), .B(micro_hash_ucr_Wx_123_), .C(_2694_), .Y(_2695_) );
NOR2X1 NOR2X1_551 ( .A(_2695_), .B(_292__bF_buf12), .Y(_125__195_) );
AOI21X1 AOI21X1_352 ( .A(micro_hash_ucr_Wx_124_), .B(_1806_), .C(micro_hash_ucr_Wx_172_), .Y(_2696_) );
OAI21X1 OAI21X1_805 ( .A(_1806_), .B(micro_hash_ucr_Wx_124_), .C(_2696_), .Y(_2697_) );
AND2X2 AND2X2_118 ( .A(_2697_), .B(_131__bF_buf12), .Y(_125__196_) );
OAI21X1 OAI21X1_806 ( .A(_2021_), .B(micro_hash_ucr_Wx_125_), .C(_1865_), .Y(_2698_) );
AOI21X1 AOI21X1_353 ( .A(_2021_), .B(micro_hash_ucr_Wx_125_), .C(_2698_), .Y(_2699_) );
NOR2X1 NOR2X1_552 ( .A(_2699_), .B(_292__bF_buf11), .Y(_125__197_) );
OAI21X1 OAI21X1_807 ( .A(_2019_), .B(micro_hash_ucr_Wx_126_), .C(_2110_), .Y(_2700_) );
AOI21X1 AOI21X1_354 ( .A(_2019_), .B(micro_hash_ucr_Wx_126_), .C(_2700_), .Y(_2701_) );
NOR2X1 NOR2X1_553 ( .A(_2701_), .B(_292__bF_buf6), .Y(_125__198_) );
AOI21X1 AOI21X1_355 ( .A(micro_hash_ucr_Wx_127_), .B(_2266_), .C(micro_hash_ucr_Wx_175_), .Y(_2702_) );
OAI21X1 OAI21X1_808 ( .A(_2266_), .B(micro_hash_ucr_Wx_127_), .C(_2702_), .Y(_2703_) );
AND2X2 AND2X2_119 ( .A(_2703_), .B(_131__bF_buf0), .Y(_125__199_) );
AOI21X1 AOI21X1_356 ( .A(micro_hash_ucr_Wx_112_), .B(_483_), .C(micro_hash_ucr_Wx_160_), .Y(_2704_) );
OAI21X1 OAI21X1_809 ( .A(_483_), .B(micro_hash_ucr_Wx_112_), .C(_2704_), .Y(_2705_) );
AND2X2 AND2X2_120 ( .A(_2705_), .B(_131__bF_buf3), .Y(_125__184_) );
AOI21X1 AOI21X1_357 ( .A(micro_hash_ucr_Wx_113_), .B(_919_), .C(micro_hash_ucr_Wx_161_), .Y(_2706_) );
OAI21X1 OAI21X1_810 ( .A(_919_), .B(micro_hash_ucr_Wx_113_), .C(_2706_), .Y(_2707_) );
AND2X2 AND2X2_121 ( .A(_2707_), .B(_131__bF_buf8), .Y(_125__185_) );
OAI21X1 OAI21X1_811 ( .A(_921_), .B(micro_hash_ucr_Wx_114_), .C(_1020_), .Y(_2708_) );
AOI21X1 AOI21X1_358 ( .A(_921_), .B(micro_hash_ucr_Wx_114_), .C(_2708_), .Y(_2709_) );
NOR2X1 NOR2X1_554 ( .A(_2709_), .B(_292__bF_buf0), .Y(_125__186_) );
OAI21X1 OAI21X1_812 ( .A(_1259_), .B(micro_hash_ucr_Wx_115_), .C(_1339_), .Y(_2710_) );
AOI21X1 AOI21X1_359 ( .A(_1259_), .B(micro_hash_ucr_Wx_115_), .C(_2710_), .Y(_2711_) );
NOR2X1 NOR2X1_555 ( .A(_2711_), .B(_292__bF_buf12), .Y(_125__187_) );
OAI21X1 OAI21X1_813 ( .A(_1796_), .B(micro_hash_ucr_Wx_116_), .C(_1858_), .Y(_2712_) );
AOI21X1 AOI21X1_360 ( .A(_1796_), .B(micro_hash_ucr_Wx_116_), .C(_2712_), .Y(_2713_) );
NOR2X1 NOR2X1_556 ( .A(_2713_), .B(_292__bF_buf6), .Y(_125__188_) );
OAI21X1 OAI21X1_814 ( .A(_1799_), .B(micro_hash_ucr_Wx_117_), .C(_2104_), .Y(_2714_) );
AOI21X1 AOI21X1_361 ( .A(_1799_), .B(micro_hash_ucr_Wx_117_), .C(_2714_), .Y(_2715_) );
NOR2X1 NOR2X1_557 ( .A(_2715_), .B(_292__bF_buf11), .Y(_125__189_) );
OAI21X1 OAI21X1_815 ( .A(_2204_), .B(micro_hash_ucr_Wx_118_), .C(_2102_), .Y(_2716_) );
AOI21X1 AOI21X1_362 ( .A(_2204_), .B(micro_hash_ucr_Wx_118_), .C(_2716_), .Y(_2717_) );
NOR2X1 NOR2X1_558 ( .A(_2717_), .B(_292__bF_buf9), .Y(_125__190_) );
INVX1 INVX1_331 ( .A(micro_hash_ucr_Wx_79_), .Y(_2718_) );
AOI21X1 AOI21X1_363 ( .A(micro_hash_ucr_Wx_119_), .B(_2718_), .C(micro_hash_ucr_Wx_167_), .Y(_2719_) );
OAI21X1 OAI21X1_816 ( .A(_2718_), .B(micro_hash_ucr_Wx_119_), .C(_2719_), .Y(_2720_) );
AND2X2 AND2X2_122 ( .A(_2720_), .B(_131__bF_buf0), .Y(_125__191_) );
OAI21X1 OAI21X1_817 ( .A(_461_), .B(micro_hash_ucr_Wx_80_), .C(_516_), .Y(_2721_) );
AOI21X1 AOI21X1_364 ( .A(_461_), .B(micro_hash_ucr_Wx_80_), .C(_2721_), .Y(_2722_) );
NOR2X1 NOR2X1_559 ( .A(_2722_), .B(_292__bF_buf8), .Y(_125__152_) );
OAI21X1 OAI21X1_818 ( .A(_631_), .B(micro_hash_ucr_Wx_81_), .C(_709_), .Y(_2723_) );
AOI21X1 AOI21X1_365 ( .A(_631_), .B(micro_hash_ucr_Wx_81_), .C(_2723_), .Y(_2724_) );
NOR2X1 NOR2X1_560 ( .A(_2724_), .B(_292__bF_buf0), .Y(_125__153_) );
OAI21X1 OAI21X1_819 ( .A(_884_), .B(micro_hash_ucr_Wx_82_), .C(_983_), .Y(_2725_) );
AOI21X1 AOI21X1_366 ( .A(_884_), .B(micro_hash_ucr_Wx_82_), .C(_2725_), .Y(_2726_) );
NOR2X1 NOR2X1_561 ( .A(_2726_), .B(_292__bF_buf0), .Y(_125__154_) );
OAI21X1 OAI21X1_820 ( .A(_1229_), .B(micro_hash_ucr_Wx_83_), .C(_1309_), .Y(_2727_) );
AOI21X1 AOI21X1_367 ( .A(_1229_), .B(micro_hash_ucr_Wx_83_), .C(_2727_), .Y(_2728_) );
NOR2X1 NOR2X1_562 ( .A(_2728_), .B(_292__bF_buf12), .Y(_125__155_) );
XNOR2X1 XNOR2X1_205 ( .A(micro_hash_ucr_Wx_44_), .B(micro_hash_ucr_Wx_84_), .Y(_2729_) );
AOI21X1 AOI21X1_368 ( .A(_1555_), .B(_2729_), .C(_292__bF_buf11), .Y(_125__156_) );
OAI21X1 OAI21X1_821 ( .A(_1769_), .B(micro_hash_ucr_Wx_85_), .C(_1838_), .Y(_2730_) );
AOI21X1 AOI21X1_369 ( .A(_1769_), .B(micro_hash_ucr_Wx_85_), .C(_2730_), .Y(_2731_) );
NOR2X1 NOR2X1_563 ( .A(_2731_), .B(_292__bF_buf11), .Y(_125__157_) );
OAI21X1 OAI21X1_822 ( .A(_1977_), .B(micro_hash_ucr_Wx_86_), .C(_2069_), .Y(_2732_) );
AOI21X1 AOI21X1_370 ( .A(_1977_), .B(micro_hash_ucr_Wx_86_), .C(_2732_), .Y(_2733_) );
NOR2X1 NOR2X1_564 ( .A(_2733_), .B(_292__bF_buf6), .Y(_125__158_) );
XNOR2X1 XNOR2X1_206 ( .A(micro_hash_ucr_Wx_47_), .B(micro_hash_ucr_Wx_87_), .Y(_2734_) );
AOI21X1 AOI21X1_371 ( .A(_2295_), .B(_2734_), .C(_292__bF_buf9), .Y(_125__159_) );
AOI21X1 AOI21X1_372 ( .A(micro_hash_ucr_Wx_96_), .B(_471_), .C(micro_hash_ucr_Wx_144_), .Y(_2735_) );
OAI21X1 OAI21X1_823 ( .A(_471_), .B(micro_hash_ucr_Wx_96_), .C(_2735_), .Y(_2736_) );
AND2X2 AND2X2_123 ( .A(_2736_), .B(_131__bF_buf3), .Y(_125__168_) );
OAI21X1 OAI21X1_824 ( .A(_900_), .B(micro_hash_ucr_Wx_97_), .C(_722_), .Y(_2737_) );
AOI21X1 AOI21X1_373 ( .A(_900_), .B(micro_hash_ucr_Wx_97_), .C(_2737_), .Y(_2738_) );
NOR2X1 NOR2X1_565 ( .A(_2738_), .B(_292__bF_buf8), .Y(_125__169_) );
OAI21X1 OAI21X1_825 ( .A(_903_), .B(micro_hash_ucr_Wx_98_), .C(_999_), .Y(_2739_) );
AOI21X1 AOI21X1_374 ( .A(_903_), .B(micro_hash_ucr_Wx_98_), .C(_2739_), .Y(_2740_) );
NOR2X1 NOR2X1_566 ( .A(_2740_), .B(_292__bF_buf3), .Y(_125__170_) );
OAI21X1 OAI21X1_826 ( .A(_1170_), .B(micro_hash_ucr_Wx_99_), .C(_1327_), .Y(_2741_) );
AOI21X1 AOI21X1_375 ( .A(_1170_), .B(micro_hash_ucr_Wx_99_), .C(_2741_), .Y(_2742_) );
NOR2X1 NOR2X1_567 ( .A(_2742_), .B(_292__bF_buf12), .Y(_125__171_) );
OAI21X1 OAI21X1_827 ( .A(_1718_), .B(micro_hash_ucr_Wx_100_), .C(_1850_), .Y(_2743_) );
AOI21X1 AOI21X1_376 ( .A(_1718_), .B(micro_hash_ucr_Wx_100_), .C(_2743_), .Y(_2744_) );
NOR2X1 NOR2X1_568 ( .A(_2744_), .B(_292__bF_buf11), .Y(_125__172_) );
OAI21X1 OAI21X1_828 ( .A(_1996_), .B(micro_hash_ucr_Wx_101_), .C(_2087_), .Y(_2745_) );
AOI21X1 AOI21X1_377 ( .A(_1996_), .B(micro_hash_ucr_Wx_101_), .C(_2745_), .Y(_2746_) );
NOR2X1 NOR2X1_569 ( .A(_2746_), .B(_292__bF_buf6), .Y(_125__173_) );
OAI21X1 OAI21X1_829 ( .A(_1994_), .B(micro_hash_ucr_Wx_102_), .C(_2085_), .Y(_2747_) );
AOI21X1 AOI21X1_378 ( .A(_1994_), .B(micro_hash_ucr_Wx_102_), .C(_2747_), .Y(_2748_) );
NOR2X1 NOR2X1_570 ( .A(_2748_), .B(_292__bF_buf9), .Y(_125__174_) );
AOI21X1 AOI21X1_379 ( .A(micro_hash_ucr_Wx_103_), .B(_2254_), .C(micro_hash_ucr_Wx_151_), .Y(_2749_) );
OAI21X1 OAI21X1_830 ( .A(_2254_), .B(micro_hash_ucr_Wx_103_), .C(_2749_), .Y(_2750_) );
AND2X2 AND2X2_124 ( .A(_2750_), .B(_131__bF_buf0), .Y(_125__175_) );
OAI21X1 OAI21X1_831 ( .A(_467_), .B(micro_hash_ucr_Wx_88_), .C(_523_), .Y(_2751_) );
AOI21X1 AOI21X1_380 ( .A(_467_), .B(micro_hash_ucr_Wx_88_), .C(_2751_), .Y(_2752_) );
NOR2X1 NOR2X1_571 ( .A(_2752_), .B(_292__bF_buf1), .Y(_125__160_) );
OAI21X1 OAI21X1_832 ( .A(_637_), .B(micro_hash_ucr_Wx_89_), .C(_715_), .Y(_2753_) );
AOI21X1 AOI21X1_381 ( .A(_637_), .B(micro_hash_ucr_Wx_89_), .C(_2753_), .Y(_2754_) );
NOR2X1 NOR2X1_572 ( .A(_2754_), .B(_292__bF_buf0), .Y(_125__161_) );
OAI21X1 OAI21X1_833 ( .A(_891_), .B(micro_hash_ucr_Wx_90_), .C(_991_), .Y(_2755_) );
AOI21X1 AOI21X1_382 ( .A(_891_), .B(micro_hash_ucr_Wx_90_), .C(_2755_), .Y(_2756_) );
NOR2X1 NOR2X1_573 ( .A(_2756_), .B(_292__bF_buf0), .Y(_125__162_) );
OAI21X1 OAI21X1_834 ( .A(_1237_), .B(micro_hash_ucr_Wx_91_), .C(_1319_), .Y(_2757_) );
AOI21X1 AOI21X1_383 ( .A(_1237_), .B(micro_hash_ucr_Wx_91_), .C(_2757_), .Y(_2758_) );
NOR2X1 NOR2X1_574 ( .A(_2758_), .B(_292__bF_buf12), .Y(_125__163_) );
OAI21X1 OAI21X1_835 ( .A(_1776_), .B(micro_hash_ucr_Wx_92_), .C(_1563_), .Y(_2759_) );
AOI21X1 AOI21X1_384 ( .A(_1776_), .B(micro_hash_ucr_Wx_92_), .C(_2759_), .Y(_2760_) );
NOR2X1 NOR2X1_575 ( .A(_2760_), .B(_292__bF_buf6), .Y(_125__164_) );
OAI21X1 OAI21X1_836 ( .A(_1778_), .B(micro_hash_ucr_Wx_93_), .C(_2078_), .Y(_2761_) );
AOI21X1 AOI21X1_385 ( .A(_1778_), .B(micro_hash_ucr_Wx_93_), .C(_2761_), .Y(_2762_) );
NOR2X1 NOR2X1_576 ( .A(_2762_), .B(_292__bF_buf11), .Y(_125__165_) );
AOI21X1 AOI21X1_386 ( .A(micro_hash_ucr_Wx_94_), .B(_1985_), .C(micro_hash_ucr_Wx_142_), .Y(_2763_) );
OAI21X1 OAI21X1_837 ( .A(_1985_), .B(micro_hash_ucr_Wx_94_), .C(_2763_), .Y(_2764_) );
AND2X2 AND2X2_125 ( .A(_2764_), .B(_131__bF_buf10), .Y(_125__166_) );
XNOR2X1 XNOR2X1_207 ( .A(micro_hash_ucr_Wx_55_), .B(micro_hash_ucr_Wx_95_), .Y(_2765_) );
AOI21X1 AOI21X1_387 ( .A(_2300_), .B(_2765_), .C(_292__bF_buf9), .Y(_125__167_) );
OAI21X1 OAI21X1_838 ( .A(_449_), .B(micro_hash_ucr_Wx_56_), .C(_503_), .Y(_2766_) );
AOI21X1 AOI21X1_388 ( .A(_449_), .B(micro_hash_ucr_Wx_56_), .C(_2766_), .Y(_2767_) );
NOR2X1 NOR2X1_577 ( .A(_2767_), .B(_292__bF_buf1), .Y(_125__128_) );
OAI21X1 OAI21X1_839 ( .A(_610_), .B(micro_hash_ucr_Wx_57_), .C(_685_), .Y(_2768_) );
AOI21X1 AOI21X1_389 ( .A(_610_), .B(micro_hash_ucr_Wx_57_), .C(_2768_), .Y(_2769_) );
NOR2X1 NOR2X1_578 ( .A(_2769_), .B(_292__bF_buf0), .Y(_125__129_) );
OAI21X1 OAI21X1_840 ( .A(_842_), .B(micro_hash_ucr_Wx_58_), .C(_953_), .Y(_2770_) );
AOI21X1 AOI21X1_390 ( .A(_842_), .B(micro_hash_ucr_Wx_58_), .C(_2770_), .Y(_2771_) );
NOR2X1 NOR2X1_579 ( .A(_2771_), .B(_292__bF_buf3), .Y(_125__130_) );
OAI21X1 OAI21X1_841 ( .A(_1199_), .B(micro_hash_ucr_Wx_59_), .C(_1289_), .Y(_2772_) );
AOI21X1 AOI21X1_391 ( .A(_1199_), .B(micro_hash_ucr_Wx_59_), .C(_2772_), .Y(_2773_) );
NOR2X1 NOR2X1_580 ( .A(_2773_), .B(_292__bF_buf12), .Y(_125__131_) );
OAI21X1 OAI21X1_842 ( .A(_1451_), .B(micro_hash_ucr_Wx_60_), .C(_1532_), .Y(_2774_) );
AOI21X1 AOI21X1_392 ( .A(_1451_), .B(micro_hash_ucr_Wx_60_), .C(_2774_), .Y(_2775_) );
NOR2X1 NOR2X1_581 ( .A(_2775_), .B(_292__bF_buf11), .Y(_125__132_) );
OAI21X1 OAI21X1_843 ( .A(_1744_), .B(micro_hash_ucr_Wx_61_), .C(_2045_), .Y(_2776_) );
AOI21X1 AOI21X1_393 ( .A(_1744_), .B(micro_hash_ucr_Wx_61_), .C(_2776_), .Y(_2777_) );
NOR2X1 NOR2X1_582 ( .A(_2777_), .B(_292__bF_buf6), .Y(_125__133_) );
AOI21X1 AOI21X1_394 ( .A(micro_hash_ucr_Wx_62_), .B(_1957_), .C(micro_hash_ucr_Wx_110_), .Y(_2778_) );
OAI21X1 OAI21X1_844 ( .A(_1957_), .B(micro_hash_ucr_Wx_62_), .C(_2778_), .Y(_2779_) );
AND2X2 AND2X2_126 ( .A(_2779_), .B(_131__bF_buf0), .Y(_125__134_) );
XNOR2X1 XNOR2X1_208 ( .A(micro_hash_ucr_Wx_23_), .B(micro_hash_ucr_Wx_63_), .Y(_2780_) );
AOI21X1 AOI21X1_395 ( .A(_2282_), .B(_2780_), .C(_292__bF_buf9), .Y(_125__135_) );
OAI21X1 OAI21X1_845 ( .A(_455_), .B(micro_hash_ucr_Wx_72_), .C(_512_), .Y(_2781_) );
AOI21X1 AOI21X1_396 ( .A(_455_), .B(micro_hash_ucr_Wx_72_), .C(_2781_), .Y(_2782_) );
NOR2X1 NOR2X1_583 ( .A(_2782_), .B(_292__bF_buf1), .Y(_125__144_) );
OAI21X1 OAI21X1_846 ( .A(_625_), .B(micro_hash_ucr_Wx_73_), .C(_702_), .Y(_2783_) );
AOI21X1 AOI21X1_397 ( .A(_625_), .B(micro_hash_ucr_Wx_73_), .C(_2783_), .Y(_2784_) );
NOR2X1 NOR2X1_584 ( .A(_2784_), .B(_292__bF_buf0), .Y(_125__145_) );
OAI21X1 OAI21X1_847 ( .A(_835_), .B(micro_hash_ucr_Wx_74_), .C(_971_), .Y(_2785_) );
AOI21X1 AOI21X1_398 ( .A(_835_), .B(micro_hash_ucr_Wx_74_), .C(_2785_), .Y(_2786_) );
NOR2X1 NOR2X1_585 ( .A(_2786_), .B(_292__bF_buf0), .Y(_125__146_) );
OAI21X1 OAI21X1_848 ( .A(_1218_), .B(micro_hash_ucr_Wx_75_), .C(_1154_), .Y(_2787_) );
AOI21X1 AOI21X1_399 ( .A(_1218_), .B(micro_hash_ucr_Wx_75_), .C(_2787_), .Y(_2788_) );
NOR2X1 NOR2X1_586 ( .A(_2788_), .B(_292__bF_buf12), .Y(_125__147_) );
OAI21X1 OAI21X1_849 ( .A(_1762_), .B(micro_hash_ucr_Wx_76_), .C(_1703_), .Y(_2789_) );
AOI21X1 AOI21X1_400 ( .A(_1762_), .B(micro_hash_ucr_Wx_76_), .C(_2789_), .Y(_2790_) );
NOR2X1 NOR2X1_587 ( .A(_2790_), .B(_292__bF_buf11), .Y(_125__148_) );
OAI21X1 OAI21X1_850 ( .A(_1972_), .B(micro_hash_ucr_Wx_77_), .C(_1705_), .Y(_2791_) );
AOI21X1 AOI21X1_401 ( .A(_1972_), .B(micro_hash_ucr_Wx_77_), .C(_2791_), .Y(_2792_) );
NOR2X1 NOR2X1_588 ( .A(_2792_), .B(_292__bF_buf11), .Y(_125__149_) );
OAI21X1 OAI21X1_851 ( .A(_1970_), .B(micro_hash_ucr_Wx_78_), .C(_2062_), .Y(_2793_) );
AOI21X1 AOI21X1_402 ( .A(_1970_), .B(micro_hash_ucr_Wx_78_), .C(_2793_), .Y(_2794_) );
NOR2X1 NOR2X1_589 ( .A(_2794_), .B(_292__bF_buf9), .Y(_125__150_) );
XNOR2X1 XNOR2X1_209 ( .A(micro_hash_ucr_Wx_39_), .B(micro_hash_ucr_Wx_79_), .Y(_2795_) );
AOI21X1 AOI21X1_403 ( .A(_2621_), .B(_2795_), .C(_292__bF_buf9), .Y(_125__151_) );
OAI21X1 OAI21X1_852 ( .A(_431_), .B(micro_hash_ucr_Wx_64_), .C(_507_), .Y(_2796_) );
AOI21X1 AOI21X1_404 ( .A(_431_), .B(micro_hash_ucr_Wx_64_), .C(_2796_), .Y(_2797_) );
NOR2X1 NOR2X1_590 ( .A(_2797_), .B(_292__bF_buf1), .Y(_125__136_) );
OAI21X1 OAI21X1_853 ( .A(_616_), .B(micro_hash_ucr_Wx_65_), .C(_961_), .Y(_2798_) );
AOI21X1 AOI21X1_405 ( .A(_616_), .B(micro_hash_ucr_Wx_65_), .C(_2798_), .Y(_2799_) );
NOR2X1 NOR2X1_591 ( .A(_2799_), .B(_292__bF_buf0), .Y(_125__137_) );
OAI21X1 OAI21X1_854 ( .A(_870_), .B(micro_hash_ucr_Wx_66_), .C(_963_), .Y(_2800_) );
AOI21X1 AOI21X1_406 ( .A(_870_), .B(micro_hash_ucr_Wx_66_), .C(_2800_), .Y(_2801_) );
NOR2X1 NOR2X1_592 ( .A(_2801_), .B(_292__bF_buf3), .Y(_125__138_) );
OAI21X1 OAI21X1_855 ( .A(_1209_), .B(micro_hash_ucr_Wx_67_), .C(_1298_), .Y(_2802_) );
AOI21X1 AOI21X1_407 ( .A(_1209_), .B(micro_hash_ucr_Wx_67_), .C(_2802_), .Y(_2803_) );
NOR2X1 NOR2X1_593 ( .A(_2803_), .B(_292__bF_buf12), .Y(_125__139_) );
XNOR2X1 XNOR2X1_210 ( .A(micro_hash_ucr_Wx_28_), .B(micro_hash_ucr_Wx_68_), .Y(_2804_) );
AOI21X1 AOI21X1_408 ( .A(_1828_), .B(_2804_), .C(_292__bF_buf11), .Y(_125__140_) );
OAI21X1 OAI21X1_856 ( .A(_1755_), .B(micro_hash_ucr_Wx_69_), .C(_2054_), .Y(_2805_) );
AOI21X1 AOI21X1_409 ( .A(_1755_), .B(micro_hash_ucr_Wx_69_), .C(_2805_), .Y(_2806_) );
NOR2X1 NOR2X1_594 ( .A(_2806_), .B(_292__bF_buf11), .Y(_125__141_) );
OAI21X1 OAI21X1_857 ( .A(_1963_), .B(micro_hash_ucr_Wx_70_), .C(_2052_), .Y(_2807_) );
AOI21X1 AOI21X1_410 ( .A(_1963_), .B(micro_hash_ucr_Wx_70_), .C(_2807_), .Y(_2808_) );
NOR2X1 NOR2X1_595 ( .A(_2808_), .B(_292__bF_buf9), .Y(_125__142_) );
AOI21X1 AOI21X1_411 ( .A(micro_hash_ucr_Wx_71_), .B(_2231_), .C(micro_hash_ucr_Wx_119_), .Y(_2809_) );
OAI21X1 OAI21X1_858 ( .A(_2231_), .B(micro_hash_ucr_Wx_71_), .C(_2809_), .Y(_2810_) );
AND2X2 AND2X2_127 ( .A(_2810_), .B(_131__bF_buf0), .Y(_125__143_) );
AND2X2 AND2X2_128 ( .A(_131__bF_buf8), .B(concatenador_data_out_104_), .Y(_125__104_) );
AND2X2 AND2X2_129 ( .A(_131__bF_buf11), .B(concatenador_data_out_105_), .Y(_125__105_) );
AND2X2 AND2X2_130 ( .A(_131__bF_buf8), .B(concatenador_data_out_106_), .Y(_125__106_) );
AND2X2 AND2X2_131 ( .A(_131__bF_buf9), .B(concatenador_data_out_107_), .Y(_125__107_) );
AND2X2 AND2X2_132 ( .A(_131__bF_buf7), .B(concatenador_data_out_108_), .Y(_125__108_) );
AND2X2 AND2X2_133 ( .A(_131__bF_buf7), .B(concatenador_data_out_109_), .Y(_125__109_) );
AND2X2 AND2X2_134 ( .A(_131__bF_buf11), .B(concatenador_data_out_110_), .Y(_125__110_) );
AND2X2 AND2X2_135 ( .A(_131__bF_buf4), .B(concatenador_data_out_111_), .Y(_125__111_) );
AND2X2 AND2X2_136 ( .A(_131__bF_buf3), .B(concatenador_data_out_120_), .Y(_125__120_) );
AND2X2 AND2X2_137 ( .A(_131__bF_buf9), .B(concatenador_data_out_121_), .Y(_125__121_) );
AND2X2 AND2X2_138 ( .A(_131__bF_buf8), .B(concatenador_data_out_122_), .Y(_125__122_) );
AND2X2 AND2X2_139 ( .A(_131__bF_buf5), .B(concatenador_data_out_123_), .Y(_125__123_) );
AND2X2 AND2X2_140 ( .A(_131__bF_buf2), .B(concatenador_data_out_124_), .Y(_125__124_) );
AND2X2 AND2X2_141 ( .A(_131__bF_buf5), .B(concatenador_data_out_125_), .Y(_125__125_) );
AND2X2 AND2X2_142 ( .A(_131__bF_buf4), .B(concatenador_data_out_126_), .Y(_125__126_) );
AND2X2 AND2X2_143 ( .A(_131__bF_buf4), .B(concatenador_data_out_127_), .Y(_125__127_) );
AND2X2 AND2X2_144 ( .A(_131__bF_buf12), .B(concatenador_data_out_112_), .Y(_125__112_) );
AND2X2 AND2X2_145 ( .A(_131__bF_buf11), .B(concatenador_data_out_113_), .Y(_125__113_) );
AND2X2 AND2X2_146 ( .A(_131__bF_buf8), .B(concatenador_data_out_114_), .Y(_125__114_) );
AND2X2 AND2X2_147 ( .A(_131__bF_buf9), .B(concatenador_data_out_115_), .Y(_125__115_) );
AND2X2 AND2X2_148 ( .A(_131__bF_buf5), .B(concatenador_data_out_116_), .Y(_125__116_) );
AND2X2 AND2X2_149 ( .A(_131__bF_buf7), .B(concatenador_data_out_117_), .Y(_125__117_) );
AND2X2 AND2X2_150 ( .A(_131__bF_buf2), .B(concatenador_data_out_118_), .Y(_125__118_) );
AND2X2 AND2X2_151 ( .A(_131__bF_buf1), .B(concatenador_data_out_119_), .Y(_125__119_) );
AND2X2 AND2X2_152 ( .A(_131__bF_buf12), .B(concatenador_data_out_80_), .Y(_125__80_) );
AND2X2 AND2X2_153 ( .A(_131__bF_buf9), .B(concatenador_data_out_81_), .Y(_125__81_) );
AND2X2 AND2X2_154 ( .A(_131__bF_buf8), .B(concatenador_data_out_82_), .Y(_125__82_) );
AND2X2 AND2X2_155 ( .A(_131__bF_buf9), .B(concatenador_data_out_83_), .Y(_125__83_) );
AND2X2 AND2X2_156 ( .A(_131__bF_buf2), .B(concatenador_data_out_84_), .Y(_125__84_) );
AND2X2 AND2X2_157 ( .A(_131__bF_buf12), .B(concatenador_data_out_85_), .Y(_125__85_) );
AND2X2 AND2X2_158 ( .A(_131__bF_buf11), .B(concatenador_data_out_86_), .Y(_125__86_) );
AND2X2 AND2X2_159 ( .A(_131__bF_buf1), .B(concatenador_data_out_87_), .Y(_125__87_) );
AND2X2 AND2X2_160 ( .A(_131__bF_buf8), .B(concatenador_data_out_96_), .Y(_125__96_) );
AND2X2 AND2X2_161 ( .A(_131__bF_buf11), .B(concatenador_data_out_97_), .Y(_125__97_) );
AND2X2 AND2X2_162 ( .A(_131__bF_buf8), .B(concatenador_data_out_98_), .Y(_125__98_) );
AND2X2 AND2X2_163 ( .A(_131__bF_buf5), .B(concatenador_data_out_99_), .Y(_125__99_) );
AND2X2 AND2X2_164 ( .A(_131__bF_buf2), .B(concatenador_data_out_100_), .Y(_125__100_) );
AND2X2 AND2X2_165 ( .A(_131__bF_buf10), .B(concatenador_data_out_101_), .Y(_125__101_) );
AND2X2 AND2X2_166 ( .A(_131__bF_buf7), .B(concatenador_data_out_102_), .Y(_125__102_) );
AND2X2 AND2X2_167 ( .A(_131__bF_buf1), .B(concatenador_data_out_103_), .Y(_125__103_) );
AND2X2 AND2X2_168 ( .A(_131__bF_buf12), .B(concatenador_data_out_88_), .Y(_125__88_) );
AND2X2 AND2X2_169 ( .A(_131__bF_buf8), .B(concatenador_data_out_89_), .Y(_125__89_) );
AND2X2 AND2X2_170 ( .A(_131__bF_buf8), .B(concatenador_data_out_90_), .Y(_125__90_) );
AND2X2 AND2X2_171 ( .A(_131__bF_buf5), .B(concatenador_data_out_91_), .Y(_125__91_) );
AND2X2 AND2X2_172 ( .A(_131__bF_buf5), .B(concatenador_data_out_92_), .Y(_125__92_) );
AND2X2 AND2X2_173 ( .A(_131__bF_buf11), .B(concatenador_data_out_93_), .Y(_125__93_) );
AND2X2 AND2X2_174 ( .A(_131__bF_buf7), .B(concatenador_data_out_94_), .Y(_125__94_) );
AND2X2 AND2X2_175 ( .A(_131__bF_buf1), .B(concatenador_data_out_95_), .Y(_125__95_) );
AND2X2 AND2X2_176 ( .A(_131__bF_buf5), .B(concatenador_data_out_56_), .Y(_125__56_) );
AND2X2 AND2X2_177 ( .A(_131__bF_buf12), .B(concatenador_data_out_57_), .Y(_125__57_) );
AND2X2 AND2X2_178 ( .A(_131__bF_buf8), .B(concatenador_data_out_58_), .Y(_125__58_) );
AND2X2 AND2X2_179 ( .A(_131__bF_buf9), .B(concatenador_data_out_59_), .Y(_125__59_) );
AND2X2 AND2X2_180 ( .A(_131__bF_buf11), .B(concatenador_data_out_60_), .Y(_125__60_) );
AND2X2 AND2X2_181 ( .A(_131__bF_buf7), .B(concatenador_data_out_61_), .Y(_125__61_) );
AND2X2 AND2X2_182 ( .A(_131__bF_buf2), .B(concatenador_data_out_62_), .Y(_125__62_) );
AND2X2 AND2X2_183 ( .A(_131__bF_buf1), .B(concatenador_data_out_63_), .Y(_125__63_) );
AND2X2 AND2X2_184 ( .A(_131__bF_buf12), .B(concatenador_data_out_72_), .Y(_125__72_) );
AND2X2 AND2X2_185 ( .A(_131__bF_buf9), .B(concatenador_data_out_73_), .Y(_125__73_) );
AND2X2 AND2X2_186 ( .A(_131__bF_buf8), .B(concatenador_data_out_74_), .Y(_125__74_) );
AND2X2 AND2X2_187 ( .A(_131__bF_buf5), .B(concatenador_data_out_75_), .Y(_125__75_) );
AND2X2 AND2X2_188 ( .A(_131__bF_buf5), .B(concatenador_data_out_76_), .Y(_125__76_) );
AND2X2 AND2X2_189 ( .A(_131__bF_buf11), .B(concatenador_data_out_77_), .Y(_125__77_) );
AND2X2 AND2X2_190 ( .A(_131__bF_buf7), .B(concatenador_data_out_78_), .Y(_125__78_) );
AND2X2 AND2X2_191 ( .A(_131__bF_buf4), .B(concatenador_data_out_79_), .Y(_125__79_) );
AND2X2 AND2X2_192 ( .A(_131__bF_buf9), .B(concatenador_data_out_64_), .Y(_125__64_) );
AND2X2 AND2X2_193 ( .A(_131__bF_buf9), .B(concatenador_data_out_65_), .Y(_125__65_) );
AND2X2 AND2X2_194 ( .A(_131__bF_buf8), .B(concatenador_data_out_66_), .Y(_125__66_) );
AND2X2 AND2X2_195 ( .A(_131__bF_buf5), .B(concatenador_data_out_67_), .Y(_125__67_) );
AND2X2 AND2X2_196 ( .A(_131__bF_buf11), .B(concatenador_data_out_68_), .Y(_125__68_) );
AND2X2 AND2X2_197 ( .A(_131__bF_buf11), .B(concatenador_data_out_69_), .Y(_125__69_) );
AND2X2 AND2X2_198 ( .A(_131__bF_buf4), .B(concatenador_data_out_70_), .Y(_125__70_) );
AND2X2 AND2X2_199 ( .A(_131__bF_buf1), .B(concatenador_data_out_71_), .Y(_125__71_) );
AND2X2 AND2X2_200 ( .A(_131__bF_buf12), .B(concatenador_data_out_32_), .Y(_125__32_) );
AND2X2 AND2X2_201 ( .A(_131__bF_buf5), .B(concatenador_data_out_33_), .Y(_125__33_) );
AND2X2 AND2X2_202 ( .A(_131__bF_buf9), .B(concatenador_data_out_34_), .Y(_125__34_) );
AND2X2 AND2X2_203 ( .A(_131__bF_buf9), .B(concatenador_data_out_35_), .Y(_125__35_) );
AND2X2 AND2X2_204 ( .A(_131__bF_buf5), .B(concatenador_data_out_36_), .Y(_125__36_) );
AND2X2 AND2X2_205 ( .A(_131__bF_buf11), .B(concatenador_data_out_37_), .Y(_125__37_) );
AND2X2 AND2X2_206 ( .A(_131__bF_buf11), .B(concatenador_data_out_38_), .Y(_125__38_) );
AND2X2 AND2X2_207 ( .A(_131__bF_buf2), .B(concatenador_data_out_39_), .Y(_125__39_) );
AND2X2 AND2X2_208 ( .A(_131__bF_buf12), .B(concatenador_data_out_48_), .Y(_125__48_) );
AND2X2 AND2X2_209 ( .A(_131__bF_buf9), .B(concatenador_data_out_49_), .Y(_125__49_) );
AND2X2 AND2X2_210 ( .A(_131__bF_buf11), .B(concatenador_data_out_50_), .Y(_125__50_) );
AND2X2 AND2X2_211 ( .A(_131__bF_buf9), .B(concatenador_data_out_51_), .Y(_125__51_) );
AND2X2 AND2X2_212 ( .A(_131__bF_buf5), .B(concatenador_data_out_52_), .Y(_125__52_) );
AND2X2 AND2X2_213 ( .A(_131__bF_buf2), .B(concatenador_data_out_53_), .Y(_125__53_) );
AND2X2 AND2X2_214 ( .A(_131__bF_buf1), .B(concatenador_data_out_54_), .Y(_125__54_) );
AND2X2 AND2X2_215 ( .A(_131__bF_buf1), .B(concatenador_data_out_55_), .Y(_125__55_) );
AND2X2 AND2X2_216 ( .A(_131__bF_buf12), .B(concatenador_data_out_40_), .Y(_125__40_) );
AND2X2 AND2X2_217 ( .A(_131__bF_buf12), .B(concatenador_data_out_41_), .Y(_125__41_) );
AND2X2 AND2X2_218 ( .A(_131__bF_buf5), .B(concatenador_data_out_42_), .Y(_125__42_) );
AND2X2 AND2X2_219 ( .A(_131__bF_buf9), .B(concatenador_data_out_43_), .Y(_125__43_) );
AND2X2 AND2X2_220 ( .A(_131__bF_buf11), .B(concatenador_data_out_44_), .Y(_125__44_) );
AND2X2 AND2X2_221 ( .A(_131__bF_buf2), .B(concatenador_data_out_45_), .Y(_125__45_) );
AND2X2 AND2X2_222 ( .A(_131__bF_buf7), .B(concatenador_data_out_46_), .Y(_125__46_) );
AND2X2 AND2X2_223 ( .A(_131__bF_buf1), .B(concatenador_data_out_47_), .Y(_125__47_) );
AND2X2 AND2X2_224 ( .A(_131__bF_buf4), .B(concatenador_data_out_8_), .Y(_125__8_) );
AND2X2 AND2X2_225 ( .A(_131__bF_buf7), .B(concatenador_data_out_9_), .Y(_125__9_) );
AND2X2 AND2X2_226 ( .A(_131__bF_buf7), .B(concatenador_data_out_10_), .Y(_125__10_) );
AND2X2 AND2X2_227 ( .A(_131__bF_buf2), .B(concatenador_data_out_11_), .Y(_125__11_) );
AND2X2 AND2X2_228 ( .A(_131__bF_buf7), .B(concatenador_data_out_12_), .Y(_125__12_) );
AND2X2 AND2X2_229 ( .A(_131__bF_buf4), .B(concatenador_data_out_13_), .Y(_125__13_) );
AND2X2 AND2X2_230 ( .A(_131__bF_buf4), .B(concatenador_data_out_14_), .Y(_125__14_) );
AND2X2 AND2X2_231 ( .A(_131__bF_buf1), .B(concatenador_data_out_15_), .Y(_125__15_) );
AND2X2 AND2X2_232 ( .A(_131__bF_buf1), .B(concatenador_data_out_24_), .Y(_125__24_) );
AND2X2 AND2X2_233 ( .A(_131__bF_buf7), .B(concatenador_data_out_25_), .Y(_125__25_) );
AND2X2 AND2X2_234 ( .A(_131__bF_buf2), .B(concatenador_data_out_26_), .Y(_125__26_) );
AND2X2 AND2X2_235 ( .A(_131__bF_buf2), .B(concatenador_data_out_27_), .Y(_125__27_) );
AND2X2 AND2X2_236 ( .A(_131__bF_buf1), .B(concatenador_data_out_28_), .Y(_125__28_) );
AND2X2 AND2X2_237 ( .A(_131__bF_buf1), .B(concatenador_data_out_29_), .Y(_125__29_) );
AND2X2 AND2X2_238 ( .A(_131__bF_buf0), .B(concatenador_data_out_30_), .Y(_125__30_) );
AND2X2 AND2X2_239 ( .A(_131__bF_buf6), .B(concatenador_data_out_31_), .Y(_125__31_) );
AND2X2 AND2X2_240 ( .A(_131__bF_buf4), .B(concatenador_data_out_16_), .Y(_125__16_) );
AND2X2 AND2X2_241 ( .A(_131__bF_buf7), .B(concatenador_data_out_17_), .Y(_125__17_) );
AND2X2 AND2X2_242 ( .A(_131__bF_buf2), .B(concatenador_data_out_18_), .Y(_125__18_) );
AND2X2 AND2X2_243 ( .A(_131__bF_buf4), .B(concatenador_data_out_19_), .Y(_125__19_) );
AND2X2 AND2X2_244 ( .A(_131__bF_buf4), .B(concatenador_data_out_20_), .Y(_125__20_) );
AND2X2 AND2X2_245 ( .A(_131__bF_buf0), .B(concatenador_data_out_21_), .Y(_125__21_) );
AND2X2 AND2X2_246 ( .A(_131__bF_buf6), .B(concatenador_data_out_22_), .Y(_125__22_) );
AND2X2 AND2X2_247 ( .A(_131__bF_buf0), .B(concatenador_data_out_23_), .Y(_125__23_) );
AND2X2 AND2X2_248 ( .A(_131__bF_buf4), .B(concatenador_data_out_0_), .Y(_125__0_) );
AND2X2 AND2X2_249 ( .A(_131__bF_buf4), .B(concatenador_data_out_1_), .Y(_125__1_) );
AND2X2 AND2X2_250 ( .A(_131__bF_buf2), .B(concatenador_data_out_2_), .Y(_125__2_) );
AND2X2 AND2X2_251 ( .A(_131__bF_buf2), .B(concatenador_data_out_3_), .Y(_125__3_) );
AND2X2 AND2X2_252 ( .A(_131__bF_buf7), .B(concatenador_data_out_4_), .Y(_125__4_) );
AND2X2 AND2X2_253 ( .A(_131__bF_buf4), .B(concatenador_data_out_5_), .Y(_125__5_) );
AND2X2 AND2X2_254 ( .A(_131__bF_buf1), .B(concatenador_data_out_6_), .Y(_125__6_) );
AND2X2 AND2X2_255 ( .A(_131__bF_buf0), .B(concatenador_data_out_7_), .Y(_125__7_) );
NOR2X1 NOR2X1_596 ( .A(_2441__bF_buf2), .B(_292__bF_buf2), .Y(_199_) );
NOR2X1 NOR2X1_597 ( .A(_1078__bF_buf1), .B(_292__bF_buf7), .Y(_194_) );
NOR2X1 NOR2X1_598 ( .A(_4199__bF_buf2), .B(_292__bF_buf8), .Y(_196_) );
NOR2X1 NOR2X1_599 ( .A(_4201__bF_buf1), .B(_292__bF_buf7), .Y(_195_) );
NOR2X1 NOR2X1_600 ( .A(_4204_), .B(_292__bF_buf7), .Y(_191_) );
NOR2X1 NOR2X1_601 ( .A(_279_), .B(_292__bF_buf7), .Y(_193_) );
NOR2X1 NOR2X1_602 ( .A(_278__bF_buf0), .B(_292__bF_buf7), .Y(_192_) );
NOR2X1 NOR2X1_603 ( .A(_4210__bF_buf1), .B(_292__bF_buf7), .Y(_188_) );
NOR2X1 NOR2X1_604 ( .A(_4207__bF_buf4), .B(_292__bF_buf7), .Y(_190_) );
NOR2X1 NOR2X1_605 ( .A(_4208_), .B(_292__bF_buf7), .Y(_189_) );
NOR2X1 NOR2X1_606 ( .A(_4212_), .B(_292__bF_buf4), .Y(_184_) );
NOR2X1 NOR2X1_607 ( .A(_269_), .B(_292__bF_buf7), .Y(_187_) );
NOR2X1 NOR2X1_608 ( .A(_4211__bF_buf1), .B(_292__bF_buf7), .Y(_185_) );
NOR2X1 NOR2X1_609 ( .A(_742__bF_buf0), .B(_292__bF_buf4), .Y(_181_) );
NOR2X1 NOR2X1_610 ( .A(_832__bF_buf0), .B(_292__bF_buf7), .Y(_183_) );
INVX8 INVX8_79 ( .A(micro_hash_ucr_pipe55), .Y(_2811_) );
NOR2X1 NOR2X1_611 ( .A(_2811__bF_buf1), .B(_292__bF_buf4), .Y(_182_) );
NOR2X1 NOR2X1_612 ( .A(_255__bF_buf0), .B(_292__bF_buf4), .Y(_178_) );
INVX8 INVX8_80 ( .A(micro_hash_ucr_pipe53_bF_buf0), .Y(_2812_) );
NOR2X1 NOR2X1_613 ( .A(_2812_), .B(_292__bF_buf4), .Y(_180_) );
NOR2X1 NOR2X1_614 ( .A(_4214__bF_buf0), .B(_292__bF_buf4), .Y(_179_) );
NOR2X1 NOR2X1_615 ( .A(_4217__bF_buf3), .B(_292__bF_buf4), .Y(_174_) );
NOR2X1 NOR2X1_616 ( .A(_4215__bF_buf2), .B(_292__bF_buf4), .Y(_177_) );
NOR2X1 NOR2X1_617 ( .A(_304_), .B(_292__bF_buf4), .Y(_176_) );
NOR2X1 NOR2X1_618 ( .A(_336_), .B(_292__bF_buf4), .Y(_171_) );
NOR2X1 NOR2X1_619 ( .A(_249__bF_buf2), .B(_292__bF_buf4), .Y(_173_) );
NOR2X1 NOR2X1_620 ( .A(_4218__bF_buf3), .B(_292__bF_buf8), .Y(_172_) );
NOR2X1 NOR2X1_621 ( .A(_4220__bF_buf2), .B(_292__bF_buf4), .Y(_168_) );
NOR2X1 NOR2X1_622 ( .A(_4219__bF_buf0), .B(_292__bF_buf4), .Y(_170_) );
NOR2X1 NOR2X1_623 ( .A(_242__bF_buf0), .B(_292__bF_buf4), .Y(_169_) );
INVX8 INVX8_81 ( .A(micro_hash_ucr_pipe39), .Y(_2813_) );
NOR2X1 NOR2X1_624 ( .A(_2813__bF_buf1), .B(_292__bF_buf8), .Y(_165_) );
INVX4 INVX4_46 ( .A(micro_hash_ucr_pipe41_bF_buf0), .Y(_2814_) );
NOR2X1 NOR2X1_625 ( .A(_2814_), .B(_292__bF_buf8), .Y(_167_) );
NOR2X1 NOR2X1_626 ( .A(_296__bF_buf3), .B(_292__bF_buf8), .Y(_166_) );
NOR2X1 NOR2X1_627 ( .A(_4224__bF_buf3), .B(_292__bF_buf1), .Y(_161_) );
NOR2X1 NOR2X1_628 ( .A(_701__bF_buf2), .B(_292__bF_buf8), .Y(_163_) );
INVX8 INVX8_82 ( .A(micro_hash_ucr_pipe37_bF_buf3), .Y(_2815_) );
NOR2X1 NOR2X1_629 ( .A(_2815_), .B(_292__bF_buf1), .Y(_162_) );
NOR2X1 NOR2X1_630 ( .A(_318_), .B(_292__bF_buf1), .Y(_158_) );
NOR2X1 NOR2X1_631 ( .A(_230__bF_buf1), .B(_292__bF_buf8), .Y(_160_) );
NOR2X1 NOR2X1_632 ( .A(_4225__bF_buf3), .B(_292__bF_buf7), .Y(_159_) );
NOR2X1 NOR2X1_633 ( .A(_4228__bF_buf4), .B(_292__bF_buf1), .Y(_155_) );
NOR2X1 NOR2X1_634 ( .A(_4226__bF_buf2), .B(_292__bF_buf1), .Y(_157_) );
NOR2X1 NOR2X1_635 ( .A(_317__bF_buf0), .B(_292__bF_buf1), .Y(_156_) );
NOR2X1 NOR2X1_636 ( .A(_4229_), .B(_292__bF_buf5), .Y(_151_) );
NOR2X1 NOR2X1_637 ( .A(_219_), .B(_292__bF_buf6), .Y(_154_) );
NOR2X1 NOR2X1_638 ( .A(_220__bF_buf2), .B(_292__bF_buf6), .Y(_152_) );
NOR2X1 NOR2X1_639 ( .A(_4233__bF_buf1), .B(_292__bF_buf5), .Y(_148_) );
NOR2X1 NOR2X1_640 ( .A(_4230__bF_buf1), .B(_292__bF_buf5), .Y(_150_) );
NOR2X1 NOR2X1_641 ( .A(_389__bF_buf3), .B(_292__bF_buf5), .Y(_149_) );
NOR2X1 NOR2X1_642 ( .A(_4236__bF_buf0), .B(_292__bF_buf10), .Y(_145_) );
NOR2X1 NOR2X1_643 ( .A(_4234__bF_buf0), .B(_292__bF_buf5), .Y(_147_) );
NOR2X1 NOR2X1_644 ( .A(_4262__bF_buf4), .B(_292__bF_buf5), .Y(_146_) );
NOR2X1 NOR2X1_645 ( .A(_624__bF_buf3), .B(_292__bF_buf10), .Y(_141_) );
NOR2X1 NOR2X1_646 ( .A(_4237__bF_buf2), .B(_292__bF_buf10), .Y(_144_) );
INVX8 INVX8_83 ( .A(micro_hash_ucr_pipe19), .Y(_2816_) );
NOR2X1 NOR2X1_647 ( .A(_2816_), .B(_292__bF_buf10), .Y(_143_) );
NOR2X1 NOR2X1_648 ( .A(_4240_), .B(_292__bF_buf7), .Y(_138_) );
NOR2X1 NOR2X1_649 ( .A(_4238__bF_buf3), .B(_292__bF_buf10), .Y(_140_) );
NOR2X1 NOR2X1_650 ( .A(_4239__bF_buf0), .B(_292__bF_buf10), .Y(_139_) );
NOR2X1 NOR2X1_651 ( .A(_4258_), .B(_292__bF_buf2), .Y(_135_) );
NOR2X1 NOR2X1_652 ( .A(_4241__bF_buf3), .B(_292__bF_buf2), .Y(_137_) );
NOR2X1 NOR2X1_653 ( .A(_4242_), .B(_292__bF_buf2), .Y(_136_) );
NOR2X1 NOR2X1_654 ( .A(_4255_), .B(_292__bF_buf10), .Y(_132_) );
NOR2X1 NOR2X1_655 ( .A(_4277_), .B(_292__bF_buf2), .Y(_134_) );
NOR2X1 NOR2X1_656 ( .A(_4243_), .B(_292__bF_buf2), .Y(_133_) );
NOR2X1 NOR2X1_657 ( .A(_4252_), .B(_292__bF_buf10), .Y(_200_) );
NOR2X1 NOR2X1_658 ( .A(_438_), .B(_292__bF_buf10), .Y(_202_) );
NOR2X1 NOR2X1_659 ( .A(_4254_), .B(_292__bF_buf10), .Y(_201_) );
AND2X2 AND2X2_256 ( .A(_131__bF_buf6), .B(micro_hash_ucr_pipe3), .Y(_175_) );
AND2X2 AND2X2_257 ( .A(_131__bF_buf13), .B(micro_hash_ucr_pipe5), .Y(_197_) );
AND2X2 AND2X2_258 ( .A(_131__bF_buf6), .B(micro_hash_ucr_pipe4), .Y(_186_) );
AND2X2 AND2X2_259 ( .A(_131__bF_buf6), .B(micro_hash_ucr_pipe0), .Y(_142_) );
AND2X2 AND2X2_260 ( .A(_131__bF_buf6), .B(micro_hash_ucr_pipe2), .Y(_164_) );
AND2X2 AND2X2_261 ( .A(_131__bF_buf6), .B(micro_hash_ucr_pipe1), .Y(_153_) );
NAND2X1 NAND2X1_345 ( .A(_330_), .B(_2391_), .Y(_2817_) );
NAND2X1 NAND2X1_346 ( .A(micro_hash_ucr_b_0_bF_buf3_), .B(micro_hash_ucr_c_0_bF_buf0_), .Y(_2818_) );
NAND2X1 NAND2X1_347 ( .A(_2818_), .B(_2817_), .Y(_2819_) );
INVX8 INVX8_84 ( .A(_2819_), .Y(_2820_) );
NOR2X1 NOR2X1_660 ( .A(_4218__bF_buf2), .B(_331_), .Y(_2821_) );
NOR2X1 NOR2X1_661 ( .A(_4219__bF_buf3), .B(_331_), .Y(_2822_) );
NOR3X1 NOR3X1_19 ( .A(micro_hash_ucr_pipe7), .B(micro_hash_ucr_pipe8), .C(_4252_), .Y(_2823_) );
NOR2X1 NOR2X1_662 ( .A(micro_hash_ucr_pipe9), .B(H_0_), .Y(_2824_) );
AOI22X1 AOI22X1_15 ( .A(_2823_), .B(_2824_), .C(_4273_), .D(_2819_), .Y(_2825_) );
INVX1 INVX1_332 ( .A(_4261_), .Y(_2826_) );
AND2X2 AND2X2_262 ( .A(_2826_), .B(_2825_), .Y(_2827_) );
OAI22X1 OAI22X1_24 ( .A(_4248_), .B(_2825_), .C(_2827_), .D(micro_hash_ucr_a_0_bF_buf3_), .Y(_2828_) );
OAI21X1 OAI21X1_859 ( .A(_205_), .B(_2819_), .C(_2828_), .Y(_2829_) );
OAI21X1 OAI21X1_860 ( .A(_2819_), .B(_4238__bF_buf0), .C(_624__bF_buf2), .Y(_2830_) );
AOI21X1 AOI21X1_412 ( .A(_4238__bF_buf0), .B(_2829_), .C(_2830_), .Y(_2831_) );
OAI21X1 OAI21X1_861 ( .A(_624__bF_buf2), .B(micro_hash_ucr_a_0_bF_buf2_), .C(_2816_), .Y(_2832_) );
AOI21X1 AOI21X1_413 ( .A(micro_hash_ucr_pipe19), .B(_2820__bF_buf3), .C(micro_hash_ucr_pipe20_bF_buf0), .Y(_2833_) );
OAI21X1 OAI21X1_862 ( .A(_2831_), .B(_2832_), .C(_2833_), .Y(_2834_) );
OAI21X1 OAI21X1_863 ( .A(micro_hash_ucr_a_0_bF_buf1_), .B(_4237__bF_buf0), .C(_2834_), .Y(_2835_) );
AND2X2 AND2X2_263 ( .A(_2835_), .B(_4236__bF_buf3), .Y(_2836_) );
NOR2X1 NOR2X1_663 ( .A(_4236__bF_buf3), .B(_2820__bF_buf3), .Y(_2837_) );
OAI21X1 OAI21X1_864 ( .A(_2836_), .B(_2837_), .C(_4262__bF_buf2), .Y(_2838_) );
OAI21X1 OAI21X1_865 ( .A(micro_hash_ucr_a_0_bF_buf0_), .B(_4262__bF_buf0), .C(_2838_), .Y(_2839_) );
AOI21X1 AOI21X1_414 ( .A(micro_hash_ucr_pipe23), .B(_2820__bF_buf3), .C(micro_hash_ucr_pipe24_bF_buf3), .Y(_2840_) );
OAI21X1 OAI21X1_866 ( .A(_2839_), .B(micro_hash_ucr_pipe23), .C(_2840_), .Y(_2841_) );
AOI21X1 AOI21X1_415 ( .A(micro_hash_ucr_pipe24_bF_buf2), .B(_331_), .C(micro_hash_ucr_pipe25_bF_buf2), .Y(_2842_) );
AND2X2 AND2X2_264 ( .A(_2841_), .B(_2842_), .Y(_2843_) );
OAI21X1 OAI21X1_867 ( .A(_2819_), .B(_389__bF_buf0), .C(_4230__bF_buf1), .Y(_2844_) );
OAI22X1 OAI22X1_25 ( .A(micro_hash_ucr_a_0_bF_buf3_), .B(_4230__bF_buf0), .C(_2843_), .D(_2844_), .Y(_2845_) );
AOI21X1 AOI21X1_416 ( .A(micro_hash_ucr_pipe27_bF_buf1), .B(_2820__bF_buf3), .C(micro_hash_ucr_pipe28_bF_buf0), .Y(_2846_) );
OAI21X1 OAI21X1_868 ( .A(_2845_), .B(micro_hash_ucr_pipe27_bF_buf1), .C(_2846_), .Y(_2847_) );
AOI21X1 AOI21X1_417 ( .A(micro_hash_ucr_pipe28_bF_buf0), .B(_331_), .C(micro_hash_ucr_pipe29), .Y(_2848_) );
AOI22X1 AOI22X1_16 ( .A(micro_hash_ucr_pipe29), .B(_2820__bF_buf3), .C(_2847_), .D(_2848_), .Y(_2849_) );
AOI21X1 AOI21X1_418 ( .A(micro_hash_ucr_a_0_bF_buf2_), .B(micro_hash_ucr_pipe30_bF_buf0), .C(micro_hash_ucr_pipe31_bF_buf3), .Y(_2850_) );
OAI21X1 OAI21X1_869 ( .A(_2849_), .B(micro_hash_ucr_pipe30_bF_buf0), .C(_2850_), .Y(_2851_) );
OAI21X1 OAI21X1_870 ( .A(_317__bF_buf3), .B(_2820__bF_buf2), .C(_2851_), .Y(_2852_) );
NAND2X1 NAND2X1_348 ( .A(_4226__bF_buf3), .B(_2852_), .Y(_2853_) );
OAI21X1 OAI21X1_871 ( .A(micro_hash_ucr_a_0_bF_buf1_), .B(_4226__bF_buf3), .C(_2853_), .Y(_2854_) );
NAND2X1 NAND2X1_349 ( .A(micro_hash_ucr_pipe33_bF_buf3), .B(_2820__bF_buf1), .Y(_2855_) );
OAI21X1 OAI21X1_872 ( .A(_2854_), .B(micro_hash_ucr_pipe33_bF_buf2), .C(_2855_), .Y(_2856_) );
OAI21X1 OAI21X1_873 ( .A(_331_), .B(_4225__bF_buf0), .C(_230__bF_buf2), .Y(_2857_) );
AOI21X1 AOI21X1_419 ( .A(_4225__bF_buf0), .B(_2856_), .C(_2857_), .Y(_2858_) );
NOR2X1 NOR2X1_664 ( .A(_230__bF_buf0), .B(_2820__bF_buf1), .Y(_2859_) );
OAI21X1 OAI21X1_874 ( .A(_2858_), .B(_2859_), .C(_4224__bF_buf2), .Y(_2860_) );
AOI21X1 AOI21X1_420 ( .A(micro_hash_ucr_pipe36_bF_buf0), .B(_331_), .C(micro_hash_ucr_pipe37_bF_buf2), .Y(_2861_) );
OAI21X1 OAI21X1_875 ( .A(_2819_), .B(_2815_), .C(_701__bF_buf0), .Y(_2862_) );
AOI21X1 AOI21X1_421 ( .A(_2861_), .B(_2860_), .C(_2862_), .Y(_2863_) );
NOR2X1 NOR2X1_665 ( .A(micro_hash_ucr_a_0_bF_buf0_), .B(_701__bF_buf3), .Y(_2864_) );
OAI21X1 OAI21X1_876 ( .A(_2863_), .B(_2864_), .C(_2813__bF_buf2), .Y(_2865_) );
NAND2X1 NAND2X1_350 ( .A(micro_hash_ucr_pipe39), .B(_2819_), .Y(_2866_) );
NAND3X1 NAND3X1_101 ( .A(_296__bF_buf0), .B(_2866_), .C(_2865_), .Y(_2867_) );
AOI21X1 AOI21X1_422 ( .A(micro_hash_ucr_pipe40_bF_buf0), .B(micro_hash_ucr_a_0_bF_buf3_), .C(micro_hash_ucr_pipe41_bF_buf2), .Y(_2868_) );
OAI21X1 OAI21X1_877 ( .A(_2820__bF_buf1), .B(_2814_), .C(_4220__bF_buf3), .Y(_2869_) );
AOI21X1 AOI21X1_423 ( .A(_2868_), .B(_2867_), .C(_2869_), .Y(_2870_) );
NOR2X1 NOR2X1_666 ( .A(_4220__bF_buf2), .B(_331_), .Y(_2871_) );
OAI21X1 OAI21X1_878 ( .A(_2870_), .B(_2871_), .C(_242__bF_buf2), .Y(_2872_) );
NAND2X1 NAND2X1_351 ( .A(micro_hash_ucr_pipe43), .B(_2820__bF_buf1), .Y(_2873_) );
AOI21X1 AOI21X1_424 ( .A(_2873_), .B(_2872_), .C(micro_hash_ucr_pipe44_bF_buf2), .Y(_2874_) );
OAI21X1 OAI21X1_879 ( .A(_2874_), .B(_2822_), .C(_336_), .Y(_2875_) );
NAND2X1 NAND2X1_352 ( .A(micro_hash_ucr_pipe45), .B(_2820__bF_buf1), .Y(_2876_) );
AOI21X1 AOI21X1_425 ( .A(_2876_), .B(_2875_), .C(micro_hash_ucr_pipe46_bF_buf1), .Y(_2877_) );
OAI21X1 OAI21X1_880 ( .A(_2877_), .B(_2821_), .C(_249__bF_buf1), .Y(_2878_) );
AOI21X1 AOI21X1_426 ( .A(micro_hash_ucr_pipe47), .B(_2820__bF_buf0), .C(micro_hash_ucr_pipe48_bF_buf4), .Y(_2879_) );
OAI21X1 OAI21X1_881 ( .A(_4217__bF_buf2), .B(micro_hash_ucr_a_0_bF_buf2_), .C(_304_), .Y(_2880_) );
AOI21X1 AOI21X1_427 ( .A(_2879_), .B(_2878_), .C(_2880_), .Y(_2881_) );
OAI21X1 OAI21X1_882 ( .A(_2819_), .B(_304_), .C(_4215__bF_buf0), .Y(_2882_) );
OAI22X1 OAI22X1_26 ( .A(_4215__bF_buf0), .B(micro_hash_ucr_a_0_bF_buf1_), .C(_2881_), .D(_2882_), .Y(_2883_) );
OAI21X1 OAI21X1_883 ( .A(_2820__bF_buf0), .B(_255__bF_buf1), .C(_4214__bF_buf4), .Y(_2884_) );
AOI21X1 AOI21X1_428 ( .A(_255__bF_buf1), .B(_2883_), .C(_2884_), .Y(_2885_) );
NOR2X1 NOR2X1_667 ( .A(_4214__bF_buf4), .B(_331_), .Y(_2886_) );
OAI21X1 OAI21X1_884 ( .A(_2885_), .B(_2886_), .C(_2812_), .Y(_2887_) );
AOI21X1 AOI21X1_429 ( .A(micro_hash_ucr_pipe53_bF_buf1), .B(_2820__bF_buf0), .C(micro_hash_ucr_pipe54_bF_buf4), .Y(_2888_) );
OAI21X1 OAI21X1_885 ( .A(_742__bF_buf1), .B(micro_hash_ucr_a_0_bF_buf0_), .C(_2811__bF_buf2), .Y(_2889_) );
AOI21X1 AOI21X1_430 ( .A(_2888_), .B(_2887_), .C(_2889_), .Y(_2890_) );
OAI21X1 OAI21X1_886 ( .A(_2819_), .B(_2811__bF_buf2), .C(_832__bF_buf4), .Y(_2891_) );
OAI22X1 OAI22X1_27 ( .A(_832__bF_buf4), .B(micro_hash_ucr_a_0_bF_buf3_), .C(_2890_), .D(_2891_), .Y(_2892_) );
NAND2X1 NAND2X1_353 ( .A(micro_hash_ucr_pipe57_bF_buf2), .B(_2820__bF_buf0), .Y(_2893_) );
OAI21X1 OAI21X1_887 ( .A(_2892_), .B(micro_hash_ucr_pipe57_bF_buf2), .C(_2893_), .Y(_2894_) );
NAND2X1 NAND2X1_354 ( .A(micro_hash_ucr_pipe58_bF_buf3), .B(_331_), .Y(_2895_) );
OAI21X1 OAI21X1_888 ( .A(_2894_), .B(micro_hash_ucr_pipe58_bF_buf3), .C(_2895_), .Y(_2896_) );
NAND2X1 NAND2X1_355 ( .A(micro_hash_ucr_pipe59), .B(_2820__bF_buf2), .Y(_2897_) );
OAI21X1 OAI21X1_889 ( .A(_2896_), .B(micro_hash_ucr_pipe59), .C(_2897_), .Y(_2898_) );
NAND2X1 NAND2X1_356 ( .A(micro_hash_ucr_pipe60_bF_buf4), .B(_331_), .Y(_2899_) );
OAI21X1 OAI21X1_890 ( .A(_2898_), .B(micro_hash_ucr_pipe60_bF_buf4), .C(_2899_), .Y(_2900_) );
NAND2X1 NAND2X1_357 ( .A(micro_hash_ucr_pipe61_bF_buf3), .B(_2820__bF_buf2), .Y(_2901_) );
OAI21X1 OAI21X1_891 ( .A(_2900_), .B(micro_hash_ucr_pipe61_bF_buf3), .C(_2901_), .Y(_2902_) );
NAND2X1 NAND2X1_358 ( .A(micro_hash_ucr_pipe62_bF_buf0), .B(_331_), .Y(_2903_) );
OAI21X1 OAI21X1_892 ( .A(_2902_), .B(micro_hash_ucr_pipe62_bF_buf0), .C(_2903_), .Y(_2904_) );
AOI21X1 AOI21X1_431 ( .A(micro_hash_ucr_pipe63_bF_buf3), .B(_2820__bF_buf2), .C(micro_hash_ucr_pipe64_bF_buf1), .Y(_2905_) );
OAI21X1 OAI21X1_893 ( .A(_2904_), .B(micro_hash_ucr_pipe63_bF_buf3), .C(_2905_), .Y(_2906_) );
AOI21X1 AOI21X1_432 ( .A(micro_hash_ucr_pipe64_bF_buf1), .B(_331_), .C(micro_hash_ucr_pipe65_bF_buf4), .Y(_2907_) );
AOI22X1 AOI22X1_17 ( .A(micro_hash_ucr_pipe65_bF_buf4), .B(_2820__bF_buf2), .C(_2906_), .D(_2907_), .Y(_2908_) );
AOI21X1 AOI21X1_433 ( .A(micro_hash_ucr_pipe66_bF_buf0), .B(micro_hash_ucr_a_0_bF_buf2_), .C(micro_hash_ucr_pipe67), .Y(_2909_) );
OAI21X1 OAI21X1_894 ( .A(_2908_), .B(micro_hash_ucr_pipe66_bF_buf0), .C(_2909_), .Y(_2910_) );
NAND2X1 NAND2X1_359 ( .A(micro_hash_ucr_pipe67), .B(_2819_), .Y(_2911_) );
AOI21X1 AOI21X1_434 ( .A(_2911_), .B(_2910_), .C(micro_hash_ucr_pipe68), .Y(_2912_) );
OAI21X1 OAI21X1_895 ( .A(_4199__bF_buf4), .B(micro_hash_ucr_a_0_bF_buf1_), .C(_344_), .Y(_2913_) );
OAI22X1 OAI22X1_28 ( .A(_2181_), .B(_2819_), .C(_2912_), .D(_2913_), .Y(_126__0_) );
NAND2X1 NAND2X1_360 ( .A(_2448_), .B(_591__bF_buf0), .Y(_2914_) );
NAND2X1 NAND2X1_361 ( .A(micro_hash_ucr_b_1_bF_buf3_), .B(micro_hash_ucr_c_1_bF_buf1_), .Y(_2915_) );
NAND2X1 NAND2X1_362 ( .A(_2915_), .B(_2914_), .Y(_2916_) );
NOR2X1 NOR2X1_668 ( .A(_4211__bF_buf1), .B(_2514__bF_buf1), .Y(_2917_) );
NOR2X1 NOR2X1_669 ( .A(_832__bF_buf0), .B(_2514__bF_buf1), .Y(_2918_) );
NOR2X1 NOR2X1_670 ( .A(_296__bF_buf3), .B(_2514__bF_buf3), .Y(_2919_) );
NAND2X1 NAND2X1_363 ( .A(micro_hash_ucr_a_1_), .B(micro_hash_ucr_pipe34_bF_buf1), .Y(_2920_) );
NAND2X1 NAND2X1_364 ( .A(micro_hash_ucr_pipe28_bF_buf2), .B(_2514__bF_buf1), .Y(_2921_) );
OAI21X1 OAI21X1_896 ( .A(micro_hash_ucr_pipe7), .B(micro_hash_ucr_pipe6), .C(_438_), .Y(_2922_) );
AOI21X1 AOI21X1_435 ( .A(_4255_), .B(_2922_), .C(micro_hash_ucr_pipe10), .Y(_2923_) );
NAND2X1 NAND2X1_365 ( .A(micro_hash_ucr_pipe7), .B(_438_), .Y(_2924_) );
NAND3X1 NAND3X1_102 ( .A(_4255_), .B(_4277_), .C(_2924_), .Y(_2925_) );
NOR2X1 NOR2X1_671 ( .A(micro_hash_ucr_pipe9), .B(H_1_), .Y(_2926_) );
AOI22X1 AOI22X1_18 ( .A(_2823_), .B(_2926_), .C(_2925_), .D(_2916_), .Y(_2927_) );
OAI22X1 OAI22X1_29 ( .A(micro_hash_ucr_a_1_), .B(_2923_), .C(_2927_), .D(_4244_), .Y(_2928_) );
OAI21X1 OAI21X1_897 ( .A(_4277_), .B(_2916_), .C(_2928_), .Y(_2929_) );
NAND2X1 NAND2X1_366 ( .A(micro_hash_ucr_pipe12_bF_buf3), .B(_2514__bF_buf2), .Y(_2930_) );
OAI21X1 OAI21X1_898 ( .A(_2929_), .B(micro_hash_ucr_pipe12_bF_buf3), .C(_2930_), .Y(_2931_) );
INVX8 INVX8_85 ( .A(_2916_), .Y(_2932_) );
NAND2X1 NAND2X1_367 ( .A(micro_hash_ucr_pipe13), .B(_2932__bF_buf1), .Y(_2933_) );
OAI21X1 OAI21X1_899 ( .A(_2931_), .B(micro_hash_ucr_pipe13), .C(_2933_), .Y(_2934_) );
NAND2X1 NAND2X1_368 ( .A(micro_hash_ucr_pipe14), .B(_2514__bF_buf2), .Y(_2935_) );
OAI21X1 OAI21X1_900 ( .A(_2934_), .B(micro_hash_ucr_pipe14), .C(_2935_), .Y(_2936_) );
NAND2X1 NAND2X1_369 ( .A(micro_hash_ucr_pipe15), .B(_2932__bF_buf1), .Y(_2937_) );
OAI21X1 OAI21X1_901 ( .A(_2936_), .B(micro_hash_ucr_pipe15), .C(_2937_), .Y(_2938_) );
NAND2X1 NAND2X1_370 ( .A(micro_hash_ucr_pipe16), .B(_2514__bF_buf2), .Y(_2939_) );
OAI21X1 OAI21X1_902 ( .A(_2938_), .B(micro_hash_ucr_pipe16), .C(_2939_), .Y(_2940_) );
NAND2X1 NAND2X1_371 ( .A(micro_hash_ucr_pipe17), .B(_2932__bF_buf1), .Y(_2941_) );
OAI21X1 OAI21X1_903 ( .A(_2940_), .B(micro_hash_ucr_pipe17), .C(_2941_), .Y(_2942_) );
NAND2X1 NAND2X1_372 ( .A(micro_hash_ucr_pipe18_bF_buf4), .B(_2514__bF_buf2), .Y(_2943_) );
OAI21X1 OAI21X1_904 ( .A(_2942_), .B(micro_hash_ucr_pipe18_bF_buf4), .C(_2943_), .Y(_2944_) );
NAND2X1 NAND2X1_373 ( .A(micro_hash_ucr_pipe19), .B(_2932__bF_buf1), .Y(_2945_) );
OAI21X1 OAI21X1_905 ( .A(_2944_), .B(micro_hash_ucr_pipe19), .C(_2945_), .Y(_2946_) );
AOI21X1 AOI21X1_436 ( .A(micro_hash_ucr_pipe20_bF_buf2), .B(_2514__bF_buf0), .C(micro_hash_ucr_pipe21), .Y(_2947_) );
OAI21X1 OAI21X1_906 ( .A(_2946_), .B(micro_hash_ucr_pipe20_bF_buf2), .C(_2947_), .Y(_2948_) );
AOI21X1 AOI21X1_437 ( .A(micro_hash_ucr_pipe21), .B(_2932__bF_buf1), .C(micro_hash_ucr_pipe22_bF_buf2), .Y(_2949_) );
AOI22X1 AOI22X1_19 ( .A(_2514__bF_buf0), .B(micro_hash_ucr_pipe22_bF_buf2), .C(_2948_), .D(_2949_), .Y(_2950_) );
OAI21X1 OAI21X1_907 ( .A(_2916_), .B(_4234__bF_buf0), .C(_4233__bF_buf4), .Y(_2951_) );
AOI21X1 AOI21X1_438 ( .A(_4234__bF_buf0), .B(_2950_), .C(_2951_), .Y(_2952_) );
OAI21X1 OAI21X1_908 ( .A(_4233__bF_buf2), .B(micro_hash_ucr_a_1_), .C(_389__bF_buf3), .Y(_2953_) );
AOI21X1 AOI21X1_439 ( .A(micro_hash_ucr_pipe25_bF_buf0), .B(_2932__bF_buf2), .C(micro_hash_ucr_pipe26_bF_buf1), .Y(_2954_) );
OAI21X1 OAI21X1_909 ( .A(_2952_), .B(_2953_), .C(_2954_), .Y(_2955_) );
NAND2X1 NAND2X1_374 ( .A(micro_hash_ucr_pipe26_bF_buf1), .B(_2514__bF_buf0), .Y(_2956_) );
AOI21X1 AOI21X1_440 ( .A(_2956_), .B(_2955_), .C(micro_hash_ucr_pipe27_bF_buf1), .Y(_2957_) );
NOR2X1 NOR2X1_672 ( .A(_4229_), .B(_2932__bF_buf2), .Y(_2958_) );
OAI21X1 OAI21X1_910 ( .A(_2957_), .B(_2958_), .C(_220__bF_buf1), .Y(_2959_) );
NAND3X1 NAND3X1_103 ( .A(_219_), .B(_2921_), .C(_2959_), .Y(_2960_) );
NAND2X1 NAND2X1_375 ( .A(micro_hash_ucr_pipe29), .B(_2932__bF_buf0), .Y(_2961_) );
AOI21X1 AOI21X1_441 ( .A(_2961_), .B(_2960_), .C(micro_hash_ucr_pipe30_bF_buf3), .Y(_2962_) );
OAI21X1 OAI21X1_911 ( .A(_2514__bF_buf1), .B(_4228__bF_buf1), .C(_317__bF_buf2), .Y(_2963_) );
AOI21X1 AOI21X1_442 ( .A(micro_hash_ucr_pipe31_bF_buf2), .B(_2916_), .C(micro_hash_ucr_pipe32_bF_buf2), .Y(_2964_) );
OAI21X1 OAI21X1_912 ( .A(_2962_), .B(_2963_), .C(_2964_), .Y(_2965_) );
NAND2X1 NAND2X1_376 ( .A(micro_hash_ucr_a_1_), .B(micro_hash_ucr_pipe32_bF_buf0), .Y(_2966_) );
AOI21X1 AOI21X1_443 ( .A(_2966_), .B(_2965_), .C(micro_hash_ucr_pipe33_bF_buf0), .Y(_2967_) );
NOR2X1 NOR2X1_673 ( .A(_318_), .B(_2916_), .Y(_2968_) );
OAI21X1 OAI21X1_913 ( .A(_2967_), .B(_2968_), .C(_4225__bF_buf4), .Y(_2969_) );
AOI21X1 AOI21X1_444 ( .A(_2920_), .B(_2969_), .C(micro_hash_ucr_pipe35), .Y(_2970_) );
NOR2X1 NOR2X1_674 ( .A(_230__bF_buf2), .B(_2916_), .Y(_2971_) );
OAI21X1 OAI21X1_914 ( .A(_2970_), .B(_2971_), .C(_4224__bF_buf3), .Y(_2972_) );
AOI21X1 AOI21X1_445 ( .A(micro_hash_ucr_a_1_), .B(micro_hash_ucr_pipe36_bF_buf3), .C(micro_hash_ucr_pipe37_bF_buf3), .Y(_2973_) );
OAI21X1 OAI21X1_915 ( .A(_2932__bF_buf0), .B(_2815_), .C(_701__bF_buf0), .Y(_2974_) );
AOI21X1 AOI21X1_446 ( .A(_2973_), .B(_2972_), .C(_2974_), .Y(_2975_) );
NOR2X1 NOR2X1_675 ( .A(_2514__bF_buf3), .B(_701__bF_buf1), .Y(_2976_) );
OAI21X1 OAI21X1_916 ( .A(_2975_), .B(_2976_), .C(_2813__bF_buf1), .Y(_2977_) );
NAND2X1 NAND2X1_377 ( .A(micro_hash_ucr_pipe39), .B(_2932__bF_buf0), .Y(_2978_) );
AOI21X1 AOI21X1_447 ( .A(_2978_), .B(_2977_), .C(micro_hash_ucr_pipe40_bF_buf1), .Y(_2979_) );
OAI21X1 OAI21X1_917 ( .A(_2979_), .B(_2919_), .C(_2814_), .Y(_2980_) );
NAND2X1 NAND2X1_378 ( .A(micro_hash_ucr_pipe41_bF_buf3), .B(_2932__bF_buf0), .Y(_2981_) );
AOI21X1 AOI21X1_448 ( .A(_2981_), .B(_2980_), .C(micro_hash_ucr_pipe42_bF_buf0), .Y(_2982_) );
OAI21X1 OAI21X1_918 ( .A(_4220__bF_buf2), .B(_2514__bF_buf3), .C(_242__bF_buf0), .Y(_2983_) );
AOI21X1 AOI21X1_449 ( .A(micro_hash_ucr_pipe43), .B(_2916_), .C(micro_hash_ucr_pipe44_bF_buf2), .Y(_2984_) );
OAI21X1 OAI21X1_919 ( .A(_2982_), .B(_2983_), .C(_2984_), .Y(_2985_) );
OAI21X1 OAI21X1_920 ( .A(_4219__bF_buf4), .B(_2514__bF_buf3), .C(_2985_), .Y(_2986_) );
OAI21X1 OAI21X1_921 ( .A(_2916_), .B(_336_), .C(_4218__bF_buf2), .Y(_2987_) );
AOI21X1 AOI21X1_450 ( .A(_336_), .B(_2986_), .C(_2987_), .Y(_2988_) );
OAI21X1 OAI21X1_922 ( .A(_4218__bF_buf2), .B(micro_hash_ucr_a_1_), .C(_249__bF_buf3), .Y(_2989_) );
AOI21X1 AOI21X1_451 ( .A(micro_hash_ucr_pipe47), .B(_2932__bF_buf3), .C(micro_hash_ucr_pipe48_bF_buf0), .Y(_2990_) );
OAI21X1 OAI21X1_923 ( .A(_2988_), .B(_2989_), .C(_2990_), .Y(_2991_) );
NAND2X1 NAND2X1_379 ( .A(micro_hash_ucr_pipe48_bF_buf0), .B(_2514__bF_buf3), .Y(_2992_) );
NAND3X1 NAND3X1_104 ( .A(_304_), .B(_2992_), .C(_2991_), .Y(_2993_) );
AOI21X1 AOI21X1_452 ( .A(micro_hash_ucr_pipe49_bF_buf1), .B(_2932__bF_buf3), .C(micro_hash_ucr_pipe50_bF_buf3), .Y(_2994_) );
OAI21X1 OAI21X1_924 ( .A(_4215__bF_buf1), .B(micro_hash_ucr_a_1_), .C(_255__bF_buf0), .Y(_2995_) );
AOI21X1 AOI21X1_453 ( .A(_2994_), .B(_2993_), .C(_2995_), .Y(_2996_) );
OAI21X1 OAI21X1_925 ( .A(_2916_), .B(_255__bF_buf2), .C(_4214__bF_buf2), .Y(_2997_) );
OAI22X1 OAI22X1_30 ( .A(_4214__bF_buf2), .B(micro_hash_ucr_a_1_), .C(_2996_), .D(_2997_), .Y(_2998_) );
OAI21X1 OAI21X1_926 ( .A(_2932__bF_buf3), .B(_2812_), .C(_742__bF_buf0), .Y(_2999_) );
AOI21X1 AOI21X1_454 ( .A(_2812_), .B(_2998_), .C(_2999_), .Y(_3000_) );
NOR2X1 NOR2X1_676 ( .A(_742__bF_buf0), .B(_2514__bF_buf1), .Y(_3001_) );
OAI21X1 OAI21X1_927 ( .A(_3000_), .B(_3001_), .C(_2811__bF_buf1), .Y(_3002_) );
NAND2X1 NAND2X1_380 ( .A(micro_hash_ucr_pipe55), .B(_2932__bF_buf3), .Y(_3003_) );
AOI21X1 AOI21X1_455 ( .A(_3003_), .B(_3002_), .C(micro_hash_ucr_pipe56_bF_buf2), .Y(_3004_) );
OAI21X1 OAI21X1_928 ( .A(_3004_), .B(_2918_), .C(_4212_), .Y(_3005_) );
NAND2X1 NAND2X1_381 ( .A(micro_hash_ucr_pipe57_bF_buf0), .B(_2932__bF_buf3), .Y(_3006_) );
AOI21X1 AOI21X1_456 ( .A(_3006_), .B(_3005_), .C(micro_hash_ucr_pipe58_bF_buf0), .Y(_3007_) );
OAI21X1 OAI21X1_929 ( .A(_3007_), .B(_2917_), .C(_269_), .Y(_3008_) );
AOI21X1 AOI21X1_457 ( .A(micro_hash_ucr_pipe59), .B(_2932__bF_buf2), .C(micro_hash_ucr_pipe60_bF_buf1), .Y(_3009_) );
OAI21X1 OAI21X1_930 ( .A(_4210__bF_buf1), .B(micro_hash_ucr_a_1_), .C(_4208_), .Y(_3010_) );
AOI21X1 AOI21X1_458 ( .A(_3009_), .B(_3008_), .C(_3010_), .Y(_3011_) );
OAI21X1 OAI21X1_931 ( .A(_2916_), .B(_4208_), .C(_4207__bF_buf4), .Y(_3012_) );
OAI22X1 OAI22X1_31 ( .A(_4207__bF_buf4), .B(micro_hash_ucr_a_1_), .C(_3011_), .D(_3012_), .Y(_3013_) );
NAND2X1 NAND2X1_382 ( .A(micro_hash_ucr_pipe63_bF_buf1), .B(_2932__bF_buf2), .Y(_3014_) );
OAI21X1 OAI21X1_932 ( .A(_3013_), .B(micro_hash_ucr_pipe63_bF_buf1), .C(_3014_), .Y(_3015_) );
NAND2X1 NAND2X1_383 ( .A(micro_hash_ucr_pipe64_bF_buf4), .B(_2514__bF_buf0), .Y(_3016_) );
OAI21X1 OAI21X1_933 ( .A(_3015_), .B(micro_hash_ucr_pipe64_bF_buf4), .C(_3016_), .Y(_3017_) );
AOI21X1 AOI21X1_459 ( .A(micro_hash_ucr_pipe65_bF_buf1), .B(_2932__bF_buf2), .C(micro_hash_ucr_pipe66_bF_buf4), .Y(_3018_) );
OAI21X1 OAI21X1_934 ( .A(_3017_), .B(micro_hash_ucr_pipe65_bF_buf1), .C(_3018_), .Y(_3019_) );
AOI21X1 AOI21X1_460 ( .A(micro_hash_ucr_pipe66_bF_buf0), .B(_2514__bF_buf0), .C(micro_hash_ucr_pipe67), .Y(_3020_) );
OAI21X1 OAI21X1_935 ( .A(_2916_), .B(_4201__bF_buf1), .C(_4199__bF_buf3), .Y(_3021_) );
AOI21X1 AOI21X1_461 ( .A(_3020_), .B(_3019_), .C(_3021_), .Y(_3022_) );
OAI21X1 OAI21X1_936 ( .A(_4199__bF_buf3), .B(micro_hash_ucr_a_1_), .C(_344_), .Y(_3023_) );
OAI22X1 OAI22X1_32 ( .A(_2181_), .B(_2916_), .C(_3022_), .D(_3023_), .Y(_126__1_) );
NAND2X1 NAND2X1_384 ( .A(micro_hash_ucr_pipe66_bF_buf4), .B(micro_hash_ucr_a_2_bF_buf0_), .Y(_3024_) );
NAND2X1 NAND2X1_385 ( .A(micro_hash_ucr_pipe58_bF_buf0), .B(micro_hash_ucr_a_2_bF_buf4_), .Y(_3025_) );
NAND2X1 NAND2X1_386 ( .A(micro_hash_ucr_pipe56_bF_buf2), .B(micro_hash_ucr_a_2_bF_buf3_), .Y(_3026_) );
NAND2X1 NAND2X1_387 ( .A(micro_hash_ucr_pipe48_bF_buf0), .B(micro_hash_ucr_a_2_bF_buf2_), .Y(_3027_) );
NAND2X1 NAND2X1_388 ( .A(micro_hash_ucr_pipe46_bF_buf4), .B(micro_hash_ucr_a_2_bF_buf1_), .Y(_3028_) );
NAND2X1 NAND2X1_389 ( .A(micro_hash_ucr_pipe44_bF_buf2), .B(micro_hash_ucr_a_2_bF_buf0_), .Y(_3029_) );
NAND2X1 NAND2X1_390 ( .A(micro_hash_ucr_pipe42_bF_buf4), .B(micro_hash_ucr_a_2_bF_buf4_), .Y(_3030_) );
NAND2X1 NAND2X1_391 ( .A(micro_hash_ucr_a_2_bF_buf3_), .B(micro_hash_ucr_pipe24_bF_buf3), .Y(_3031_) );
INVX4 INVX4_47 ( .A(micro_hash_ucr_a_2_bF_buf2_), .Y(_3032_) );
NAND2X1 NAND2X1_392 ( .A(micro_hash_ucr_pipe18_bF_buf4), .B(_3032_), .Y(_3033_) );
NAND2X1 NAND2X1_393 ( .A(micro_hash_ucr_pipe16), .B(_3032_), .Y(_3034_) );
NAND2X1 NAND2X1_394 ( .A(micro_hash_ucr_pipe14), .B(_3032_), .Y(_3035_) );
NAND2X1 NAND2X1_395 ( .A(micro_hash_ucr_pipe12_bF_buf3), .B(_3032_), .Y(_3036_) );
XNOR2X1 XNOR2X1_211 ( .A(micro_hash_ucr_b_2_bF_buf3_), .B(micro_hash_ucr_c_2_bF_buf0_), .Y(_3037_) );
INVX8 INVX8_86 ( .A(_3037__bF_buf2), .Y(_3038_) );
NAND2X1 NAND2X1_396 ( .A(micro_hash_ucr_pipe11), .B(_3038_), .Y(_3039_) );
NOR2X1 NOR2X1_677 ( .A(micro_hash_ucr_pipe9), .B(H_2_), .Y(_3040_) );
AOI22X1 AOI22X1_20 ( .A(_2823_), .B(_3040_), .C(_2925_), .D(_3037__bF_buf1), .Y(_3041_) );
OAI22X1 OAI22X1_33 ( .A(micro_hash_ucr_a_2_bF_buf1_), .B(_2923_), .C(_3041_), .D(_4244_), .Y(_3042_) );
NAND3X1 NAND3X1_105 ( .A(_4258_), .B(_3039_), .C(_3042_), .Y(_3043_) );
NAND3X1 NAND3X1_106 ( .A(_4242_), .B(_3036_), .C(_3043_), .Y(_3044_) );
NAND2X1 NAND2X1_397 ( .A(micro_hash_ucr_pipe13), .B(_3038_), .Y(_3045_) );
NAND3X1 NAND3X1_107 ( .A(_4241__bF_buf3), .B(_3045_), .C(_3044_), .Y(_3046_) );
NAND3X1 NAND3X1_108 ( .A(_4240_), .B(_3035_), .C(_3046_), .Y(_3047_) );
NAND2X1 NAND2X1_398 ( .A(micro_hash_ucr_pipe15), .B(_3038_), .Y(_3048_) );
NAND3X1 NAND3X1_109 ( .A(_4239__bF_buf3), .B(_3048_), .C(_3047_), .Y(_3049_) );
NAND3X1 NAND3X1_110 ( .A(_4238__bF_buf2), .B(_3034_), .C(_3049_), .Y(_3050_) );
NAND2X1 NAND2X1_399 ( .A(micro_hash_ucr_pipe17), .B(_3038_), .Y(_3051_) );
NAND3X1 NAND3X1_111 ( .A(_624__bF_buf1), .B(_3051_), .C(_3050_), .Y(_3052_) );
NAND3X1 NAND3X1_112 ( .A(_2816_), .B(_3033_), .C(_3052_), .Y(_3053_) );
AOI21X1 AOI21X1_462 ( .A(micro_hash_ucr_pipe19), .B(_3038_), .C(micro_hash_ucr_pipe20_bF_buf0), .Y(_3054_) );
OAI21X1 OAI21X1_937 ( .A(_4237__bF_buf0), .B(micro_hash_ucr_a_2_bF_buf0_), .C(_4236__bF_buf2), .Y(_3055_) );
AOI21X1 AOI21X1_463 ( .A(_3054_), .B(_3053_), .C(_3055_), .Y(_3056_) );
OAI21X1 OAI21X1_938 ( .A(_3037__bF_buf1), .B(_4236__bF_buf1), .C(_4262__bF_buf4), .Y(_3057_) );
OAI22X1 OAI22X1_34 ( .A(micro_hash_ucr_a_2_bF_buf4_), .B(_4262__bF_buf2), .C(_3056_), .D(_3057_), .Y(_3058_) );
NAND2X1 NAND2X1_400 ( .A(_4234__bF_buf3), .B(_3058_), .Y(_3059_) );
NAND2X1 NAND2X1_401 ( .A(micro_hash_ucr_pipe23), .B(_3037__bF_buf1), .Y(_3060_) );
NAND3X1 NAND3X1_113 ( .A(_4233__bF_buf1), .B(_3060_), .C(_3059_), .Y(_3061_) );
NAND3X1 NAND3X1_114 ( .A(_389__bF_buf1), .B(_3031_), .C(_3061_), .Y(_3062_) );
NAND2X1 NAND2X1_402 ( .A(micro_hash_ucr_pipe25_bF_buf0), .B(_3037__bF_buf1), .Y(_3063_) );
NAND3X1 NAND3X1_115 ( .A(_4230__bF_buf1), .B(_3063_), .C(_3062_), .Y(_3064_) );
AOI21X1 AOI21X1_464 ( .A(micro_hash_ucr_a_2_bF_buf3_), .B(micro_hash_ucr_pipe26_bF_buf2), .C(micro_hash_ucr_pipe27_bF_buf3), .Y(_3065_) );
OAI21X1 OAI21X1_939 ( .A(_3038_), .B(_4229_), .C(_220__bF_buf2), .Y(_3066_) );
AOI21X1 AOI21X1_465 ( .A(_3065_), .B(_3064_), .C(_3066_), .Y(_3067_) );
NOR2X1 NOR2X1_678 ( .A(_3032_), .B(_220__bF_buf2), .Y(_3068_) );
OAI21X1 OAI21X1_940 ( .A(_3067_), .B(_3068_), .C(_219_), .Y(_3069_) );
NAND2X1 NAND2X1_403 ( .A(micro_hash_ucr_pipe29), .B(_3038_), .Y(_3070_) );
AOI21X1 AOI21X1_466 ( .A(_3070_), .B(_3069_), .C(micro_hash_ucr_pipe30_bF_buf3), .Y(_3071_) );
OAI21X1 OAI21X1_941 ( .A(_3032_), .B(_4228__bF_buf0), .C(_317__bF_buf2), .Y(_3072_) );
AOI21X1 AOI21X1_467 ( .A(micro_hash_ucr_pipe31_bF_buf2), .B(_3037__bF_buf1), .C(micro_hash_ucr_pipe32_bF_buf1), .Y(_3073_) );
OAI21X1 OAI21X1_942 ( .A(_3071_), .B(_3072_), .C(_3073_), .Y(_3074_) );
NAND2X1 NAND2X1_404 ( .A(micro_hash_ucr_a_2_bF_buf2_), .B(micro_hash_ucr_pipe32_bF_buf0), .Y(_3075_) );
NAND3X1 NAND3X1_116 ( .A(_318_), .B(_3075_), .C(_3074_), .Y(_3076_) );
NAND2X1 NAND2X1_405 ( .A(micro_hash_ucr_pipe33_bF_buf0), .B(_3037__bF_buf3), .Y(_3077_) );
NAND3X1 NAND3X1_117 ( .A(_4225__bF_buf4), .B(_3077_), .C(_3076_), .Y(_3078_) );
AOI21X1 AOI21X1_468 ( .A(micro_hash_ucr_a_2_bF_buf1_), .B(micro_hash_ucr_pipe34_bF_buf3), .C(micro_hash_ucr_pipe35), .Y(_3079_) );
OAI21X1 OAI21X1_943 ( .A(_3038_), .B(_230__bF_buf2), .C(_4224__bF_buf2), .Y(_3080_) );
AOI21X1 AOI21X1_469 ( .A(_3079_), .B(_3078_), .C(_3080_), .Y(_3081_) );
NOR2X1 NOR2X1_679 ( .A(_3032_), .B(_4224__bF_buf2), .Y(_3082_) );
OAI21X1 OAI21X1_944 ( .A(_3081_), .B(_3082_), .C(_2815_), .Y(_3083_) );
AOI21X1 AOI21X1_470 ( .A(micro_hash_ucr_pipe37_bF_buf1), .B(_3038_), .C(micro_hash_ucr_pipe38_bF_buf2), .Y(_3084_) );
OAI21X1 OAI21X1_945 ( .A(_701__bF_buf1), .B(micro_hash_ucr_a_2_bF_buf0_), .C(_2813__bF_buf0), .Y(_3085_) );
AOI21X1 AOI21X1_471 ( .A(_3084_), .B(_3083_), .C(_3085_), .Y(_3086_) );
OAI21X1 OAI21X1_946 ( .A(_3037__bF_buf3), .B(_2813__bF_buf0), .C(_296__bF_buf3), .Y(_3087_) );
NAND2X1 NAND2X1_406 ( .A(micro_hash_ucr_pipe40_bF_buf1), .B(_3032_), .Y(_3088_) );
OAI21X1 OAI21X1_947 ( .A(_3086_), .B(_3087_), .C(_3088_), .Y(_3089_) );
NAND2X1 NAND2X1_407 ( .A(_2814_), .B(_3089_), .Y(_3090_) );
NAND2X1 NAND2X1_408 ( .A(micro_hash_ucr_pipe41_bF_buf3), .B(_3037__bF_buf3), .Y(_3091_) );
NAND3X1 NAND3X1_118 ( .A(_4220__bF_buf2), .B(_3091_), .C(_3090_), .Y(_3092_) );
NAND3X1 NAND3X1_119 ( .A(_242__bF_buf0), .B(_3030_), .C(_3092_), .Y(_3093_) );
NAND2X1 NAND2X1_409 ( .A(micro_hash_ucr_pipe43), .B(_3037__bF_buf3), .Y(_3094_) );
NAND3X1 NAND3X1_120 ( .A(_4219__bF_buf3), .B(_3094_), .C(_3093_), .Y(_3095_) );
NAND3X1 NAND3X1_121 ( .A(_336_), .B(_3029_), .C(_3095_), .Y(_3096_) );
NAND2X1 NAND2X1_410 ( .A(micro_hash_ucr_pipe45), .B(_3037__bF_buf3), .Y(_3097_) );
NAND3X1 NAND3X1_122 ( .A(_4218__bF_buf2), .B(_3097_), .C(_3096_), .Y(_3098_) );
NAND3X1 NAND3X1_123 ( .A(_249__bF_buf3), .B(_3028_), .C(_3098_), .Y(_3099_) );
NAND2X1 NAND2X1_411 ( .A(micro_hash_ucr_pipe47), .B(_3037__bF_buf2), .Y(_3100_) );
NAND3X1 NAND3X1_124 ( .A(_4217__bF_buf3), .B(_3100_), .C(_3099_), .Y(_3101_) );
AOI21X1 AOI21X1_472 ( .A(_3027_), .B(_3101_), .C(micro_hash_ucr_pipe49_bF_buf1), .Y(_3102_) );
OAI21X1 OAI21X1_948 ( .A(_3037__bF_buf2), .B(_304_), .C(_4215__bF_buf1), .Y(_3103_) );
AOI21X1 AOI21X1_473 ( .A(micro_hash_ucr_pipe50_bF_buf3), .B(_3032_), .C(micro_hash_ucr_pipe51), .Y(_3104_) );
OAI21X1 OAI21X1_949 ( .A(_3102_), .B(_3103_), .C(_3104_), .Y(_3105_) );
AOI21X1 AOI21X1_474 ( .A(micro_hash_ucr_pipe51), .B(_3038_), .C(micro_hash_ucr_pipe52_bF_buf2), .Y(_3106_) );
NOR2X1 NOR2X1_680 ( .A(micro_hash_ucr_a_2_bF_buf4_), .B(_4214__bF_buf0), .Y(_3107_) );
AOI21X1 AOI21X1_475 ( .A(_3106_), .B(_3105_), .C(_3107_), .Y(_3108_) );
AOI21X1 AOI21X1_476 ( .A(micro_hash_ucr_pipe53_bF_buf3), .B(_3037__bF_buf2), .C(micro_hash_ucr_pipe54_bF_buf3), .Y(_3109_) );
OAI21X1 OAI21X1_950 ( .A(_3108_), .B(micro_hash_ucr_pipe53_bF_buf3), .C(_3109_), .Y(_3110_) );
NAND2X1 NAND2X1_412 ( .A(micro_hash_ucr_pipe54_bF_buf3), .B(micro_hash_ucr_a_2_bF_buf3_), .Y(_3111_) );
NAND3X1 NAND3X1_125 ( .A(_2811__bF_buf1), .B(_3111_), .C(_3110_), .Y(_3112_) );
NAND2X1 NAND2X1_413 ( .A(micro_hash_ucr_pipe55), .B(_3037__bF_buf2), .Y(_3113_) );
NAND3X1 NAND3X1_126 ( .A(_832__bF_buf0), .B(_3113_), .C(_3112_), .Y(_3114_) );
NAND3X1 NAND3X1_127 ( .A(_4212_), .B(_3026_), .C(_3114_), .Y(_3115_) );
NAND2X1 NAND2X1_414 ( .A(micro_hash_ucr_pipe57_bF_buf1), .B(_3037__bF_buf0), .Y(_3116_) );
NAND3X1 NAND3X1_128 ( .A(_4211__bF_buf1), .B(_3116_), .C(_3115_), .Y(_3117_) );
NAND3X1 NAND3X1_129 ( .A(_269_), .B(_3025_), .C(_3117_), .Y(_3118_) );
NAND2X1 NAND2X1_415 ( .A(micro_hash_ucr_pipe59), .B(_3037__bF_buf0), .Y(_3119_) );
NAND3X1 NAND3X1_130 ( .A(_4210__bF_buf1), .B(_3119_), .C(_3118_), .Y(_3120_) );
AOI21X1 AOI21X1_477 ( .A(micro_hash_ucr_pipe60_bF_buf1), .B(micro_hash_ucr_a_2_bF_buf2_), .C(micro_hash_ucr_pipe61_bF_buf2), .Y(_3121_) );
NOR2X1 NOR2X1_681 ( .A(_4208_), .B(_3038_), .Y(_3122_) );
AOI21X1 AOI21X1_478 ( .A(_3121_), .B(_3120_), .C(_3122_), .Y(_3123_) );
AOI21X1 AOI21X1_479 ( .A(micro_hash_ucr_pipe62_bF_buf0), .B(_3032_), .C(micro_hash_ucr_pipe63_bF_buf1), .Y(_3124_) );
OAI21X1 OAI21X1_951 ( .A(_3123_), .B(micro_hash_ucr_pipe62_bF_buf0), .C(_3124_), .Y(_3125_) );
AOI21X1 AOI21X1_480 ( .A(micro_hash_ucr_pipe63_bF_buf0), .B(_3038_), .C(micro_hash_ucr_pipe64_bF_buf4), .Y(_3126_) );
NOR2X1 NOR2X1_682 ( .A(micro_hash_ucr_a_2_bF_buf1_), .B(_278__bF_buf0), .Y(_3127_) );
AOI21X1 AOI21X1_481 ( .A(_3126_), .B(_3125_), .C(_3127_), .Y(_3128_) );
NAND2X1 NAND2X1_416 ( .A(micro_hash_ucr_pipe65_bF_buf2), .B(_3037__bF_buf0), .Y(_3129_) );
OAI21X1 OAI21X1_952 ( .A(_3128_), .B(micro_hash_ucr_pipe65_bF_buf2), .C(_3129_), .Y(_3130_) );
OAI21X1 OAI21X1_953 ( .A(_3130_), .B(micro_hash_ucr_pipe66_bF_buf4), .C(_3024_), .Y(_3131_) );
OAI21X1 OAI21X1_954 ( .A(_3037__bF_buf0), .B(_4201__bF_buf3), .C(_4199__bF_buf0), .Y(_3132_) );
AOI21X1 AOI21X1_482 ( .A(_4201__bF_buf3), .B(_3131_), .C(_3132_), .Y(_3133_) );
OAI21X1 OAI21X1_955 ( .A(_4199__bF_buf3), .B(micro_hash_ucr_a_2_bF_buf0_), .C(_344_), .Y(_3134_) );
NAND2X1 NAND2X1_417 ( .A(_3038_), .B(_198_), .Y(_3135_) );
OAI21X1 OAI21X1_956 ( .A(_3133_), .B(_3134_), .C(_3135_), .Y(_126__2_) );
NOR2X1 NOR2X1_683 ( .A(micro_hash_ucr_c_3_bF_buf2_), .B(micro_hash_ucr_b_3_bF_buf3_), .Y(_3136_) );
NOR2X1 NOR2X1_684 ( .A(_4200_), .B(_2468_), .Y(_3137_) );
NOR2X1 NOR2X1_685 ( .A(_3136_), .B(_3137_), .Y(_3138_) );
NAND2X1 NAND2X1_418 ( .A(_3138__bF_buf3), .B(_198_), .Y(_3139_) );
NAND2X1 NAND2X1_419 ( .A(micro_hash_ucr_pipe66_bF_buf4), .B(micro_hash_ucr_a_3_bF_buf3_), .Y(_3140_) );
NAND2X1 NAND2X1_420 ( .A(micro_hash_ucr_pipe64_bF_buf1), .B(micro_hash_ucr_a_3_bF_buf2_), .Y(_3141_) );
NAND2X1 NAND2X1_421 ( .A(micro_hash_ucr_pipe62_bF_buf2), .B(micro_hash_ucr_a_3_bF_buf1_), .Y(_3142_) );
NAND2X1 NAND2X1_422 ( .A(micro_hash_ucr_pipe60_bF_buf4), .B(micro_hash_ucr_a_3_bF_buf0_), .Y(_3143_) );
NAND2X1 NAND2X1_423 ( .A(micro_hash_ucr_pipe58_bF_buf0), .B(micro_hash_ucr_a_3_bF_buf3_), .Y(_3144_) );
NAND2X1 NAND2X1_424 ( .A(micro_hash_ucr_pipe52_bF_buf2), .B(_2531_), .Y(_3145_) );
NAND2X1 NAND2X1_425 ( .A(micro_hash_ucr_pipe50_bF_buf3), .B(_2531_), .Y(_3146_) );
NAND2X1 NAND2X1_426 ( .A(micro_hash_ucr_pipe48_bF_buf2), .B(_2531_), .Y(_3147_) );
NAND2X1 NAND2X1_427 ( .A(micro_hash_ucr_pipe22_bF_buf3), .B(_2531_), .Y(_3148_) );
NAND2X1 NAND2X1_428 ( .A(micro_hash_ucr_pipe20_bF_buf0), .B(_2531_), .Y(_3149_) );
NAND2X1 NAND2X1_429 ( .A(micro_hash_ucr_a_3_bF_buf2_), .B(micro_hash_ucr_pipe14), .Y(_3150_) );
NAND2X1 NAND2X1_430 ( .A(micro_hash_ucr_a_3_bF_buf1_), .B(micro_hash_ucr_pipe12_bF_buf0), .Y(_3151_) );
INVX1 INVX1_333 ( .A(_4244_), .Y(_3152_) );
NAND3X1 NAND3X1_131 ( .A(_2532_), .B(_4253_), .C(_4267_), .Y(_3153_) );
OAI21X1 OAI21X1_957 ( .A(_4272_), .B(_3138__bF_buf3), .C(_3153_), .Y(_3154_) );
AOI22X1 AOI22X1_21 ( .A(_2531_), .B(_4257_), .C(_3154_), .D(_3152_), .Y(_3155_) );
AOI21X1 AOI21X1_483 ( .A(micro_hash_ucr_pipe11), .B(_3138__bF_buf3), .C(_3155_), .Y(_3156_) );
OAI21X1 OAI21X1_958 ( .A(_3156_), .B(micro_hash_ucr_pipe12_bF_buf0), .C(_3151_), .Y(_3157_) );
OAI21X1 OAI21X1_959 ( .A(_3137_), .B(_3136_), .C(micro_hash_ucr_pipe13), .Y(_3158_) );
OAI21X1 OAI21X1_960 ( .A(_3157_), .B(micro_hash_ucr_pipe13), .C(_3158_), .Y(_3159_) );
OAI21X1 OAI21X1_961 ( .A(_3159_), .B(micro_hash_ucr_pipe14), .C(_3150_), .Y(_3160_) );
INVX4 INVX4_48 ( .A(_3138__bF_buf2), .Y(_3161_) );
OAI21X1 OAI21X1_962 ( .A(_3161_), .B(_4240_), .C(_4239__bF_buf1), .Y(_3162_) );
AOI21X1 AOI21X1_484 ( .A(_4240_), .B(_3160_), .C(_3162_), .Y(_3163_) );
OAI21X1 OAI21X1_963 ( .A(_4239__bF_buf1), .B(micro_hash_ucr_a_3_bF_buf0_), .C(_4238__bF_buf2), .Y(_3164_) );
AOI21X1 AOI21X1_485 ( .A(micro_hash_ucr_pipe17), .B(_3138__bF_buf3), .C(micro_hash_ucr_pipe18_bF_buf4), .Y(_3165_) );
OAI21X1 OAI21X1_964 ( .A(_3163_), .B(_3164_), .C(_3165_), .Y(_3166_) );
NAND2X1 NAND2X1_431 ( .A(micro_hash_ucr_pipe18_bF_buf1), .B(_2531_), .Y(_3167_) );
AOI21X1 AOI21X1_486 ( .A(_3167_), .B(_3166_), .C(micro_hash_ucr_pipe19), .Y(_3168_) );
NOR2X1 NOR2X1_686 ( .A(_2816_), .B(_3138__bF_buf3), .Y(_3169_) );
OAI21X1 OAI21X1_965 ( .A(_3168_), .B(_3169_), .C(_4237__bF_buf0), .Y(_3170_) );
AOI21X1 AOI21X1_487 ( .A(_3149_), .B(_3170_), .C(micro_hash_ucr_pipe21), .Y(_3171_) );
NOR2X1 NOR2X1_687 ( .A(_4236__bF_buf3), .B(_3138__bF_buf2), .Y(_3172_) );
OAI21X1 OAI21X1_966 ( .A(_3171_), .B(_3172_), .C(_4262__bF_buf2), .Y(_3173_) );
NAND3X1 NAND3X1_132 ( .A(_4234__bF_buf3), .B(_3148_), .C(_3173_), .Y(_3174_) );
AOI21X1 AOI21X1_488 ( .A(micro_hash_ucr_pipe23), .B(_3138__bF_buf2), .C(micro_hash_ucr_pipe24_bF_buf3), .Y(_3175_) );
OAI21X1 OAI21X1_967 ( .A(_4233__bF_buf2), .B(micro_hash_ucr_a_3_bF_buf3_), .C(_389__bF_buf2), .Y(_3176_) );
AOI21X1 AOI21X1_489 ( .A(_3175_), .B(_3174_), .C(_3176_), .Y(_3177_) );
OAI21X1 OAI21X1_968 ( .A(_3161_), .B(_389__bF_buf2), .C(_4230__bF_buf0), .Y(_3178_) );
OAI22X1 OAI22X1_35 ( .A(micro_hash_ucr_a_3_bF_buf2_), .B(_4230__bF_buf0), .C(_3177_), .D(_3178_), .Y(_3179_) );
AOI21X1 AOI21X1_490 ( .A(micro_hash_ucr_pipe27_bF_buf0), .B(_3138__bF_buf2), .C(micro_hash_ucr_pipe28_bF_buf0), .Y(_3180_) );
OAI21X1 OAI21X1_969 ( .A(_3179_), .B(micro_hash_ucr_pipe27_bF_buf0), .C(_3180_), .Y(_3181_) );
AOI21X1 AOI21X1_491 ( .A(micro_hash_ucr_pipe28_bF_buf0), .B(_2531_), .C(micro_hash_ucr_pipe29), .Y(_3182_) );
OAI21X1 OAI21X1_970 ( .A(_3161_), .B(_219_), .C(_4228__bF_buf2), .Y(_3183_) );
AOI21X1 AOI21X1_492 ( .A(_3182_), .B(_3181_), .C(_3183_), .Y(_3184_) );
NOR2X1 NOR2X1_688 ( .A(micro_hash_ucr_a_3_bF_buf1_), .B(_4228__bF_buf2), .Y(_3185_) );
OAI21X1 OAI21X1_971 ( .A(_3184_), .B(_3185_), .C(_317__bF_buf1), .Y(_3186_) );
OAI21X1 OAI21X1_972 ( .A(_3137_), .B(_3136_), .C(micro_hash_ucr_pipe31_bF_buf3), .Y(_3187_) );
NAND3X1 NAND3X1_133 ( .A(_4226__bF_buf3), .B(_3187_), .C(_3186_), .Y(_3188_) );
AOI21X1 AOI21X1_493 ( .A(micro_hash_ucr_a_3_bF_buf0_), .B(micro_hash_ucr_pipe32_bF_buf2), .C(micro_hash_ucr_pipe33_bF_buf3), .Y(_3189_) );
OAI21X1 OAI21X1_973 ( .A(_3138__bF_buf0), .B(_318_), .C(_4225__bF_buf3), .Y(_3190_) );
AOI21X1 AOI21X1_494 ( .A(_3189_), .B(_3188_), .C(_3190_), .Y(_3191_) );
NOR2X1 NOR2X1_689 ( .A(_2531_), .B(_4225__bF_buf3), .Y(_3192_) );
OAI21X1 OAI21X1_974 ( .A(_3191_), .B(_3192_), .C(_230__bF_buf3), .Y(_3193_) );
AOI21X1 AOI21X1_495 ( .A(micro_hash_ucr_pipe35), .B(_3138__bF_buf0), .C(micro_hash_ucr_pipe36_bF_buf2), .Y(_3194_) );
OAI21X1 OAI21X1_975 ( .A(_4224__bF_buf0), .B(micro_hash_ucr_a_3_bF_buf3_), .C(_2815_), .Y(_3195_) );
AOI21X1 AOI21X1_496 ( .A(_3194_), .B(_3193_), .C(_3195_), .Y(_3196_) );
OAI21X1 OAI21X1_976 ( .A(_3161_), .B(_2815_), .C(_701__bF_buf3), .Y(_3197_) );
OAI22X1 OAI22X1_36 ( .A(micro_hash_ucr_a_3_bF_buf2_), .B(_701__bF_buf3), .C(_3196_), .D(_3197_), .Y(_3198_) );
NOR2X1 NOR2X1_690 ( .A(micro_hash_ucr_pipe39), .B(_3198_), .Y(_3199_) );
OAI21X1 OAI21X1_977 ( .A(_3161_), .B(_2813__bF_buf3), .C(_296__bF_buf0), .Y(_3200_) );
AOI21X1 AOI21X1_497 ( .A(micro_hash_ucr_pipe40_bF_buf0), .B(_2531_), .C(micro_hash_ucr_pipe41_bF_buf2), .Y(_3201_) );
OAI21X1 OAI21X1_978 ( .A(_3199_), .B(_3200_), .C(_3201_), .Y(_3202_) );
AOI21X1 AOI21X1_498 ( .A(micro_hash_ucr_pipe41_bF_buf2), .B(_3138__bF_buf0), .C(micro_hash_ucr_pipe42_bF_buf4), .Y(_3203_) );
AOI22X1 AOI22X1_22 ( .A(micro_hash_ucr_pipe42_bF_buf4), .B(_2531_), .C(_3202_), .D(_3203_), .Y(_3204_) );
OAI21X1 OAI21X1_979 ( .A(_3161_), .B(_242__bF_buf1), .C(_4219__bF_buf0), .Y(_3205_) );
AOI21X1 AOI21X1_499 ( .A(_242__bF_buf1), .B(_3204_), .C(_3205_), .Y(_3206_) );
OAI21X1 OAI21X1_980 ( .A(_4219__bF_buf0), .B(micro_hash_ucr_a_3_bF_buf1_), .C(_336_), .Y(_3207_) );
AOI21X1 AOI21X1_500 ( .A(micro_hash_ucr_pipe45), .B(_3138__bF_buf0), .C(micro_hash_ucr_pipe46_bF_buf1), .Y(_3208_) );
OAI21X1 OAI21X1_981 ( .A(_3206_), .B(_3207_), .C(_3208_), .Y(_3209_) );
NAND2X1 NAND2X1_432 ( .A(micro_hash_ucr_pipe46_bF_buf4), .B(_2531_), .Y(_3210_) );
AOI21X1 AOI21X1_501 ( .A(_3210_), .B(_3209_), .C(micro_hash_ucr_pipe47), .Y(_3211_) );
NOR2X1 NOR2X1_691 ( .A(_249__bF_buf3), .B(_3138__bF_buf1), .Y(_3212_) );
OAI21X1 OAI21X1_982 ( .A(_3211_), .B(_3212_), .C(_4217__bF_buf3), .Y(_3213_) );
NAND3X1 NAND3X1_134 ( .A(_304_), .B(_3147_), .C(_3213_), .Y(_3214_) );
NAND2X1 NAND2X1_433 ( .A(micro_hash_ucr_pipe49_bF_buf2), .B(_3138__bF_buf1), .Y(_3215_) );
NAND3X1 NAND3X1_135 ( .A(_4215__bF_buf2), .B(_3215_), .C(_3214_), .Y(_3216_) );
NAND3X1 NAND3X1_136 ( .A(_255__bF_buf0), .B(_3146_), .C(_3216_), .Y(_3217_) );
NAND2X1 NAND2X1_434 ( .A(micro_hash_ucr_pipe51), .B(_3138__bF_buf1), .Y(_3218_) );
NAND3X1 NAND3X1_137 ( .A(_4214__bF_buf0), .B(_3218_), .C(_3217_), .Y(_3219_) );
NAND3X1 NAND3X1_138 ( .A(_2812_), .B(_3145_), .C(_3219_), .Y(_3220_) );
AOI21X1 AOI21X1_502 ( .A(micro_hash_ucr_pipe53_bF_buf3), .B(_3138__bF_buf1), .C(micro_hash_ucr_pipe54_bF_buf3), .Y(_3221_) );
OAI21X1 OAI21X1_983 ( .A(_742__bF_buf0), .B(micro_hash_ucr_a_3_bF_buf0_), .C(_2811__bF_buf0), .Y(_3222_) );
AOI21X1 AOI21X1_503 ( .A(_3221_), .B(_3220_), .C(_3222_), .Y(_3223_) );
OAI21X1 OAI21X1_984 ( .A(_3161_), .B(_2811__bF_buf0), .C(_832__bF_buf2), .Y(_3224_) );
NAND2X1 NAND2X1_435 ( .A(micro_hash_ucr_pipe56_bF_buf2), .B(_2531_), .Y(_3225_) );
OAI21X1 OAI21X1_985 ( .A(_3223_), .B(_3224_), .C(_3225_), .Y(_3226_) );
NAND2X1 NAND2X1_436 ( .A(_4212_), .B(_3226_), .Y(_3227_) );
OAI21X1 OAI21X1_986 ( .A(_3137_), .B(_3136_), .C(micro_hash_ucr_pipe57_bF_buf1), .Y(_3228_) );
NAND3X1 NAND3X1_139 ( .A(_4211__bF_buf0), .B(_3228_), .C(_3227_), .Y(_3229_) );
NAND3X1 NAND3X1_140 ( .A(_269_), .B(_3144_), .C(_3229_), .Y(_3230_) );
OAI21X1 OAI21X1_987 ( .A(_3137_), .B(_3136_), .C(micro_hash_ucr_pipe59), .Y(_3231_) );
NAND3X1 NAND3X1_141 ( .A(_4210__bF_buf1), .B(_3231_), .C(_3230_), .Y(_3232_) );
NAND3X1 NAND3X1_142 ( .A(_4208_), .B(_3143_), .C(_3232_), .Y(_3233_) );
OAI21X1 OAI21X1_988 ( .A(_3137_), .B(_3136_), .C(micro_hash_ucr_pipe61_bF_buf3), .Y(_3234_) );
NAND3X1 NAND3X1_143 ( .A(_4207__bF_buf4), .B(_3234_), .C(_3233_), .Y(_3235_) );
NAND3X1 NAND3X1_144 ( .A(_4204_), .B(_3142_), .C(_3235_), .Y(_3236_) );
OAI21X1 OAI21X1_989 ( .A(_3137_), .B(_3136_), .C(micro_hash_ucr_pipe63_bF_buf3), .Y(_3237_) );
NAND3X1 NAND3X1_145 ( .A(_278__bF_buf0), .B(_3237_), .C(_3236_), .Y(_3238_) );
NAND3X1 NAND3X1_146 ( .A(_279_), .B(_3141_), .C(_3238_), .Y(_3239_) );
OAI21X1 OAI21X1_990 ( .A(_3137_), .B(_3136_), .C(micro_hash_ucr_pipe65_bF_buf1), .Y(_3240_) );
NAND3X1 NAND3X1_147 ( .A(_1078__bF_buf1), .B(_3240_), .C(_3239_), .Y(_3241_) );
NAND2X1 NAND2X1_437 ( .A(_3140_), .B(_3241_), .Y(_3242_) );
OAI21X1 OAI21X1_991 ( .A(_3161_), .B(_4201__bF_buf1), .C(_4199__bF_buf3), .Y(_3243_) );
AOI21X1 AOI21X1_504 ( .A(_4201__bF_buf1), .B(_3242_), .C(_3243_), .Y(_3244_) );
OAI21X1 OAI21X1_992 ( .A(_4199__bF_buf3), .B(micro_hash_ucr_a_3_bF_buf3_), .C(_344_), .Y(_3245_) );
OAI21X1 OAI21X1_993 ( .A(_3244_), .B(_3245_), .C(_3139_), .Y(_126__3_) );
XNOR2X1 XNOR2X1_212 ( .A(micro_hash_ucr_b_4_), .B(micro_hash_ucr_c_4_), .Y(_3246_) );
INVX8 INVX8_87 ( .A(_3246__bF_buf2), .Y(_3247_) );
NAND2X1 NAND2X1_438 ( .A(_3247_), .B(_198_), .Y(_3248_) );
NAND2X1 NAND2X1_439 ( .A(micro_hash_ucr_pipe66_bF_buf4), .B(micro_hash_ucr_a_4_bF_buf3_), .Y(_3249_) );
NAND2X1 NAND2X1_440 ( .A(micro_hash_ucr_pipe64_bF_buf4), .B(micro_hash_ucr_a_4_bF_buf2_), .Y(_3250_) );
NAND2X1 NAND2X1_441 ( .A(micro_hash_ucr_pipe56_bF_buf2), .B(micro_hash_ucr_a_4_bF_buf1_), .Y(_3251_) );
NAND2X1 NAND2X1_442 ( .A(micro_hash_ucr_pipe54_bF_buf3), .B(micro_hash_ucr_a_4_bF_buf0_), .Y(_3252_) );
NAND2X1 NAND2X1_443 ( .A(micro_hash_ucr_pipe52_bF_buf2), .B(micro_hash_ucr_a_4_bF_buf3_), .Y(_3253_) );
NAND2X1 NAND2X1_444 ( .A(micro_hash_ucr_pipe36_bF_buf3), .B(_2546_), .Y(_3254_) );
NAND2X1 NAND2X1_445 ( .A(micro_hash_ucr_pipe34_bF_buf1), .B(_2546_), .Y(_3255_) );
NAND2X1 NAND2X1_446 ( .A(micro_hash_ucr_pipe24_bF_buf3), .B(_2546_), .Y(_3256_) );
NAND2X1 NAND2X1_447 ( .A(micro_hash_ucr_pipe22_bF_buf3), .B(_2546_), .Y(_3257_) );
NAND2X1 NAND2X1_448 ( .A(micro_hash_ucr_a_4_bF_buf2_), .B(micro_hash_ucr_pipe16), .Y(_3258_) );
NAND2X1 NAND2X1_449 ( .A(micro_hash_ucr_a_4_bF_buf1_), .B(micro_hash_ucr_pipe14), .Y(_3259_) );
NOR2X1 NOR2X1_692 ( .A(micro_hash_ucr_a_4_bF_buf0_), .B(_2923_), .Y(_3260_) );
OAI21X1 OAI21X1_994 ( .A(_4256_), .B(micro_hash_ucr_pipe11), .C(_3246__bF_buf0), .Y(_3261_) );
NAND3X1 NAND3X1_148 ( .A(_4255_), .B(_2543_), .C(_2823_), .Y(_3262_) );
AOI21X1 AOI21X1_505 ( .A(_3261_), .B(_3262_), .C(_4244_), .Y(_3263_) );
OAI22X1 OAI22X1_37 ( .A(_4277_), .B(_3246__bF_buf0), .C(_3263_), .D(_3260_), .Y(_3264_) );
NAND2X1 NAND2X1_450 ( .A(micro_hash_ucr_pipe12_bF_buf3), .B(_2546_), .Y(_3265_) );
OAI21X1 OAI21X1_995 ( .A(_3264_), .B(micro_hash_ucr_pipe12_bF_buf3), .C(_3265_), .Y(_3266_) );
NOR2X1 NOR2X1_693 ( .A(micro_hash_ucr_pipe13), .B(_3266_), .Y(_3267_) );
NOR2X1 NOR2X1_694 ( .A(_4242_), .B(_3246__bF_buf0), .Y(_3268_) );
OAI21X1 OAI21X1_996 ( .A(_3267_), .B(_3268_), .C(_4241__bF_buf3), .Y(_3269_) );
NAND3X1 NAND3X1_149 ( .A(_4240_), .B(_3259_), .C(_3269_), .Y(_3270_) );
NAND2X1 NAND2X1_451 ( .A(micro_hash_ucr_pipe15), .B(_3246__bF_buf0), .Y(_3271_) );
NAND3X1 NAND3X1_150 ( .A(_4239__bF_buf3), .B(_3271_), .C(_3270_), .Y(_3272_) );
NAND3X1 NAND3X1_151 ( .A(_4238__bF_buf2), .B(_3258_), .C(_3272_), .Y(_3273_) );
NAND2X1 NAND2X1_452 ( .A(micro_hash_ucr_pipe17), .B(_3246__bF_buf2), .Y(_3274_) );
NAND3X1 NAND3X1_152 ( .A(_624__bF_buf1), .B(_3274_), .C(_3273_), .Y(_3275_) );
AOI21X1 AOI21X1_506 ( .A(micro_hash_ucr_a_4_bF_buf3_), .B(micro_hash_ucr_pipe18_bF_buf1), .C(micro_hash_ucr_pipe19), .Y(_3276_) );
OAI21X1 OAI21X1_997 ( .A(_3247_), .B(_2816_), .C(_4237__bF_buf0), .Y(_3277_) );
AOI21X1 AOI21X1_507 ( .A(_3276_), .B(_3275_), .C(_3277_), .Y(_3278_) );
NOR2X1 NOR2X1_695 ( .A(_2546_), .B(_4237__bF_buf2), .Y(_3279_) );
OAI21X1 OAI21X1_998 ( .A(_3278_), .B(_3279_), .C(_4236__bF_buf2), .Y(_3280_) );
NAND2X1 NAND2X1_453 ( .A(micro_hash_ucr_pipe21), .B(_3247_), .Y(_3281_) );
NAND3X1 NAND3X1_153 ( .A(_4262__bF_buf4), .B(_3281_), .C(_3280_), .Y(_3282_) );
NAND3X1 NAND3X1_154 ( .A(_4234__bF_buf3), .B(_3257_), .C(_3282_), .Y(_3283_) );
NAND2X1 NAND2X1_454 ( .A(micro_hash_ucr_pipe23), .B(_3247_), .Y(_3284_) );
NAND3X1 NAND3X1_155 ( .A(_4233__bF_buf4), .B(_3284_), .C(_3283_), .Y(_3285_) );
NAND3X1 NAND3X1_156 ( .A(_389__bF_buf1), .B(_3256_), .C(_3285_), .Y(_3286_) );
AOI21X1 AOI21X1_508 ( .A(micro_hash_ucr_pipe25_bF_buf0), .B(_3247_), .C(micro_hash_ucr_pipe26_bF_buf1), .Y(_3287_) );
OAI21X1 OAI21X1_999 ( .A(_4230__bF_buf1), .B(micro_hash_ucr_a_4_bF_buf2_), .C(_4229_), .Y(_3288_) );
AOI21X1 AOI21X1_509 ( .A(_3287_), .B(_3286_), .C(_3288_), .Y(_3289_) );
OAI21X1 OAI21X1_1000 ( .A(_3246__bF_buf1), .B(_4229_), .C(_220__bF_buf2), .Y(_3290_) );
OAI22X1 OAI22X1_38 ( .A(micro_hash_ucr_a_4_bF_buf1_), .B(_220__bF_buf1), .C(_3289_), .D(_3290_), .Y(_3291_) );
NAND2X1 NAND2X1_455 ( .A(_219_), .B(_3291_), .Y(_3292_) );
NAND2X1 NAND2X1_456 ( .A(micro_hash_ucr_pipe29), .B(_3246__bF_buf1), .Y(_3293_) );
NAND3X1 NAND3X1_157 ( .A(_4228__bF_buf0), .B(_3293_), .C(_3292_), .Y(_3294_) );
AOI21X1 AOI21X1_510 ( .A(micro_hash_ucr_a_4_bF_buf0_), .B(micro_hash_ucr_pipe30_bF_buf3), .C(micro_hash_ucr_pipe31_bF_buf2), .Y(_3295_) );
OAI21X1 OAI21X1_1001 ( .A(_3247_), .B(_317__bF_buf2), .C(_4226__bF_buf1), .Y(_3296_) );
AOI21X1 AOI21X1_511 ( .A(_3295_), .B(_3294_), .C(_3296_), .Y(_3297_) );
NOR2X1 NOR2X1_696 ( .A(_2546_), .B(_4226__bF_buf2), .Y(_3298_) );
OAI21X1 OAI21X1_1002 ( .A(_3297_), .B(_3298_), .C(_318_), .Y(_3299_) );
NAND2X1 NAND2X1_457 ( .A(micro_hash_ucr_pipe33_bF_buf1), .B(_3247_), .Y(_3300_) );
NAND3X1 NAND3X1_158 ( .A(_4225__bF_buf4), .B(_3300_), .C(_3299_), .Y(_3301_) );
NAND3X1 NAND3X1_159 ( .A(_230__bF_buf1), .B(_3255_), .C(_3301_), .Y(_3302_) );
NAND2X1 NAND2X1_458 ( .A(micro_hash_ucr_pipe35), .B(_3247_), .Y(_3303_) );
NAND3X1 NAND3X1_160 ( .A(_4224__bF_buf3), .B(_3303_), .C(_3302_), .Y(_3304_) );
NAND3X1 NAND3X1_161 ( .A(_2815_), .B(_3254_), .C(_3304_), .Y(_3305_) );
AOI21X1 AOI21X1_512 ( .A(micro_hash_ucr_pipe37_bF_buf3), .B(_3247_), .C(micro_hash_ucr_pipe38_bF_buf0), .Y(_3306_) );
OAI21X1 OAI21X1_1003 ( .A(_701__bF_buf0), .B(micro_hash_ucr_a_4_bF_buf3_), .C(_2813__bF_buf0), .Y(_3307_) );
AOI21X1 AOI21X1_513 ( .A(_3306_), .B(_3305_), .C(_3307_), .Y(_3308_) );
OAI21X1 OAI21X1_1004 ( .A(_3246__bF_buf1), .B(_2813__bF_buf0), .C(_296__bF_buf1), .Y(_3309_) );
OAI22X1 OAI22X1_39 ( .A(_296__bF_buf3), .B(micro_hash_ucr_a_4_bF_buf2_), .C(_3308_), .D(_3309_), .Y(_3310_) );
AOI21X1 AOI21X1_514 ( .A(micro_hash_ucr_pipe41_bF_buf0), .B(_3247_), .C(micro_hash_ucr_pipe42_bF_buf1), .Y(_3311_) );
OAI21X1 OAI21X1_1005 ( .A(_3310_), .B(micro_hash_ucr_pipe41_bF_buf0), .C(_3311_), .Y(_3312_) );
AOI21X1 AOI21X1_515 ( .A(micro_hash_ucr_pipe42_bF_buf0), .B(_2546_), .C(micro_hash_ucr_pipe43), .Y(_3313_) );
AOI22X1 AOI22X1_23 ( .A(micro_hash_ucr_pipe43), .B(_3247_), .C(_3312_), .D(_3313_), .Y(_3314_) );
AOI21X1 AOI21X1_516 ( .A(micro_hash_ucr_pipe44_bF_buf3), .B(micro_hash_ucr_a_4_bF_buf1_), .C(micro_hash_ucr_pipe45), .Y(_3315_) );
OAI21X1 OAI21X1_1006 ( .A(_3314_), .B(micro_hash_ucr_pipe44_bF_buf3), .C(_3315_), .Y(_3316_) );
AOI21X1 AOI21X1_517 ( .A(micro_hash_ucr_pipe45), .B(_3246__bF_buf1), .C(micro_hash_ucr_pipe46_bF_buf3), .Y(_3317_) );
AOI22X1 AOI22X1_24 ( .A(micro_hash_ucr_pipe46_bF_buf3), .B(micro_hash_ucr_a_4_bF_buf0_), .C(_3316_), .D(_3317_), .Y(_3318_) );
AOI21X1 AOI21X1_518 ( .A(micro_hash_ucr_pipe47), .B(_3247_), .C(micro_hash_ucr_pipe48_bF_buf0), .Y(_3319_) );
OAI21X1 OAI21X1_1007 ( .A(_3318_), .B(micro_hash_ucr_pipe47), .C(_3319_), .Y(_3320_) );
AOI21X1 AOI21X1_519 ( .A(micro_hash_ucr_pipe48_bF_buf0), .B(_2546_), .C(micro_hash_ucr_pipe49_bF_buf1), .Y(_3321_) );
OAI21X1 OAI21X1_1008 ( .A(_3246__bF_buf3), .B(_304_), .C(_4215__bF_buf1), .Y(_3322_) );
AOI21X1 AOI21X1_520 ( .A(_3321_), .B(_3320_), .C(_3322_), .Y(_3323_) );
NOR2X1 NOR2X1_697 ( .A(micro_hash_ucr_a_4_bF_buf3_), .B(_4215__bF_buf1), .Y(_3324_) );
OAI21X1 OAI21X1_1009 ( .A(_3323_), .B(_3324_), .C(_255__bF_buf0), .Y(_3325_) );
NAND2X1 NAND2X1_459 ( .A(micro_hash_ucr_pipe51), .B(_3246__bF_buf3), .Y(_3326_) );
NAND3X1 NAND3X1_162 ( .A(_4214__bF_buf0), .B(_3326_), .C(_3325_), .Y(_3327_) );
NAND3X1 NAND3X1_163 ( .A(_2812_), .B(_3253_), .C(_3327_), .Y(_3328_) );
NAND2X1 NAND2X1_460 ( .A(micro_hash_ucr_pipe53_bF_buf3), .B(_3246__bF_buf3), .Y(_3329_) );
NAND3X1 NAND3X1_164 ( .A(_742__bF_buf0), .B(_3329_), .C(_3328_), .Y(_3330_) );
NAND3X1 NAND3X1_165 ( .A(_2811__bF_buf1), .B(_3252_), .C(_3330_), .Y(_3331_) );
NAND2X1 NAND2X1_461 ( .A(micro_hash_ucr_pipe55), .B(_3246__bF_buf3), .Y(_3332_) );
NAND3X1 NAND3X1_166 ( .A(_832__bF_buf0), .B(_3332_), .C(_3331_), .Y(_3333_) );
NAND3X1 NAND3X1_167 ( .A(_4212_), .B(_3251_), .C(_3333_), .Y(_3334_) );
NAND2X1 NAND2X1_462 ( .A(micro_hash_ucr_pipe57_bF_buf0), .B(_3246__bF_buf3), .Y(_3335_) );
NAND3X1 NAND3X1_168 ( .A(_4211__bF_buf1), .B(_3335_), .C(_3334_), .Y(_3336_) );
AOI21X1 AOI21X1_521 ( .A(micro_hash_ucr_pipe58_bF_buf0), .B(micro_hash_ucr_a_4_bF_buf2_), .C(micro_hash_ucr_pipe59), .Y(_3337_) );
NOR2X1 NOR2X1_698 ( .A(_269_), .B(_3247_), .Y(_3338_) );
AOI21X1 AOI21X1_522 ( .A(_3337_), .B(_3336_), .C(_3338_), .Y(_3339_) );
AOI21X1 AOI21X1_523 ( .A(micro_hash_ucr_pipe60_bF_buf1), .B(_2546_), .C(micro_hash_ucr_pipe61_bF_buf2), .Y(_3340_) );
OAI21X1 OAI21X1_1010 ( .A(_3339_), .B(micro_hash_ucr_pipe60_bF_buf1), .C(_3340_), .Y(_3341_) );
AOI21X1 AOI21X1_524 ( .A(micro_hash_ucr_pipe61_bF_buf2), .B(_3247_), .C(micro_hash_ucr_pipe62_bF_buf0), .Y(_3342_) );
NOR2X1 NOR2X1_699 ( .A(micro_hash_ucr_a_4_bF_buf1_), .B(_4207__bF_buf4), .Y(_3343_) );
AOI21X1 AOI21X1_525 ( .A(_3342_), .B(_3341_), .C(_3343_), .Y(_3344_) );
NAND2X1 NAND2X1_463 ( .A(micro_hash_ucr_pipe63_bF_buf0), .B(_3246__bF_buf2), .Y(_3345_) );
OAI21X1 OAI21X1_1011 ( .A(_3344_), .B(micro_hash_ucr_pipe63_bF_buf0), .C(_3345_), .Y(_3346_) );
OAI21X1 OAI21X1_1012 ( .A(_3346_), .B(micro_hash_ucr_pipe64_bF_buf4), .C(_3250_), .Y(_3347_) );
NAND2X1 NAND2X1_464 ( .A(micro_hash_ucr_pipe65_bF_buf2), .B(_3246__bF_buf2), .Y(_3348_) );
OAI21X1 OAI21X1_1013 ( .A(_3347_), .B(micro_hash_ucr_pipe65_bF_buf2), .C(_3348_), .Y(_3349_) );
OAI21X1 OAI21X1_1014 ( .A(_3349_), .B(micro_hash_ucr_pipe66_bF_buf4), .C(_3249_), .Y(_3350_) );
OAI21X1 OAI21X1_1015 ( .A(_3246__bF_buf2), .B(_4201__bF_buf3), .C(_4199__bF_buf3), .Y(_3351_) );
AOI21X1 AOI21X1_526 ( .A(_4201__bF_buf3), .B(_3350_), .C(_3351_), .Y(_3352_) );
OAI21X1 OAI21X1_1016 ( .A(_4199__bF_buf3), .B(micro_hash_ucr_a_4_bF_buf0_), .C(_344_), .Y(_3353_) );
OAI21X1 OAI21X1_1017 ( .A(_3352_), .B(_3353_), .C(_3248_), .Y(_126__4_) );
XNOR2X1 XNOR2X1_213 ( .A(micro_hash_ucr_b_5_bF_buf3_), .B(micro_hash_ucr_c_5_), .Y(_3354_) );
INVX8 INVX8_88 ( .A(_3354__bF_buf2), .Y(_3355_) );
NAND2X1 NAND2X1_465 ( .A(_3355_), .B(_198_), .Y(_3356_) );
NAND2X1 NAND2X1_466 ( .A(micro_hash_ucr_pipe62_bF_buf0), .B(micro_hash_ucr_a_5_bF_buf3_), .Y(_3357_) );
NAND2X1 NAND2X1_467 ( .A(micro_hash_ucr_pipe60_bF_buf1), .B(micro_hash_ucr_a_5_bF_buf2_), .Y(_3358_) );
NAND2X1 NAND2X1_468 ( .A(micro_hash_ucr_pipe58_bF_buf0), .B(micro_hash_ucr_a_5_bF_buf1_), .Y(_3359_) );
NAND2X1 NAND2X1_469 ( .A(micro_hash_ucr_pipe56_bF_buf2), .B(micro_hash_ucr_a_5_bF_buf0_), .Y(_3360_) );
NAND2X1 NAND2X1_470 ( .A(micro_hash_ucr_pipe50_bF_buf3), .B(_2551_), .Y(_3361_) );
NAND2X1 NAND2X1_471 ( .A(micro_hash_ucr_pipe44_bF_buf0), .B(micro_hash_ucr_a_5_bF_buf3_), .Y(_3362_) );
NAND2X1 NAND2X1_472 ( .A(micro_hash_ucr_pipe42_bF_buf0), .B(micro_hash_ucr_a_5_bF_buf2_), .Y(_3363_) );
NAND2X1 NAND2X1_473 ( .A(micro_hash_ucr_pipe40_bF_buf3), .B(micro_hash_ucr_a_5_bF_buf1_), .Y(_3364_) );
NAND2X1 NAND2X1_474 ( .A(micro_hash_ucr_pipe34_bF_buf1), .B(_2551_), .Y(_3365_) );
NAND2X1 NAND2X1_475 ( .A(micro_hash_ucr_a_5_bF_buf0_), .B(micro_hash_ucr_pipe28_bF_buf1), .Y(_3366_) );
NAND2X1 NAND2X1_476 ( .A(micro_hash_ucr_pipe18_bF_buf4), .B(_2551_), .Y(_3367_) );
NAND2X1 NAND2X1_477 ( .A(micro_hash_ucr_pipe16), .B(_2551_), .Y(_3368_) );
NAND2X1 NAND2X1_478 ( .A(micro_hash_ucr_pipe14), .B(_2551_), .Y(_3369_) );
NAND2X1 NAND2X1_479 ( .A(micro_hash_ucr_pipe12_bF_buf0), .B(_2551_), .Y(_3370_) );
NAND2X1 NAND2X1_480 ( .A(micro_hash_ucr_pipe11), .B(_3355_), .Y(_3371_) );
NAND2X1 NAND2X1_481 ( .A(_2551_), .B(_4257_), .Y(_3372_) );
NOR2X1 NOR2X1_700 ( .A(micro_hash_ucr_pipe9), .B(H_5_), .Y(_3373_) );
AOI22X1 AOI22X1_25 ( .A(_2823_), .B(_3373_), .C(_2925_), .D(_3354__bF_buf3), .Y(_3374_) );
OAI21X1 OAI21X1_1018 ( .A(_3374_), .B(_4244_), .C(_3372_), .Y(_3375_) );
NAND3X1 NAND3X1_169 ( .A(_4258_), .B(_3371_), .C(_3375_), .Y(_3376_) );
NAND3X1 NAND3X1_170 ( .A(_4242_), .B(_3370_), .C(_3376_), .Y(_3377_) );
NAND2X1 NAND2X1_482 ( .A(micro_hash_ucr_pipe13), .B(_3355_), .Y(_3378_) );
NAND3X1 NAND3X1_171 ( .A(_4241__bF_buf3), .B(_3378_), .C(_3377_), .Y(_3379_) );
NAND3X1 NAND3X1_172 ( .A(_4240_), .B(_3369_), .C(_3379_), .Y(_3380_) );
NAND2X1 NAND2X1_483 ( .A(micro_hash_ucr_pipe15), .B(_3355_), .Y(_3381_) );
NAND3X1 NAND3X1_173 ( .A(_4239__bF_buf3), .B(_3381_), .C(_3380_), .Y(_3382_) );
NAND3X1 NAND3X1_174 ( .A(_4238__bF_buf2), .B(_3368_), .C(_3382_), .Y(_3383_) );
NAND2X1 NAND2X1_484 ( .A(micro_hash_ucr_pipe17), .B(_3355_), .Y(_3384_) );
NAND3X1 NAND3X1_175 ( .A(_624__bF_buf1), .B(_3384_), .C(_3383_), .Y(_3385_) );
NAND3X1 NAND3X1_176 ( .A(_2816_), .B(_3367_), .C(_3385_), .Y(_3386_) );
AOI21X1 AOI21X1_527 ( .A(micro_hash_ucr_pipe19), .B(_3355_), .C(micro_hash_ucr_pipe20_bF_buf0), .Y(_3387_) );
OAI21X1 OAI21X1_1019 ( .A(_4237__bF_buf2), .B(micro_hash_ucr_a_5_bF_buf3_), .C(_4236__bF_buf2), .Y(_3388_) );
AOI21X1 AOI21X1_528 ( .A(_3387_), .B(_3386_), .C(_3388_), .Y(_3389_) );
OAI21X1 OAI21X1_1020 ( .A(_3354__bF_buf3), .B(_4236__bF_buf1), .C(_4262__bF_buf4), .Y(_3390_) );
NAND2X1 NAND2X1_485 ( .A(micro_hash_ucr_pipe22_bF_buf2), .B(_2551_), .Y(_3391_) );
OAI21X1 OAI21X1_1021 ( .A(_3389_), .B(_3390_), .C(_3391_), .Y(_3392_) );
NAND2X1 NAND2X1_486 ( .A(micro_hash_ucr_pipe23), .B(_3355_), .Y(_3393_) );
OAI21X1 OAI21X1_1022 ( .A(_3392_), .B(micro_hash_ucr_pipe23), .C(_3393_), .Y(_3394_) );
OAI21X1 OAI21X1_1023 ( .A(_2551_), .B(_4233__bF_buf4), .C(_389__bF_buf1), .Y(_3395_) );
AOI21X1 AOI21X1_529 ( .A(_4233__bF_buf4), .B(_3394_), .C(_3395_), .Y(_3396_) );
OAI21X1 OAI21X1_1024 ( .A(_3355_), .B(_389__bF_buf3), .C(_4230__bF_buf4), .Y(_3397_) );
NAND2X1 NAND2X1_487 ( .A(micro_hash_ucr_a_5_bF_buf2_), .B(micro_hash_ucr_pipe26_bF_buf2), .Y(_3398_) );
OAI21X1 OAI21X1_1025 ( .A(_3396_), .B(_3397_), .C(_3398_), .Y(_3399_) );
NAND2X1 NAND2X1_488 ( .A(micro_hash_ucr_pipe27_bF_buf2), .B(_3354__bF_buf2), .Y(_3400_) );
OAI21X1 OAI21X1_1026 ( .A(_3399_), .B(micro_hash_ucr_pipe27_bF_buf2), .C(_3400_), .Y(_3401_) );
OAI21X1 OAI21X1_1027 ( .A(_3401_), .B(micro_hash_ucr_pipe28_bF_buf1), .C(_3366_), .Y(_3402_) );
OAI21X1 OAI21X1_1028 ( .A(_3354__bF_buf2), .B(_219_), .C(_4228__bF_buf3), .Y(_3403_) );
AOI21X1 AOI21X1_530 ( .A(_219_), .B(_3402_), .C(_3403_), .Y(_3404_) );
OAI21X1 OAI21X1_1029 ( .A(_4228__bF_buf4), .B(micro_hash_ucr_a_5_bF_buf1_), .C(_317__bF_buf0), .Y(_3405_) );
AOI21X1 AOI21X1_531 ( .A(micro_hash_ucr_pipe31_bF_buf0), .B(_3355_), .C(micro_hash_ucr_pipe32_bF_buf4), .Y(_3406_) );
OAI21X1 OAI21X1_1030 ( .A(_3404_), .B(_3405_), .C(_3406_), .Y(_3407_) );
NAND2X1 NAND2X1_489 ( .A(micro_hash_ucr_pipe32_bF_buf4), .B(_2551_), .Y(_3408_) );
NAND3X1 NAND3X1_177 ( .A(_318_), .B(_3408_), .C(_3407_), .Y(_3409_) );
NAND2X1 NAND2X1_490 ( .A(micro_hash_ucr_pipe33_bF_buf1), .B(_3355_), .Y(_3410_) );
NAND3X1 NAND3X1_178 ( .A(_4225__bF_buf1), .B(_3410_), .C(_3409_), .Y(_3411_) );
NAND3X1 NAND3X1_179 ( .A(_230__bF_buf1), .B(_3365_), .C(_3411_), .Y(_3412_) );
NAND2X1 NAND2X1_491 ( .A(micro_hash_ucr_pipe35), .B(_3355_), .Y(_3413_) );
AOI21X1 AOI21X1_532 ( .A(_3413_), .B(_3412_), .C(micro_hash_ucr_pipe36_bF_buf1), .Y(_3414_) );
OAI21X1 OAI21X1_1031 ( .A(_2551_), .B(_4224__bF_buf3), .C(_2815_), .Y(_3415_) );
AOI21X1 AOI21X1_533 ( .A(micro_hash_ucr_pipe37_bF_buf3), .B(_3354__bF_buf2), .C(micro_hash_ucr_pipe38_bF_buf0), .Y(_3416_) );
OAI21X1 OAI21X1_1032 ( .A(_3414_), .B(_3415_), .C(_3416_), .Y(_3417_) );
NAND2X1 NAND2X1_492 ( .A(micro_hash_ucr_a_5_bF_buf0_), .B(micro_hash_ucr_pipe38_bF_buf0), .Y(_3418_) );
NAND3X1 NAND3X1_180 ( .A(_2813__bF_buf1), .B(_3418_), .C(_3417_), .Y(_3419_) );
NAND2X1 NAND2X1_493 ( .A(micro_hash_ucr_pipe39), .B(_3354__bF_buf0), .Y(_3420_) );
NAND3X1 NAND3X1_181 ( .A(_296__bF_buf3), .B(_3420_), .C(_3419_), .Y(_3421_) );
NAND3X1 NAND3X1_182 ( .A(_2814_), .B(_3364_), .C(_3421_), .Y(_3422_) );
NAND2X1 NAND2X1_494 ( .A(micro_hash_ucr_pipe41_bF_buf3), .B(_3354__bF_buf0), .Y(_3423_) );
NAND3X1 NAND3X1_183 ( .A(_4220__bF_buf2), .B(_3423_), .C(_3422_), .Y(_3424_) );
NAND3X1 NAND3X1_184 ( .A(_242__bF_buf0), .B(_3363_), .C(_3424_), .Y(_3425_) );
NAND2X1 NAND2X1_495 ( .A(micro_hash_ucr_pipe43), .B(_3354__bF_buf0), .Y(_3426_) );
NAND3X1 NAND3X1_185 ( .A(_4219__bF_buf4), .B(_3426_), .C(_3425_), .Y(_3427_) );
AOI21X1 AOI21X1_534 ( .A(_3362_), .B(_3427_), .C(micro_hash_ucr_pipe45), .Y(_3428_) );
OAI21X1 OAI21X1_1033 ( .A(_3354__bF_buf0), .B(_336_), .C(_4218__bF_buf2), .Y(_3429_) );
AOI21X1 AOI21X1_535 ( .A(micro_hash_ucr_pipe46_bF_buf1), .B(_2551_), .C(micro_hash_ucr_pipe47), .Y(_3430_) );
OAI21X1 OAI21X1_1034 ( .A(_3428_), .B(_3429_), .C(_3430_), .Y(_3431_) );
AOI21X1 AOI21X1_536 ( .A(micro_hash_ucr_pipe47), .B(_3355_), .C(micro_hash_ucr_pipe48_bF_buf2), .Y(_3432_) );
NAND2X1 NAND2X1_496 ( .A(_3432_), .B(_3431_), .Y(_3433_) );
NAND2X1 NAND2X1_497 ( .A(micro_hash_ucr_pipe48_bF_buf2), .B(_2551_), .Y(_3434_) );
NAND3X1 NAND3X1_186 ( .A(_304_), .B(_3434_), .C(_3433_), .Y(_3435_) );
NAND2X1 NAND2X1_498 ( .A(micro_hash_ucr_pipe49_bF_buf1), .B(_3355_), .Y(_3436_) );
NAND3X1 NAND3X1_187 ( .A(_4215__bF_buf2), .B(_3436_), .C(_3435_), .Y(_3437_) );
NAND3X1 NAND3X1_188 ( .A(_255__bF_buf0), .B(_3361_), .C(_3437_), .Y(_3438_) );
NAND2X1 NAND2X1_499 ( .A(micro_hash_ucr_pipe51), .B(_3355_), .Y(_3439_) );
AOI21X1 AOI21X1_537 ( .A(_3439_), .B(_3438_), .C(micro_hash_ucr_pipe52_bF_buf2), .Y(_3440_) );
OAI21X1 OAI21X1_1035 ( .A(_4214__bF_buf0), .B(_2551_), .C(_2812_), .Y(_3441_) );
AOI21X1 AOI21X1_538 ( .A(micro_hash_ucr_pipe53_bF_buf3), .B(_3354__bF_buf1), .C(micro_hash_ucr_pipe54_bF_buf3), .Y(_3442_) );
OAI21X1 OAI21X1_1036 ( .A(_3440_), .B(_3441_), .C(_3442_), .Y(_3443_) );
NAND2X1 NAND2X1_500 ( .A(micro_hash_ucr_pipe54_bF_buf3), .B(micro_hash_ucr_a_5_bF_buf3_), .Y(_3444_) );
NAND3X1 NAND3X1_189 ( .A(_2811__bF_buf1), .B(_3444_), .C(_3443_), .Y(_3445_) );
NAND2X1 NAND2X1_501 ( .A(micro_hash_ucr_pipe55), .B(_3354__bF_buf1), .Y(_3446_) );
NAND3X1 NAND3X1_190 ( .A(_832__bF_buf0), .B(_3446_), .C(_3445_), .Y(_3447_) );
NAND3X1 NAND3X1_191 ( .A(_4212_), .B(_3360_), .C(_3447_), .Y(_3448_) );
NAND2X1 NAND2X1_502 ( .A(micro_hash_ucr_pipe57_bF_buf0), .B(_3354__bF_buf1), .Y(_3449_) );
NAND3X1 NAND3X1_192 ( .A(_4211__bF_buf1), .B(_3449_), .C(_3448_), .Y(_3450_) );
NAND3X1 NAND3X1_193 ( .A(_269_), .B(_3359_), .C(_3450_), .Y(_3451_) );
NAND2X1 NAND2X1_503 ( .A(micro_hash_ucr_pipe59), .B(_3354__bF_buf1), .Y(_3452_) );
NAND3X1 NAND3X1_194 ( .A(_4210__bF_buf1), .B(_3452_), .C(_3451_), .Y(_3453_) );
NAND3X1 NAND3X1_195 ( .A(_4208_), .B(_3358_), .C(_3453_), .Y(_3454_) );
NAND2X1 NAND2X1_504 ( .A(micro_hash_ucr_pipe61_bF_buf2), .B(_3354__bF_buf3), .Y(_3455_) );
NAND3X1 NAND3X1_196 ( .A(_4207__bF_buf4), .B(_3455_), .C(_3454_), .Y(_3456_) );
AOI21X1 AOI21X1_539 ( .A(_3357_), .B(_3456_), .C(micro_hash_ucr_pipe63_bF_buf0), .Y(_3457_) );
OAI21X1 OAI21X1_1037 ( .A(_3354__bF_buf3), .B(_4204_), .C(_278__bF_buf0), .Y(_3458_) );
AOI21X1 AOI21X1_540 ( .A(micro_hash_ucr_pipe64_bF_buf4), .B(_2551_), .C(micro_hash_ucr_pipe65_bF_buf1), .Y(_3459_) );
OAI21X1 OAI21X1_1038 ( .A(_3457_), .B(_3458_), .C(_3459_), .Y(_3460_) );
AOI21X1 AOI21X1_541 ( .A(micro_hash_ucr_pipe65_bF_buf2), .B(_3355_), .C(micro_hash_ucr_pipe66_bF_buf4), .Y(_3461_) );
NOR2X1 NOR2X1_701 ( .A(micro_hash_ucr_a_5_bF_buf2_), .B(_1078__bF_buf1), .Y(_3462_) );
AOI21X1 AOI21X1_542 ( .A(_3461_), .B(_3460_), .C(_3462_), .Y(_3463_) );
OAI21X1 OAI21X1_1039 ( .A(_3354__bF_buf3), .B(_4201__bF_buf3), .C(_4199__bF_buf0), .Y(_3464_) );
AOI21X1 AOI21X1_543 ( .A(_4201__bF_buf3), .B(_3463_), .C(_3464_), .Y(_3465_) );
OAI21X1 OAI21X1_1040 ( .A(_4199__bF_buf0), .B(micro_hash_ucr_a_5_bF_buf1_), .C(_344_), .Y(_3466_) );
OAI21X1 OAI21X1_1041 ( .A(_3465_), .B(_3466_), .C(_3356_), .Y(_126__5_) );
NOR2X1 NOR2X1_702 ( .A(micro_hash_ucr_b_6_bF_buf0_), .B(micro_hash_ucr_c_6_), .Y(_3467_) );
NOR2X1 NOR2X1_703 ( .A(_399__bF_buf2), .B(_2434_), .Y(_3468_) );
NOR2X1 NOR2X1_704 ( .A(_3467_), .B(_3468_), .Y(_3469_) );
INVX8 INVX8_89 ( .A(_3469_), .Y(_3470_) );
NAND2X1 NAND2X1_505 ( .A(micro_hash_ucr_pipe62_bF_buf3), .B(micro_hash_ucr_a_6_bF_buf0_), .Y(_3471_) );
NAND2X1 NAND2X1_506 ( .A(micro_hash_ucr_pipe60_bF_buf2), .B(micro_hash_ucr_a_6_bF_buf3_), .Y(_3472_) );
NAND2X1 NAND2X1_507 ( .A(micro_hash_ucr_pipe58_bF_buf2), .B(micro_hash_ucr_a_6_bF_buf2_), .Y(_3473_) );
NAND2X1 NAND2X1_508 ( .A(micro_hash_ucr_pipe42_bF_buf3), .B(micro_hash_ucr_a_6_bF_buf1_), .Y(_3474_) );
NAND2X1 NAND2X1_509 ( .A(micro_hash_ucr_pipe40_bF_buf0), .B(micro_hash_ucr_a_6_bF_buf0_), .Y(_3475_) );
NAND2X1 NAND2X1_510 ( .A(micro_hash_ucr_a_6_bF_buf3_), .B(micro_hash_ucr_pipe38_bF_buf1), .Y(_3476_) );
NAND2X1 NAND2X1_511 ( .A(micro_hash_ucr_a_6_bF_buf2_), .B(micro_hash_ucr_pipe36_bF_buf2), .Y(_3477_) );
NOR2X1 NOR2X1_705 ( .A(_400_), .B(_4228__bF_buf1), .Y(_3478_) );
NOR2X1 NOR2X1_706 ( .A(_400_), .B(_220__bF_buf4), .Y(_3479_) );
AOI21X1 AOI21X1_544 ( .A(_4263_), .B(_2826_), .C(micro_hash_ucr_a_6_bF_buf1_), .Y(_3480_) );
NOR2X1 NOR2X1_707 ( .A(micro_hash_ucr_pipe9), .B(H_6_), .Y(_3481_) );
NAND2X1 NAND2X1_512 ( .A(_2816_), .B(_4274_), .Y(_3482_) );
AOI22X1 AOI22X1_26 ( .A(_2823_), .B(_3481_), .C(_3482_), .D(_3470_), .Y(_3483_) );
AOI21X1 AOI21X1_545 ( .A(micro_hash_ucr_a_6_bF_buf0_), .B(_4250_), .C(_3483_), .Y(_3484_) );
OAI22X1 OAI22X1_40 ( .A(_207_), .B(_3470_), .C(_3484_), .D(_3480_), .Y(_3485_) );
OAI21X1 OAI21X1_1042 ( .A(_3470_), .B(_4236__bF_buf1), .C(_4262__bF_buf4), .Y(_3486_) );
AOI21X1 AOI21X1_546 ( .A(_4236__bF_buf1), .B(_3485_), .C(_3486_), .Y(_3487_) );
OAI21X1 OAI21X1_1043 ( .A(_4262__bF_buf0), .B(micro_hash_ucr_a_6_bF_buf3_), .C(_4234__bF_buf1), .Y(_3488_) );
AOI21X1 AOI21X1_547 ( .A(micro_hash_ucr_pipe23), .B(_3469_), .C(micro_hash_ucr_pipe24_bF_buf3), .Y(_3489_) );
OAI21X1 OAI21X1_1044 ( .A(_3487_), .B(_3488_), .C(_3489_), .Y(_3490_) );
OAI21X1 OAI21X1_1045 ( .A(micro_hash_ucr_a_6_bF_buf2_), .B(_4233__bF_buf2), .C(_3490_), .Y(_3491_) );
AND2X2 AND2X2_265 ( .A(_3491_), .B(_389__bF_buf2), .Y(_3492_) );
NOR2X1 NOR2X1_708 ( .A(_389__bF_buf2), .B(_3469_), .Y(_3493_) );
OAI21X1 OAI21X1_1046 ( .A(_3492_), .B(_3493_), .C(_4230__bF_buf0), .Y(_3494_) );
OAI21X1 OAI21X1_1047 ( .A(micro_hash_ucr_a_6_bF_buf1_), .B(_4230__bF_buf0), .C(_3494_), .Y(_3495_) );
OR2X2 OR2X2_26 ( .A(_3495_), .B(micro_hash_ucr_pipe27_bF_buf0), .Y(_3496_) );
NAND2X1 NAND2X1_513 ( .A(micro_hash_ucr_pipe27_bF_buf0), .B(_3469_), .Y(_3497_) );
AOI21X1 AOI21X1_548 ( .A(_3497_), .B(_3496_), .C(micro_hash_ucr_pipe28_bF_buf0), .Y(_3498_) );
OAI21X1 OAI21X1_1048 ( .A(_3498_), .B(_3479_), .C(_219_), .Y(_3499_) );
NAND2X1 NAND2X1_514 ( .A(micro_hash_ucr_pipe29), .B(_3469_), .Y(_3500_) );
AOI21X1 AOI21X1_549 ( .A(_3500_), .B(_3499_), .C(micro_hash_ucr_pipe30_bF_buf0), .Y(_3501_) );
OAI21X1 OAI21X1_1049 ( .A(_3501_), .B(_3478_), .C(_317__bF_buf3), .Y(_3502_) );
AOI21X1 AOI21X1_550 ( .A(micro_hash_ucr_pipe31_bF_buf1), .B(_3469_), .C(micro_hash_ucr_pipe32_bF_buf2), .Y(_3503_) );
OAI21X1 OAI21X1_1050 ( .A(_4226__bF_buf3), .B(micro_hash_ucr_a_6_bF_buf0_), .C(_318_), .Y(_3504_) );
AOI21X1 AOI21X1_551 ( .A(_3503_), .B(_3502_), .C(_3504_), .Y(_3505_) );
OAI21X1 OAI21X1_1051 ( .A(_3470_), .B(_318_), .C(_4225__bF_buf2), .Y(_3506_) );
OAI22X1 OAI22X1_41 ( .A(micro_hash_ucr_a_6_bF_buf3_), .B(_4225__bF_buf2), .C(_3505_), .D(_3506_), .Y(_3507_) );
NOR2X1 NOR2X1_709 ( .A(micro_hash_ucr_pipe35), .B(_3507_), .Y(_3508_) );
NOR2X1 NOR2X1_710 ( .A(_230__bF_buf0), .B(_3470_), .Y(_3509_) );
OAI21X1 OAI21X1_1052 ( .A(_3508_), .B(_3509_), .C(_4224__bF_buf0), .Y(_3510_) );
NAND3X1 NAND3X1_197 ( .A(_2815_), .B(_3477_), .C(_3510_), .Y(_3511_) );
OAI21X1 OAI21X1_1053 ( .A(_3468_), .B(_3467_), .C(micro_hash_ucr_pipe37_bF_buf2), .Y(_3512_) );
NAND3X1 NAND3X1_198 ( .A(_701__bF_buf3), .B(_3512_), .C(_3511_), .Y(_3513_) );
NAND3X1 NAND3X1_199 ( .A(_2813__bF_buf3), .B(_3476_), .C(_3513_), .Y(_3514_) );
OAI21X1 OAI21X1_1054 ( .A(_3468_), .B(_3467_), .C(micro_hash_ucr_pipe39), .Y(_3515_) );
NAND3X1 NAND3X1_200 ( .A(_296__bF_buf0), .B(_3515_), .C(_3514_), .Y(_3516_) );
NAND3X1 NAND3X1_201 ( .A(_2814_), .B(_3475_), .C(_3516_), .Y(_3517_) );
OAI21X1 OAI21X1_1055 ( .A(_3468_), .B(_3467_), .C(micro_hash_ucr_pipe41_bF_buf2), .Y(_3518_) );
NAND3X1 NAND3X1_202 ( .A(_4220__bF_buf3), .B(_3518_), .C(_3517_), .Y(_3519_) );
NAND3X1 NAND3X1_203 ( .A(_242__bF_buf3), .B(_3474_), .C(_3519_), .Y(_3520_) );
OAI21X1 OAI21X1_1056 ( .A(_3468_), .B(_3467_), .C(micro_hash_ucr_pipe43), .Y(_3521_) );
NAND3X1 NAND3X1_204 ( .A(_4219__bF_buf4), .B(_3521_), .C(_3520_), .Y(_3522_) );
AOI21X1 AOI21X1_552 ( .A(micro_hash_ucr_pipe44_bF_buf3), .B(micro_hash_ucr_a_6_bF_buf2_), .C(micro_hash_ucr_pipe45), .Y(_3523_) );
OAI21X1 OAI21X1_1057 ( .A(_3469_), .B(_336_), .C(_4218__bF_buf1), .Y(_3524_) );
AOI21X1 AOI21X1_553 ( .A(_3523_), .B(_3522_), .C(_3524_), .Y(_3525_) );
NOR2X1 NOR2X1_711 ( .A(_4218__bF_buf1), .B(_400_), .Y(_3526_) );
OAI21X1 OAI21X1_1058 ( .A(_3525_), .B(_3526_), .C(_249__bF_buf2), .Y(_3527_) );
AOI21X1 AOI21X1_554 ( .A(micro_hash_ucr_pipe47), .B(_3469_), .C(micro_hash_ucr_pipe48_bF_buf4), .Y(_3528_) );
OAI21X1 OAI21X1_1059 ( .A(_4217__bF_buf2), .B(micro_hash_ucr_a_6_bF_buf1_), .C(_304_), .Y(_3529_) );
AOI21X1 AOI21X1_555 ( .A(_3528_), .B(_3527_), .C(_3529_), .Y(_3530_) );
OAI21X1 OAI21X1_1060 ( .A(_3470_), .B(_304_), .C(_4215__bF_buf3), .Y(_3531_) );
OAI22X1 OAI22X1_42 ( .A(_4215__bF_buf3), .B(micro_hash_ucr_a_6_bF_buf0_), .C(_3530_), .D(_3531_), .Y(_3532_) );
OAI21X1 OAI21X1_1061 ( .A(_3469_), .B(_255__bF_buf3), .C(_4214__bF_buf1), .Y(_3533_) );
AOI21X1 AOI21X1_556 ( .A(_255__bF_buf3), .B(_3532_), .C(_3533_), .Y(_3534_) );
NOR2X1 NOR2X1_712 ( .A(_4214__bF_buf4), .B(_400_), .Y(_3535_) );
OAI21X1 OAI21X1_1062 ( .A(_3534_), .B(_3535_), .C(_2812_), .Y(_3536_) );
AOI21X1 AOI21X1_557 ( .A(micro_hash_ucr_pipe53_bF_buf2), .B(_3469_), .C(micro_hash_ucr_pipe54_bF_buf1), .Y(_3537_) );
OAI21X1 OAI21X1_1063 ( .A(_742__bF_buf2), .B(micro_hash_ucr_a_6_bF_buf3_), .C(_2811__bF_buf3), .Y(_3538_) );
AOI21X1 AOI21X1_558 ( .A(_3537_), .B(_3536_), .C(_3538_), .Y(_3539_) );
OAI21X1 OAI21X1_1064 ( .A(_3470_), .B(_2811__bF_buf3), .C(_832__bF_buf1), .Y(_3540_) );
NAND2X1 NAND2X1_515 ( .A(micro_hash_ucr_pipe56_bF_buf3), .B(_400_), .Y(_3541_) );
OAI21X1 OAI21X1_1065 ( .A(_3539_), .B(_3540_), .C(_3541_), .Y(_3542_) );
NAND2X1 NAND2X1_516 ( .A(_4212_), .B(_3542_), .Y(_3543_) );
OAI21X1 OAI21X1_1066 ( .A(_4212_), .B(_3469_), .C(_3543_), .Y(_3544_) );
OAI21X1 OAI21X1_1067 ( .A(_3544_), .B(micro_hash_ucr_pipe58_bF_buf2), .C(_3473_), .Y(_3545_) );
OAI21X1 OAI21X1_1068 ( .A(_3468_), .B(_3467_), .C(micro_hash_ucr_pipe59), .Y(_3546_) );
OAI21X1 OAI21X1_1069 ( .A(_3545_), .B(micro_hash_ucr_pipe59), .C(_3546_), .Y(_3547_) );
OAI21X1 OAI21X1_1070 ( .A(_3547_), .B(micro_hash_ucr_pipe60_bF_buf2), .C(_3472_), .Y(_3548_) );
OAI21X1 OAI21X1_1071 ( .A(_3468_), .B(_3467_), .C(micro_hash_ucr_pipe61_bF_buf1), .Y(_3549_) );
OAI21X1 OAI21X1_1072 ( .A(_3548_), .B(micro_hash_ucr_pipe61_bF_buf1), .C(_3549_), .Y(_3550_) );
OAI21X1 OAI21X1_1073 ( .A(_3550_), .B(micro_hash_ucr_pipe62_bF_buf3), .C(_3471_), .Y(_3551_) );
NAND2X1 NAND2X1_517 ( .A(_4204_), .B(_3551_), .Y(_3552_) );
OAI21X1 OAI21X1_1074 ( .A(_4204_), .B(_3470_), .C(_3552_), .Y(_3553_) );
AOI21X1 AOI21X1_559 ( .A(micro_hash_ucr_pipe64_bF_buf2), .B(_400_), .C(micro_hash_ucr_pipe65_bF_buf3), .Y(_3554_) );
OAI21X1 OAI21X1_1075 ( .A(_3553_), .B(micro_hash_ucr_pipe64_bF_buf2), .C(_3554_), .Y(_3555_) );
AOI21X1 AOI21X1_560 ( .A(micro_hash_ucr_pipe65_bF_buf0), .B(_3469_), .C(micro_hash_ucr_pipe66_bF_buf2), .Y(_3556_) );
AOI22X1 AOI22X1_27 ( .A(micro_hash_ucr_pipe66_bF_buf2), .B(_400_), .C(_3555_), .D(_3556_), .Y(_3557_) );
OAI21X1 OAI21X1_1076 ( .A(_3470_), .B(_4201__bF_buf2), .C(_4199__bF_buf4), .Y(_3558_) );
AOI21X1 AOI21X1_561 ( .A(_4201__bF_buf2), .B(_3557_), .C(_3558_), .Y(_3559_) );
OAI21X1 OAI21X1_1077 ( .A(_4199__bF_buf5), .B(micro_hash_ucr_a_6_bF_buf2_), .C(_344_), .Y(_3560_) );
OAI22X1 OAI22X1_43 ( .A(_2181_), .B(_3470_), .C(_3559_), .D(_3560_), .Y(_126__6_) );
NOR2X1 NOR2X1_713 ( .A(micro_hash_ucr_b_7_bF_buf2_), .B(micro_hash_ucr_c_7_), .Y(_3561_) );
NAND2X1 NAND2X1_518 ( .A(micro_hash_ucr_b_7_bF_buf1_), .B(micro_hash_ucr_c_7_), .Y(_3562_) );
INVX4 INVX4_49 ( .A(_3562_), .Y(_3563_) );
NOR2X1 NOR2X1_714 ( .A(_3561_), .B(_3563_), .Y(_3564_) );
INVX8 INVX8_90 ( .A(_3564_), .Y(_3565_) );
INVX8 INVX8_91 ( .A(micro_hash_ucr_a_7_bF_buf0_), .Y(_3566_) );
NAND2X1 NAND2X1_519 ( .A(micro_hash_ucr_pipe60_bF_buf4), .B(_3566_), .Y(_3567_) );
NAND2X1 NAND2X1_520 ( .A(micro_hash_ucr_pipe58_bF_buf3), .B(_3566_), .Y(_3568_) );
NAND2X1 NAND2X1_521 ( .A(micro_hash_ucr_pipe50_bF_buf3), .B(_3566_), .Y(_3569_) );
NAND2X1 NAND2X1_522 ( .A(micro_hash_ucr_pipe48_bF_buf2), .B(_3566_), .Y(_3570_) );
NAND2X1 NAND2X1_523 ( .A(micro_hash_ucr_pipe42_bF_buf4), .B(micro_hash_ucr_a_7_bF_buf3_), .Y(_3571_) );
NAND2X1 NAND2X1_524 ( .A(micro_hash_ucr_pipe40_bF_buf2), .B(micro_hash_ucr_a_7_bF_buf2_), .Y(_3572_) );
NAND2X1 NAND2X1_525 ( .A(micro_hash_ucr_a_7_bF_buf1_), .B(micro_hash_ucr_pipe38_bF_buf1), .Y(_3573_) );
NAND2X1 NAND2X1_526 ( .A(micro_hash_ucr_a_7_bF_buf0_), .B(micro_hash_ucr_pipe32_bF_buf1), .Y(_3574_) );
AOI21X1 AOI21X1_562 ( .A(_4240_), .B(_4279_), .C(_3565_), .Y(_3575_) );
NOR2X1 NOR2X1_715 ( .A(H_7_), .B(_4266_), .Y(_3576_) );
AOI22X1 AOI22X1_28 ( .A(_4253_), .B(_3576_), .C(_4273_), .D(_3565_), .Y(_3577_) );
AOI21X1 AOI21X1_563 ( .A(_4260_), .B(_3577_), .C(_3575_), .Y(_3578_) );
OAI21X1 OAI21X1_1078 ( .A(_4248_), .B(_3577_), .C(micro_hash_ucr_a_7_bF_buf3_), .Y(_3579_) );
OAI21X1 OAI21X1_1079 ( .A(_3578_), .B(micro_hash_ucr_pipe16), .C(_3579_), .Y(_3580_) );
OAI21X1 OAI21X1_1080 ( .A(_3565_), .B(_4238__bF_buf1), .C(_624__bF_buf1), .Y(_3581_) );
AOI21X1 AOI21X1_564 ( .A(_4238__bF_buf1), .B(_3580_), .C(_3581_), .Y(_3582_) );
OAI21X1 OAI21X1_1081 ( .A(_624__bF_buf2), .B(micro_hash_ucr_a_7_bF_buf2_), .C(_2816_), .Y(_3583_) );
AOI21X1 AOI21X1_565 ( .A(micro_hash_ucr_pipe19), .B(_3564_), .C(micro_hash_ucr_pipe20_bF_buf2), .Y(_3584_) );
OAI21X1 OAI21X1_1082 ( .A(_3582_), .B(_3583_), .C(_3584_), .Y(_3585_) );
NAND2X1 NAND2X1_527 ( .A(micro_hash_ucr_pipe20_bF_buf0), .B(_3566_), .Y(_3586_) );
NAND3X1 NAND3X1_205 ( .A(_4236__bF_buf2), .B(_3586_), .C(_3585_), .Y(_3587_) );
AOI21X1 AOI21X1_566 ( .A(micro_hash_ucr_pipe21), .B(_3564_), .C(micro_hash_ucr_pipe22_bF_buf3), .Y(_3588_) );
OAI21X1 OAI21X1_1083 ( .A(_4262__bF_buf2), .B(micro_hash_ucr_a_7_bF_buf1_), .C(_4234__bF_buf3), .Y(_3589_) );
AOI21X1 AOI21X1_567 ( .A(_3588_), .B(_3587_), .C(_3589_), .Y(_3590_) );
OAI21X1 OAI21X1_1084 ( .A(_3565_), .B(_4234__bF_buf0), .C(_4233__bF_buf4), .Y(_3591_) );
OAI22X1 OAI22X1_44 ( .A(micro_hash_ucr_a_7_bF_buf0_), .B(_4233__bF_buf4), .C(_3590_), .D(_3591_), .Y(_3592_) );
NAND2X1 NAND2X1_528 ( .A(micro_hash_ucr_pipe25_bF_buf1), .B(_3564_), .Y(_3593_) );
OAI21X1 OAI21X1_1085 ( .A(_3592_), .B(micro_hash_ucr_pipe25_bF_buf1), .C(_3593_), .Y(_3594_) );
NAND2X1 NAND2X1_529 ( .A(micro_hash_ucr_pipe26_bF_buf1), .B(_3566_), .Y(_3595_) );
OAI21X1 OAI21X1_1086 ( .A(_3594_), .B(micro_hash_ucr_pipe26_bF_buf2), .C(_3595_), .Y(_3596_) );
NAND2X1 NAND2X1_530 ( .A(micro_hash_ucr_pipe27_bF_buf3), .B(_3564_), .Y(_3597_) );
OAI21X1 OAI21X1_1087 ( .A(_3596_), .B(micro_hash_ucr_pipe27_bF_buf2), .C(_3597_), .Y(_3598_) );
NAND2X1 NAND2X1_531 ( .A(micro_hash_ucr_pipe28_bF_buf1), .B(_3566_), .Y(_3599_) );
OAI21X1 OAI21X1_1088 ( .A(_3598_), .B(micro_hash_ucr_pipe28_bF_buf1), .C(_3599_), .Y(_3600_) );
NAND2X1 NAND2X1_532 ( .A(micro_hash_ucr_pipe29), .B(_3564_), .Y(_3601_) );
OAI21X1 OAI21X1_1089 ( .A(_3600_), .B(micro_hash_ucr_pipe29), .C(_3601_), .Y(_3602_) );
NAND2X1 NAND2X1_533 ( .A(_4228__bF_buf0), .B(_3602_), .Y(_3603_) );
OAI21X1 OAI21X1_1090 ( .A(_3566_), .B(_4228__bF_buf0), .C(_3603_), .Y(_3604_) );
OAI21X1 OAI21X1_1091 ( .A(_3563_), .B(_3561_), .C(micro_hash_ucr_pipe31_bF_buf3), .Y(_3605_) );
OAI21X1 OAI21X1_1092 ( .A(_3604_), .B(micro_hash_ucr_pipe31_bF_buf2), .C(_3605_), .Y(_3606_) );
OAI21X1 OAI21X1_1093 ( .A(_3606_), .B(micro_hash_ucr_pipe32_bF_buf1), .C(_3574_), .Y(_3607_) );
NAND2X1 NAND2X1_534 ( .A(_318_), .B(_3607_), .Y(_3608_) );
OAI21X1 OAI21X1_1094 ( .A(_318_), .B(_3565_), .C(_3608_), .Y(_3609_) );
AOI21X1 AOI21X1_568 ( .A(micro_hash_ucr_pipe34_bF_buf1), .B(_3566_), .C(micro_hash_ucr_pipe35), .Y(_3610_) );
OAI21X1 OAI21X1_1095 ( .A(_3609_), .B(micro_hash_ucr_pipe34_bF_buf1), .C(_3610_), .Y(_3611_) );
AOI21X1 AOI21X1_569 ( .A(micro_hash_ucr_pipe35), .B(_3564_), .C(micro_hash_ucr_pipe36_bF_buf3), .Y(_3612_) );
AOI22X1 AOI22X1_29 ( .A(_3566_), .B(micro_hash_ucr_pipe36_bF_buf3), .C(_3611_), .D(_3612_), .Y(_3613_) );
OAI21X1 OAI21X1_1096 ( .A(_3563_), .B(_3561_), .C(micro_hash_ucr_pipe37_bF_buf2), .Y(_3614_) );
OAI21X1 OAI21X1_1097 ( .A(_3613_), .B(micro_hash_ucr_pipe37_bF_buf2), .C(_3614_), .Y(_3615_) );
OAI21X1 OAI21X1_1098 ( .A(_3615_), .B(micro_hash_ucr_pipe38_bF_buf1), .C(_3573_), .Y(_3616_) );
OAI21X1 OAI21X1_1099 ( .A(_3563_), .B(_3561_), .C(micro_hash_ucr_pipe39), .Y(_3617_) );
OAI21X1 OAI21X1_1100 ( .A(_3616_), .B(micro_hash_ucr_pipe39), .C(_3617_), .Y(_3618_) );
OAI21X1 OAI21X1_1101 ( .A(_3618_), .B(micro_hash_ucr_pipe40_bF_buf2), .C(_3572_), .Y(_3619_) );
OAI21X1 OAI21X1_1102 ( .A(_3563_), .B(_3561_), .C(micro_hash_ucr_pipe41_bF_buf1), .Y(_3620_) );
OAI21X1 OAI21X1_1103 ( .A(_3619_), .B(micro_hash_ucr_pipe41_bF_buf1), .C(_3620_), .Y(_3621_) );
OAI21X1 OAI21X1_1104 ( .A(_3621_), .B(micro_hash_ucr_pipe42_bF_buf4), .C(_3571_), .Y(_3622_) );
OAI21X1 OAI21X1_1105 ( .A(_3565_), .B(_242__bF_buf1), .C(_4219__bF_buf0), .Y(_3623_) );
AOI21X1 AOI21X1_570 ( .A(_242__bF_buf1), .B(_3622_), .C(_3623_), .Y(_3624_) );
OAI21X1 OAI21X1_1106 ( .A(_4219__bF_buf0), .B(micro_hash_ucr_a_7_bF_buf3_), .C(_336_), .Y(_3625_) );
AOI21X1 AOI21X1_571 ( .A(micro_hash_ucr_pipe45), .B(_3564_), .C(micro_hash_ucr_pipe46_bF_buf4), .Y(_3626_) );
OAI21X1 OAI21X1_1107 ( .A(_3624_), .B(_3625_), .C(_3626_), .Y(_3627_) );
NAND2X1 NAND2X1_535 ( .A(micro_hash_ucr_pipe46_bF_buf4), .B(_3566_), .Y(_3628_) );
AOI21X1 AOI21X1_572 ( .A(_3628_), .B(_3627_), .C(micro_hash_ucr_pipe47), .Y(_3629_) );
NOR2X1 NOR2X1_716 ( .A(_249__bF_buf3), .B(_3564_), .Y(_3630_) );
OAI21X1 OAI21X1_1108 ( .A(_3629_), .B(_3630_), .C(_4217__bF_buf3), .Y(_3631_) );
AOI21X1 AOI21X1_573 ( .A(_3570_), .B(_3631_), .C(micro_hash_ucr_pipe49_bF_buf2), .Y(_3632_) );
NOR2X1 NOR2X1_717 ( .A(_304_), .B(_3564_), .Y(_3633_) );
OAI21X1 OAI21X1_1109 ( .A(_3632_), .B(_3633_), .C(_4215__bF_buf2), .Y(_3634_) );
NAND3X1 NAND3X1_206 ( .A(_255__bF_buf2), .B(_3569_), .C(_3634_), .Y(_3635_) );
AOI21X1 AOI21X1_574 ( .A(micro_hash_ucr_pipe51), .B(_3564_), .C(micro_hash_ucr_pipe52_bF_buf0), .Y(_3636_) );
OAI21X1 OAI21X1_1110 ( .A(_4214__bF_buf2), .B(micro_hash_ucr_a_7_bF_buf2_), .C(_2812_), .Y(_3637_) );
AOI21X1 AOI21X1_575 ( .A(_3636_), .B(_3635_), .C(_3637_), .Y(_3638_) );
OAI21X1 OAI21X1_1111 ( .A(_3565_), .B(_2812_), .C(_742__bF_buf1), .Y(_3639_) );
OAI22X1 OAI22X1_45 ( .A(_742__bF_buf1), .B(micro_hash_ucr_a_7_bF_buf1_), .C(_3638_), .D(_3639_), .Y(_3640_) );
OAI21X1 OAI21X1_1112 ( .A(_3564_), .B(_2811__bF_buf2), .C(_832__bF_buf4), .Y(_3641_) );
AOI21X1 AOI21X1_576 ( .A(_2811__bF_buf2), .B(_3640_), .C(_3641_), .Y(_3642_) );
NOR2X1 NOR2X1_718 ( .A(_832__bF_buf2), .B(_3566_), .Y(_3643_) );
OAI21X1 OAI21X1_1113 ( .A(_3642_), .B(_3643_), .C(_4212_), .Y(_3644_) );
NAND2X1 NAND2X1_536 ( .A(micro_hash_ucr_pipe57_bF_buf1), .B(_3564_), .Y(_3645_) );
NAND3X1 NAND3X1_207 ( .A(_4211__bF_buf0), .B(_3645_), .C(_3644_), .Y(_3646_) );
NAND3X1 NAND3X1_208 ( .A(_269_), .B(_3568_), .C(_3646_), .Y(_3647_) );
NAND2X1 NAND2X1_537 ( .A(micro_hash_ucr_pipe59), .B(_3564_), .Y(_3648_) );
NAND3X1 NAND3X1_209 ( .A(_4210__bF_buf3), .B(_3648_), .C(_3647_), .Y(_3649_) );
NAND3X1 NAND3X1_210 ( .A(_4208_), .B(_3567_), .C(_3649_), .Y(_3650_) );
NAND2X1 NAND2X1_538 ( .A(micro_hash_ucr_pipe61_bF_buf3), .B(_3564_), .Y(_3651_) );
AOI21X1 AOI21X1_577 ( .A(_3651_), .B(_3650_), .C(micro_hash_ucr_pipe62_bF_buf2), .Y(_3652_) );
OAI21X1 OAI21X1_1114 ( .A(_4207__bF_buf2), .B(_3566_), .C(_4204_), .Y(_3653_) );
AOI21X1 AOI21X1_578 ( .A(micro_hash_ucr_pipe63_bF_buf2), .B(_3565_), .C(micro_hash_ucr_pipe64_bF_buf0), .Y(_3654_) );
OAI21X1 OAI21X1_1115 ( .A(_3652_), .B(_3653_), .C(_3654_), .Y(_3655_) );
NAND2X1 NAND2X1_539 ( .A(micro_hash_ucr_pipe64_bF_buf2), .B(micro_hash_ucr_a_7_bF_buf0_), .Y(_3656_) );
NAND3X1 NAND3X1_211 ( .A(_279_), .B(_3656_), .C(_3655_), .Y(_3657_) );
OAI21X1 OAI21X1_1116 ( .A(_3563_), .B(_3561_), .C(micro_hash_ucr_pipe65_bF_buf3), .Y(_3658_) );
NAND3X1 NAND3X1_212 ( .A(_1078__bF_buf3), .B(_3658_), .C(_3657_), .Y(_3659_) );
OAI21X1 OAI21X1_1117 ( .A(_1078__bF_buf3), .B(_3566_), .C(_3659_), .Y(_3660_) );
OAI21X1 OAI21X1_1118 ( .A(_3565_), .B(_4201__bF_buf2), .C(_4199__bF_buf4), .Y(_3661_) );
AOI21X1 AOI21X1_579 ( .A(_4201__bF_buf2), .B(_3660_), .C(_3661_), .Y(_3662_) );
OAI21X1 OAI21X1_1119 ( .A(_4199__bF_buf4), .B(micro_hash_ucr_a_7_bF_buf3_), .C(_344_), .Y(_3663_) );
OAI22X1 OAI22X1_46 ( .A(_2181_), .B(_3565_), .C(_3662_), .D(_3663_), .Y(_126__7_) );
INVX1 INVX1_334 ( .A(_4256_), .Y(_3664_) );
NOR2X1 NOR2X1_719 ( .A(micro_hash_ucr_pipe15), .B(_4280_), .Y(_3665_) );
NAND3X1 NAND3X1_213 ( .A(_4243_), .B(_4258_), .C(_4241__bF_buf2), .Y(_3666_) );
OAI21X1 OAI21X1_1120 ( .A(_3664_), .B(_3666_), .C(_3665_), .Y(_3667_) );
OR2X2 OR2X2_27 ( .A(_4268_), .B(_3666_), .Y(_3668_) );
NOR2X1 NOR2X1_720 ( .A(H_8_), .B(_3668_), .Y(_3669_) );
OAI21X1 OAI21X1_1121 ( .A(_3667_), .B(_3669_), .C(_4239__bF_buf0), .Y(_3670_) );
AOI21X1 AOI21X1_580 ( .A(_4238__bF_buf3), .B(_3670_), .C(micro_hash_ucr_pipe18_bF_buf0), .Y(_3671_) );
NAND2X1 NAND2X1_540 ( .A(_4239__bF_buf4), .B(_624__bF_buf3), .Y(_3672_) );
OAI21X1 OAI21X1_1122 ( .A(_3668_), .B(_3672_), .C(_330_), .Y(_3673_) );
NAND2X1 NAND2X1_541 ( .A(_2816_), .B(_3673_), .Y(_3674_) );
OAI21X1 OAI21X1_1123 ( .A(_3671_), .B(_3674_), .C(_4237__bF_buf3), .Y(_3675_) );
AOI21X1 AOI21X1_581 ( .A(micro_hash_ucr_pipe20_bF_buf3), .B(_330_), .C(micro_hash_ucr_pipe21), .Y(_3676_) );
AOI21X1 AOI21X1_582 ( .A(_3676_), .B(_3675_), .C(micro_hash_ucr_pipe22_bF_buf0), .Y(_3677_) );
OAI21X1 OAI21X1_1124 ( .A(_4262__bF_buf0), .B(micro_hash_ucr_b_0_bF_buf2_), .C(_4234__bF_buf2), .Y(_3678_) );
OAI21X1 OAI21X1_1125 ( .A(_3677_), .B(_3678_), .C(_4233__bF_buf3), .Y(_3679_) );
AOI21X1 AOI21X1_583 ( .A(micro_hash_ucr_pipe24_bF_buf2), .B(_330_), .C(micro_hash_ucr_pipe25_bF_buf2), .Y(_3680_) );
AOI21X1 AOI21X1_584 ( .A(_3680_), .B(_3679_), .C(micro_hash_ucr_pipe26_bF_buf3), .Y(_3681_) );
OAI21X1 OAI21X1_1126 ( .A(_4230__bF_buf2), .B(micro_hash_ucr_b_0_bF_buf1_), .C(_4229_), .Y(_3682_) );
OAI21X1 OAI21X1_1127 ( .A(_3681_), .B(_3682_), .C(_220__bF_buf4), .Y(_3683_) );
AOI21X1 AOI21X1_585 ( .A(micro_hash_ucr_pipe28_bF_buf2), .B(_330_), .C(micro_hash_ucr_pipe29), .Y(_3684_) );
AOI21X1 AOI21X1_586 ( .A(_3684_), .B(_3683_), .C(micro_hash_ucr_pipe30_bF_buf0), .Y(_3685_) );
OAI21X1 OAI21X1_1128 ( .A(_4228__bF_buf1), .B(micro_hash_ucr_b_0_bF_buf0_), .C(_317__bF_buf3), .Y(_3686_) );
OAI21X1 OAI21X1_1129 ( .A(_3685_), .B(_3686_), .C(_4226__bF_buf1), .Y(_3687_) );
AOI21X1 AOI21X1_587 ( .A(micro_hash_ucr_pipe32_bF_buf2), .B(_330_), .C(micro_hash_ucr_pipe33_bF_buf2), .Y(_3688_) );
AOI21X1 AOI21X1_588 ( .A(_3688_), .B(_3687_), .C(micro_hash_ucr_pipe34_bF_buf3), .Y(_3689_) );
OAI21X1 OAI21X1_1130 ( .A(_4225__bF_buf0), .B(micro_hash_ucr_b_0_bF_buf3_), .C(_230__bF_buf0), .Y(_3690_) );
OAI21X1 OAI21X1_1131 ( .A(_3689_), .B(_3690_), .C(_4224__bF_buf2), .Y(_3691_) );
AOI21X1 AOI21X1_589 ( .A(micro_hash_ucr_pipe36_bF_buf0), .B(_330_), .C(micro_hash_ucr_pipe37_bF_buf1), .Y(_3692_) );
AOI21X1 AOI21X1_590 ( .A(_3692_), .B(_3691_), .C(micro_hash_ucr_pipe38_bF_buf2), .Y(_3693_) );
OAI21X1 OAI21X1_1132 ( .A(_701__bF_buf3), .B(micro_hash_ucr_b_0_bF_buf2_), .C(_2813__bF_buf3), .Y(_3694_) );
OAI21X1 OAI21X1_1133 ( .A(_3693_), .B(_3694_), .C(_296__bF_buf1), .Y(_3695_) );
AOI21X1 AOI21X1_591 ( .A(micro_hash_ucr_pipe40_bF_buf1), .B(_330_), .C(micro_hash_ucr_pipe41_bF_buf3), .Y(_3696_) );
AOI21X1 AOI21X1_592 ( .A(_3696_), .B(_3695_), .C(micro_hash_ucr_pipe42_bF_buf3), .Y(_3697_) );
OAI21X1 OAI21X1_1134 ( .A(_4220__bF_buf1), .B(micro_hash_ucr_b_0_bF_buf1_), .C(_242__bF_buf2), .Y(_3698_) );
OAI21X1 OAI21X1_1135 ( .A(_3697_), .B(_3698_), .C(_4219__bF_buf3), .Y(_3699_) );
AOI21X1 AOI21X1_593 ( .A(micro_hash_ucr_pipe44_bF_buf0), .B(_330_), .C(micro_hash_ucr_pipe45), .Y(_3700_) );
AOI21X1 AOI21X1_594 ( .A(_3700_), .B(_3699_), .C(micro_hash_ucr_pipe46_bF_buf1), .Y(_3701_) );
OAI21X1 OAI21X1_1136 ( .A(_4218__bF_buf2), .B(micro_hash_ucr_b_0_bF_buf0_), .C(_249__bF_buf1), .Y(_3702_) );
OAI21X1 OAI21X1_1137 ( .A(_3701_), .B(_3702_), .C(_4217__bF_buf0), .Y(_3703_) );
AOI21X1 AOI21X1_595 ( .A(micro_hash_ucr_pipe48_bF_buf2), .B(_330_), .C(micro_hash_ucr_pipe49_bF_buf0), .Y(_3704_) );
AOI21X1 AOI21X1_596 ( .A(_3704_), .B(_3703_), .C(micro_hash_ucr_pipe50_bF_buf1), .Y(_3705_) );
OAI21X1 OAI21X1_1138 ( .A(_4215__bF_buf0), .B(micro_hash_ucr_b_0_bF_buf3_), .C(_255__bF_buf2), .Y(_3706_) );
OAI21X1 OAI21X1_1139 ( .A(_3705_), .B(_3706_), .C(_4214__bF_buf2), .Y(_3707_) );
AOI21X1 AOI21X1_597 ( .A(micro_hash_ucr_pipe52_bF_buf0), .B(_330_), .C(micro_hash_ucr_pipe53_bF_buf0), .Y(_3708_) );
AOI21X1 AOI21X1_598 ( .A(_3708_), .B(_3707_), .C(micro_hash_ucr_pipe54_bF_buf4), .Y(_3709_) );
OAI21X1 OAI21X1_1140 ( .A(_742__bF_buf1), .B(micro_hash_ucr_b_0_bF_buf2_), .C(_2811__bF_buf0), .Y(_3710_) );
OAI21X1 OAI21X1_1141 ( .A(_3709_), .B(_3710_), .C(_832__bF_buf2), .Y(_3711_) );
AOI21X1 AOI21X1_599 ( .A(micro_hash_ucr_pipe56_bF_buf0), .B(_330_), .C(micro_hash_ucr_pipe57_bF_buf2), .Y(_3712_) );
AOI21X1 AOI21X1_600 ( .A(_3712_), .B(_3711_), .C(micro_hash_ucr_pipe58_bF_buf3), .Y(_3713_) );
OAI21X1 OAI21X1_1142 ( .A(_4211__bF_buf0), .B(micro_hash_ucr_b_0_bF_buf1_), .C(_269_), .Y(_3714_) );
OAI21X1 OAI21X1_1143 ( .A(_3713_), .B(_3714_), .C(_4210__bF_buf3), .Y(_3715_) );
AOI21X1 AOI21X1_601 ( .A(micro_hash_ucr_pipe60_bF_buf3), .B(_330_), .C(micro_hash_ucr_pipe61_bF_buf0), .Y(_3716_) );
AOI21X1 AOI21X1_602 ( .A(_3716_), .B(_3715_), .C(micro_hash_ucr_pipe62_bF_buf3), .Y(_3717_) );
OAI21X1 OAI21X1_1144 ( .A(_4207__bF_buf2), .B(micro_hash_ucr_b_0_bF_buf0_), .C(_4204_), .Y(_3718_) );
OAI21X1 OAI21X1_1145 ( .A(_3717_), .B(_3718_), .C(_278__bF_buf1), .Y(_3719_) );
AOI21X1 AOI21X1_603 ( .A(micro_hash_ucr_pipe64_bF_buf0), .B(_330_), .C(micro_hash_ucr_pipe65_bF_buf0), .Y(_3720_) );
AOI21X1 AOI21X1_604 ( .A(_3720_), .B(_3719_), .C(micro_hash_ucr_pipe66_bF_buf2), .Y(_3721_) );
OAI21X1 OAI21X1_1146 ( .A(_1078__bF_buf2), .B(micro_hash_ucr_b_0_bF_buf3_), .C(_4201__bF_buf0), .Y(_3722_) );
OAI21X1 OAI21X1_1147 ( .A(_3721_), .B(_3722_), .C(_4199__bF_buf1), .Y(_3723_) );
OAI21X1 OAI21X1_1148 ( .A(_4199__bF_buf1), .B(micro_hash_ucr_b_0_bF_buf2_), .C(_3723_), .Y(_3724_) );
NOR2X1 NOR2X1_721 ( .A(_345_), .B(_3724_), .Y(_127__0_) );
NOR2X1 NOR2X1_722 ( .A(H_9_), .B(_3668_), .Y(_3725_) );
OAI21X1 OAI21X1_1149 ( .A(_3667_), .B(_3725_), .C(_4239__bF_buf4), .Y(_3726_) );
AOI21X1 AOI21X1_605 ( .A(_4238__bF_buf3), .B(_3726_), .C(micro_hash_ucr_pipe18_bF_buf2), .Y(_3727_) );
OAI21X1 OAI21X1_1150 ( .A(_3668_), .B(_3672_), .C(_2448_), .Y(_3728_) );
NAND2X1 NAND2X1_542 ( .A(_2816_), .B(_3728_), .Y(_3729_) );
OAI21X1 OAI21X1_1151 ( .A(_3727_), .B(_3729_), .C(_4237__bF_buf3), .Y(_3730_) );
AOI21X1 AOI21X1_606 ( .A(micro_hash_ucr_pipe20_bF_buf3), .B(_2448_), .C(micro_hash_ucr_pipe21), .Y(_3731_) );
AOI21X1 AOI21X1_607 ( .A(_3731_), .B(_3730_), .C(micro_hash_ucr_pipe22_bF_buf0), .Y(_3732_) );
OAI21X1 OAI21X1_1152 ( .A(_4262__bF_buf3), .B(micro_hash_ucr_b_1_bF_buf2_), .C(_4234__bF_buf0), .Y(_3733_) );
OAI21X1 OAI21X1_1153 ( .A(_3732_), .B(_3733_), .C(_4233__bF_buf3), .Y(_3734_) );
AOI21X1 AOI21X1_608 ( .A(micro_hash_ucr_pipe24_bF_buf2), .B(_2448_), .C(micro_hash_ucr_pipe25_bF_buf0), .Y(_3735_) );
AOI21X1 AOI21X1_609 ( .A(_3735_), .B(_3734_), .C(micro_hash_ucr_pipe26_bF_buf3), .Y(_3736_) );
OAI21X1 OAI21X1_1154 ( .A(_4230__bF_buf2), .B(micro_hash_ucr_b_1_bF_buf1_), .C(_4229_), .Y(_3737_) );
OAI21X1 OAI21X1_1155 ( .A(_3736_), .B(_3737_), .C(_220__bF_buf1), .Y(_3738_) );
AOI21X1 AOI21X1_610 ( .A(micro_hash_ucr_pipe28_bF_buf2), .B(_2448_), .C(micro_hash_ucr_pipe29), .Y(_3739_) );
AOI21X1 AOI21X1_611 ( .A(_3739_), .B(_3738_), .C(micro_hash_ucr_pipe30_bF_buf3), .Y(_3740_) );
OAI21X1 OAI21X1_1156 ( .A(_4228__bF_buf1), .B(micro_hash_ucr_b_1_bF_buf0_), .C(_317__bF_buf2), .Y(_3741_) );
OAI21X1 OAI21X1_1157 ( .A(_3740_), .B(_3741_), .C(_4226__bF_buf1), .Y(_3742_) );
AOI21X1 AOI21X1_612 ( .A(micro_hash_ucr_pipe32_bF_buf0), .B(_2448_), .C(micro_hash_ucr_pipe33_bF_buf0), .Y(_3743_) );
AOI21X1 AOI21X1_613 ( .A(_3743_), .B(_3742_), .C(micro_hash_ucr_pipe34_bF_buf3), .Y(_3744_) );
OAI21X1 OAI21X1_1158 ( .A(_4225__bF_buf0), .B(micro_hash_ucr_b_1_bF_buf3_), .C(_230__bF_buf2), .Y(_3745_) );
OAI21X1 OAI21X1_1159 ( .A(_3744_), .B(_3745_), .C(_4224__bF_buf2), .Y(_3746_) );
AOI21X1 AOI21X1_614 ( .A(micro_hash_ucr_pipe36_bF_buf0), .B(_2448_), .C(micro_hash_ucr_pipe37_bF_buf1), .Y(_3747_) );
AOI21X1 AOI21X1_615 ( .A(_3747_), .B(_3746_), .C(micro_hash_ucr_pipe38_bF_buf2), .Y(_3748_) );
OAI21X1 OAI21X1_1160 ( .A(_701__bF_buf0), .B(micro_hash_ucr_b_1_bF_buf2_), .C(_2813__bF_buf2), .Y(_3749_) );
OAI21X1 OAI21X1_1161 ( .A(_3748_), .B(_3749_), .C(_296__bF_buf1), .Y(_3750_) );
AOI21X1 AOI21X1_616 ( .A(micro_hash_ucr_pipe40_bF_buf1), .B(_2448_), .C(micro_hash_ucr_pipe41_bF_buf3), .Y(_3751_) );
AOI21X1 AOI21X1_617 ( .A(_3751_), .B(_3750_), .C(micro_hash_ucr_pipe42_bF_buf0), .Y(_3752_) );
OAI21X1 OAI21X1_1162 ( .A(_4220__bF_buf1), .B(micro_hash_ucr_b_1_bF_buf1_), .C(_242__bF_buf2), .Y(_3753_) );
OAI21X1 OAI21X1_1163 ( .A(_3752_), .B(_3753_), .C(_4219__bF_buf3), .Y(_3754_) );
AOI21X1 AOI21X1_618 ( .A(micro_hash_ucr_pipe44_bF_buf0), .B(_2448_), .C(micro_hash_ucr_pipe45), .Y(_3755_) );
AOI21X1 AOI21X1_619 ( .A(_3755_), .B(_3754_), .C(micro_hash_ucr_pipe46_bF_buf1), .Y(_3756_) );
OAI21X1 OAI21X1_1164 ( .A(_4218__bF_buf0), .B(micro_hash_ucr_b_1_bF_buf0_), .C(_249__bF_buf1), .Y(_3757_) );
OAI21X1 OAI21X1_1165 ( .A(_3756_), .B(_3757_), .C(_4217__bF_buf0), .Y(_3758_) );
AOI21X1 AOI21X1_620 ( .A(micro_hash_ucr_pipe48_bF_buf3), .B(_2448_), .C(micro_hash_ucr_pipe49_bF_buf0), .Y(_3759_) );
AOI21X1 AOI21X1_621 ( .A(_3759_), .B(_3758_), .C(micro_hash_ucr_pipe50_bF_buf1), .Y(_3760_) );
OAI21X1 OAI21X1_1166 ( .A(_4215__bF_buf0), .B(micro_hash_ucr_b_1_bF_buf3_), .C(_255__bF_buf1), .Y(_3761_) );
OAI21X1 OAI21X1_1167 ( .A(_3760_), .B(_3761_), .C(_4214__bF_buf4), .Y(_3762_) );
AOI21X1 AOI21X1_622 ( .A(micro_hash_ucr_pipe52_bF_buf1), .B(_2448_), .C(micro_hash_ucr_pipe53_bF_buf1), .Y(_3763_) );
AOI21X1 AOI21X1_623 ( .A(_3763_), .B(_3762_), .C(micro_hash_ucr_pipe54_bF_buf4), .Y(_3764_) );
OAI21X1 OAI21X1_1168 ( .A(_742__bF_buf1), .B(micro_hash_ucr_b_1_bF_buf2_), .C(_2811__bF_buf2), .Y(_3765_) );
OAI21X1 OAI21X1_1169 ( .A(_3764_), .B(_3765_), .C(_832__bF_buf4), .Y(_3766_) );
AOI21X1 AOI21X1_624 ( .A(micro_hash_ucr_pipe56_bF_buf0), .B(_2448_), .C(micro_hash_ucr_pipe57_bF_buf2), .Y(_3767_) );
AOI21X1 AOI21X1_625 ( .A(_3767_), .B(_3766_), .C(micro_hash_ucr_pipe58_bF_buf2), .Y(_3768_) );
OAI21X1 OAI21X1_1170 ( .A(_4211__bF_buf4), .B(micro_hash_ucr_b_1_bF_buf1_), .C(_269_), .Y(_3769_) );
OAI21X1 OAI21X1_1171 ( .A(_3768_), .B(_3769_), .C(_4210__bF_buf0), .Y(_3770_) );
AOI21X1 AOI21X1_626 ( .A(micro_hash_ucr_pipe60_bF_buf3), .B(_2448_), .C(micro_hash_ucr_pipe61_bF_buf0), .Y(_3771_) );
AOI21X1 AOI21X1_627 ( .A(_3771_), .B(_3770_), .C(micro_hash_ucr_pipe62_bF_buf1), .Y(_3772_) );
OAI21X1 OAI21X1_1172 ( .A(_4207__bF_buf2), .B(micro_hash_ucr_b_1_bF_buf0_), .C(_4204_), .Y(_3773_) );
OAI21X1 OAI21X1_1173 ( .A(_3772_), .B(_3773_), .C(_278__bF_buf1), .Y(_3774_) );
AOI21X1 AOI21X1_628 ( .A(micro_hash_ucr_pipe64_bF_buf0), .B(_2448_), .C(micro_hash_ucr_pipe65_bF_buf0), .Y(_3775_) );
AOI21X1 AOI21X1_629 ( .A(_3775_), .B(_3774_), .C(micro_hash_ucr_pipe66_bF_buf2), .Y(_3776_) );
OAI21X1 OAI21X1_1174 ( .A(_1078__bF_buf2), .B(micro_hash_ucr_b_1_bF_buf3_), .C(_4201__bF_buf0), .Y(_3777_) );
OAI21X1 OAI21X1_1175 ( .A(_3776_), .B(_3777_), .C(_4199__bF_buf1), .Y(_3778_) );
OAI21X1 OAI21X1_1176 ( .A(_4199__bF_buf2), .B(micro_hash_ucr_b_1_bF_buf2_), .C(_3778_), .Y(_3779_) );
NOR2X1 NOR2X1_723 ( .A(_345_), .B(_3779_), .Y(_127__1_) );
NOR2X1 NOR2X1_724 ( .A(H_10_), .B(_3668_), .Y(_3780_) );
OAI21X1 OAI21X1_1177 ( .A(_3667_), .B(_3780_), .C(_4239__bF_buf4), .Y(_3781_) );
AOI21X1 AOI21X1_630 ( .A(_4238__bF_buf3), .B(_3781_), .C(micro_hash_ucr_pipe18_bF_buf0), .Y(_3782_) );
OAI21X1 OAI21X1_1178 ( .A(_3668_), .B(_3672_), .C(_2464_), .Y(_3783_) );
NAND2X1 NAND2X1_543 ( .A(_2816_), .B(_3783_), .Y(_3784_) );
OAI21X1 OAI21X1_1179 ( .A(_3782_), .B(_3784_), .C(_4237__bF_buf3), .Y(_3785_) );
AOI21X1 AOI21X1_631 ( .A(micro_hash_ucr_pipe20_bF_buf3), .B(_2464_), .C(micro_hash_ucr_pipe21), .Y(_3786_) );
AOI21X1 AOI21X1_632 ( .A(_3786_), .B(_3785_), .C(micro_hash_ucr_pipe22_bF_buf0), .Y(_3787_) );
OAI21X1 OAI21X1_1180 ( .A(_4262__bF_buf0), .B(micro_hash_ucr_b_2_bF_buf2_), .C(_4234__bF_buf2), .Y(_3788_) );
OAI21X1 OAI21X1_1181 ( .A(_3787_), .B(_3788_), .C(_4233__bF_buf3), .Y(_3789_) );
AOI21X1 AOI21X1_633 ( .A(micro_hash_ucr_pipe24_bF_buf2), .B(_2464_), .C(micro_hash_ucr_pipe25_bF_buf2), .Y(_3790_) );
AOI21X1 AOI21X1_634 ( .A(_3790_), .B(_3789_), .C(micro_hash_ucr_pipe26_bF_buf3), .Y(_3791_) );
OAI21X1 OAI21X1_1182 ( .A(_4230__bF_buf2), .B(micro_hash_ucr_b_2_bF_buf1_), .C(_4229_), .Y(_3792_) );
OAI21X1 OAI21X1_1183 ( .A(_3791_), .B(_3792_), .C(_220__bF_buf1), .Y(_3793_) );
AOI21X1 AOI21X1_635 ( .A(micro_hash_ucr_pipe28_bF_buf2), .B(_2464_), .C(micro_hash_ucr_pipe29), .Y(_3794_) );
AOI21X1 AOI21X1_636 ( .A(_3794_), .B(_3793_), .C(micro_hash_ucr_pipe30_bF_buf0), .Y(_3795_) );
OAI21X1 OAI21X1_1184 ( .A(_4228__bF_buf1), .B(micro_hash_ucr_b_2_bF_buf0_), .C(_317__bF_buf3), .Y(_3796_) );
OAI21X1 OAI21X1_1185 ( .A(_3795_), .B(_3796_), .C(_4226__bF_buf1), .Y(_3797_) );
AOI21X1 AOI21X1_637 ( .A(micro_hash_ucr_pipe32_bF_buf0), .B(_2464_), .C(micro_hash_ucr_pipe33_bF_buf2), .Y(_3798_) );
AOI21X1 AOI21X1_638 ( .A(_3798_), .B(_3797_), .C(micro_hash_ucr_pipe34_bF_buf3), .Y(_3799_) );
OAI21X1 OAI21X1_1186 ( .A(_4225__bF_buf0), .B(micro_hash_ucr_b_2_bF_buf3_), .C(_230__bF_buf2), .Y(_3800_) );
OAI21X1 OAI21X1_1187 ( .A(_3799_), .B(_3800_), .C(_4224__bF_buf2), .Y(_3801_) );
AOI21X1 AOI21X1_639 ( .A(micro_hash_ucr_pipe36_bF_buf0), .B(_2464_), .C(micro_hash_ucr_pipe37_bF_buf1), .Y(_3802_) );
AOI21X1 AOI21X1_640 ( .A(_3802_), .B(_3801_), .C(micro_hash_ucr_pipe38_bF_buf2), .Y(_3803_) );
OAI21X1 OAI21X1_1188 ( .A(_701__bF_buf0), .B(micro_hash_ucr_b_2_bF_buf2_), .C(_2813__bF_buf2), .Y(_3804_) );
OAI21X1 OAI21X1_1189 ( .A(_3803_), .B(_3804_), .C(_296__bF_buf1), .Y(_3805_) );
AOI21X1 AOI21X1_641 ( .A(micro_hash_ucr_pipe40_bF_buf1), .B(_2464_), .C(micro_hash_ucr_pipe41_bF_buf3), .Y(_3806_) );
AOI21X1 AOI21X1_642 ( .A(_3806_), .B(_3805_), .C(micro_hash_ucr_pipe42_bF_buf0), .Y(_3807_) );
OAI21X1 OAI21X1_1190 ( .A(_4220__bF_buf1), .B(micro_hash_ucr_b_2_bF_buf1_), .C(_242__bF_buf2), .Y(_3808_) );
OAI21X1 OAI21X1_1191 ( .A(_3807_), .B(_3808_), .C(_4219__bF_buf3), .Y(_3809_) );
AOI21X1 AOI21X1_643 ( .A(micro_hash_ucr_pipe44_bF_buf0), .B(_2464_), .C(micro_hash_ucr_pipe45), .Y(_3810_) );
AOI21X1 AOI21X1_644 ( .A(_3810_), .B(_3809_), .C(micro_hash_ucr_pipe46_bF_buf3), .Y(_3811_) );
OAI21X1 OAI21X1_1192 ( .A(_4218__bF_buf0), .B(micro_hash_ucr_b_2_bF_buf0_), .C(_249__bF_buf0), .Y(_3812_) );
OAI21X1 OAI21X1_1193 ( .A(_3811_), .B(_3812_), .C(_4217__bF_buf0), .Y(_3813_) );
AOI21X1 AOI21X1_645 ( .A(micro_hash_ucr_pipe48_bF_buf4), .B(_2464_), .C(micro_hash_ucr_pipe49_bF_buf3), .Y(_3814_) );
AOI21X1 AOI21X1_646 ( .A(_3814_), .B(_3813_), .C(micro_hash_ucr_pipe50_bF_buf1), .Y(_3815_) );
OAI21X1 OAI21X1_1194 ( .A(_4215__bF_buf3), .B(micro_hash_ucr_b_2_bF_buf3_), .C(_255__bF_buf3), .Y(_3816_) );
OAI21X1 OAI21X1_1195 ( .A(_3815_), .B(_3816_), .C(_4214__bF_buf1), .Y(_3817_) );
AOI21X1 AOI21X1_647 ( .A(micro_hash_ucr_pipe52_bF_buf1), .B(_2464_), .C(micro_hash_ucr_pipe53_bF_buf1), .Y(_3818_) );
AOI21X1 AOI21X1_648 ( .A(_3818_), .B(_3817_), .C(micro_hash_ucr_pipe54_bF_buf1), .Y(_3819_) );
OAI21X1 OAI21X1_1196 ( .A(_742__bF_buf2), .B(micro_hash_ucr_b_2_bF_buf2_), .C(_2811__bF_buf3), .Y(_3820_) );
OAI21X1 OAI21X1_1197 ( .A(_3819_), .B(_3820_), .C(_832__bF_buf4), .Y(_3821_) );
AOI21X1 AOI21X1_649 ( .A(micro_hash_ucr_pipe56_bF_buf0), .B(_2464_), .C(micro_hash_ucr_pipe57_bF_buf3), .Y(_3822_) );
AOI21X1 AOI21X1_650 ( .A(_3822_), .B(_3821_), .C(micro_hash_ucr_pipe58_bF_buf2), .Y(_3823_) );
OAI21X1 OAI21X1_1198 ( .A(_4211__bF_buf4), .B(micro_hash_ucr_b_2_bF_buf1_), .C(_269_), .Y(_3824_) );
OAI21X1 OAI21X1_1199 ( .A(_3823_), .B(_3824_), .C(_4210__bF_buf0), .Y(_3825_) );
AOI21X1 AOI21X1_651 ( .A(micro_hash_ucr_pipe60_bF_buf3), .B(_2464_), .C(micro_hash_ucr_pipe61_bF_buf0), .Y(_3826_) );
AOI21X1 AOI21X1_652 ( .A(_3826_), .B(_3825_), .C(micro_hash_ucr_pipe62_bF_buf3), .Y(_3827_) );
OAI21X1 OAI21X1_1200 ( .A(_4207__bF_buf2), .B(micro_hash_ucr_b_2_bF_buf0_), .C(_4204_), .Y(_3828_) );
OAI21X1 OAI21X1_1201 ( .A(_3827_), .B(_3828_), .C(_278__bF_buf1), .Y(_3829_) );
AOI21X1 AOI21X1_653 ( .A(micro_hash_ucr_pipe64_bF_buf2), .B(_2464_), .C(micro_hash_ucr_pipe65_bF_buf0), .Y(_3830_) );
AOI21X1 AOI21X1_654 ( .A(_3830_), .B(_3829_), .C(micro_hash_ucr_pipe66_bF_buf2), .Y(_3831_) );
OAI21X1 OAI21X1_1202 ( .A(_1078__bF_buf2), .B(micro_hash_ucr_b_2_bF_buf3_), .C(_4201__bF_buf0), .Y(_3832_) );
OAI21X1 OAI21X1_1203 ( .A(_3831_), .B(_3832_), .C(_4199__bF_buf1), .Y(_3833_) );
OAI21X1 OAI21X1_1204 ( .A(_4199__bF_buf2), .B(micro_hash_ucr_b_2_bF_buf2_), .C(_3833_), .Y(_3834_) );
NOR2X1 NOR2X1_725 ( .A(_345_), .B(_3834_), .Y(_127__2_) );
NOR2X1 NOR2X1_726 ( .A(H_11_), .B(_3668_), .Y(_3835_) );
OAI21X1 OAI21X1_1205 ( .A(_3667_), .B(_3835_), .C(_4239__bF_buf0), .Y(_3836_) );
AOI21X1 AOI21X1_655 ( .A(_4238__bF_buf3), .B(_3836_), .C(micro_hash_ucr_pipe18_bF_buf0), .Y(_3837_) );
OAI21X1 OAI21X1_1206 ( .A(_3668_), .B(_3672_), .C(_2468_), .Y(_3838_) );
NAND2X1 NAND2X1_544 ( .A(_2816_), .B(_3838_), .Y(_3839_) );
OAI21X1 OAI21X1_1207 ( .A(_3837_), .B(_3839_), .C(_4237__bF_buf3), .Y(_3840_) );
AOI21X1 AOI21X1_656 ( .A(micro_hash_ucr_pipe20_bF_buf3), .B(_2468_), .C(micro_hash_ucr_pipe21), .Y(_3841_) );
AOI21X1 AOI21X1_657 ( .A(_3841_), .B(_3840_), .C(micro_hash_ucr_pipe22_bF_buf0), .Y(_3842_) );
OAI21X1 OAI21X1_1208 ( .A(_4262__bF_buf0), .B(micro_hash_ucr_b_3_bF_buf2_), .C(_4234__bF_buf2), .Y(_3843_) );
OAI21X1 OAI21X1_1209 ( .A(_3842_), .B(_3843_), .C(_4233__bF_buf3), .Y(_3844_) );
AOI21X1 AOI21X1_658 ( .A(micro_hash_ucr_pipe24_bF_buf2), .B(_2468_), .C(micro_hash_ucr_pipe25_bF_buf2), .Y(_3845_) );
AOI21X1 AOI21X1_659 ( .A(_3845_), .B(_3844_), .C(micro_hash_ucr_pipe26_bF_buf3), .Y(_3846_) );
OAI21X1 OAI21X1_1210 ( .A(_4230__bF_buf2), .B(micro_hash_ucr_b_3_bF_buf1_), .C(_4229_), .Y(_3847_) );
OAI21X1 OAI21X1_1211 ( .A(_3846_), .B(_3847_), .C(_220__bF_buf1), .Y(_3848_) );
AOI21X1 AOI21X1_660 ( .A(micro_hash_ucr_pipe28_bF_buf2), .B(_2468_), .C(micro_hash_ucr_pipe29), .Y(_3849_) );
AOI21X1 AOI21X1_661 ( .A(_3849_), .B(_3848_), .C(micro_hash_ucr_pipe30_bF_buf3), .Y(_3850_) );
OAI21X1 OAI21X1_1212 ( .A(_4228__bF_buf1), .B(micro_hash_ucr_b_3_bF_buf0_), .C(_317__bF_buf3), .Y(_3851_) );
OAI21X1 OAI21X1_1213 ( .A(_3850_), .B(_3851_), .C(_4226__bF_buf1), .Y(_3852_) );
AOI21X1 AOI21X1_662 ( .A(micro_hash_ucr_pipe32_bF_buf0), .B(_2468_), .C(micro_hash_ucr_pipe33_bF_buf2), .Y(_3853_) );
AOI21X1 AOI21X1_663 ( .A(_3853_), .B(_3852_), .C(micro_hash_ucr_pipe34_bF_buf3), .Y(_3854_) );
OAI21X1 OAI21X1_1214 ( .A(_4225__bF_buf3), .B(micro_hash_ucr_b_3_bF_buf3_), .C(_230__bF_buf0), .Y(_3855_) );
OAI21X1 OAI21X1_1215 ( .A(_3854_), .B(_3855_), .C(_4224__bF_buf0), .Y(_3856_) );
AOI21X1 AOI21X1_664 ( .A(micro_hash_ucr_pipe36_bF_buf0), .B(_2468_), .C(micro_hash_ucr_pipe37_bF_buf2), .Y(_3857_) );
AOI21X1 AOI21X1_665 ( .A(_3857_), .B(_3856_), .C(micro_hash_ucr_pipe38_bF_buf2), .Y(_3858_) );
OAI21X1 OAI21X1_1216 ( .A(_701__bF_buf1), .B(micro_hash_ucr_b_3_bF_buf2_), .C(_2813__bF_buf2), .Y(_3859_) );
OAI21X1 OAI21X1_1217 ( .A(_3858_), .B(_3859_), .C(_296__bF_buf1), .Y(_3860_) );
AOI21X1 AOI21X1_666 ( .A(micro_hash_ucr_pipe40_bF_buf0), .B(_2468_), .C(micro_hash_ucr_pipe41_bF_buf2), .Y(_3861_) );
AOI21X1 AOI21X1_667 ( .A(_3861_), .B(_3860_), .C(micro_hash_ucr_pipe42_bF_buf3), .Y(_3862_) );
OAI21X1 OAI21X1_1218 ( .A(_4220__bF_buf1), .B(micro_hash_ucr_b_3_bF_buf1_), .C(_242__bF_buf3), .Y(_3863_) );
OAI21X1 OAI21X1_1219 ( .A(_3862_), .B(_3863_), .C(_4219__bF_buf3), .Y(_3864_) );
AOI21X1 AOI21X1_668 ( .A(micro_hash_ucr_pipe44_bF_buf0), .B(_2468_), .C(micro_hash_ucr_pipe45), .Y(_3865_) );
AOI21X1 AOI21X1_669 ( .A(_3865_), .B(_3864_), .C(micro_hash_ucr_pipe46_bF_buf3), .Y(_3866_) );
OAI21X1 OAI21X1_1220 ( .A(_4218__bF_buf0), .B(micro_hash_ucr_b_3_bF_buf0_), .C(_249__bF_buf0), .Y(_3867_) );
OAI21X1 OAI21X1_1221 ( .A(_3866_), .B(_3867_), .C(_4217__bF_buf0), .Y(_3868_) );
AOI21X1 AOI21X1_670 ( .A(micro_hash_ucr_pipe48_bF_buf3), .B(_2468_), .C(micro_hash_ucr_pipe49_bF_buf3), .Y(_3869_) );
AOI21X1 AOI21X1_671 ( .A(_3869_), .B(_3868_), .C(micro_hash_ucr_pipe50_bF_buf1), .Y(_3870_) );
OAI21X1 OAI21X1_1222 ( .A(_4215__bF_buf0), .B(micro_hash_ucr_b_3_bF_buf3_), .C(_255__bF_buf1), .Y(_3871_) );
OAI21X1 OAI21X1_1223 ( .A(_3870_), .B(_3871_), .C(_4214__bF_buf4), .Y(_3872_) );
AOI21X1 AOI21X1_672 ( .A(micro_hash_ucr_pipe52_bF_buf1), .B(_2468_), .C(micro_hash_ucr_pipe53_bF_buf1), .Y(_3873_) );
AOI21X1 AOI21X1_673 ( .A(_3873_), .B(_3872_), .C(micro_hash_ucr_pipe54_bF_buf1), .Y(_3874_) );
OAI21X1 OAI21X1_1224 ( .A(_742__bF_buf2), .B(micro_hash_ucr_b_3_bF_buf2_), .C(_2811__bF_buf3), .Y(_3875_) );
OAI21X1 OAI21X1_1225 ( .A(_3874_), .B(_3875_), .C(_832__bF_buf4), .Y(_3876_) );
AOI21X1 AOI21X1_674 ( .A(micro_hash_ucr_pipe56_bF_buf0), .B(_2468_), .C(micro_hash_ucr_pipe57_bF_buf3), .Y(_3877_) );
AOI21X1 AOI21X1_675 ( .A(_3877_), .B(_3876_), .C(micro_hash_ucr_pipe58_bF_buf2), .Y(_3878_) );
OAI21X1 OAI21X1_1226 ( .A(_4211__bF_buf4), .B(micro_hash_ucr_b_3_bF_buf1_), .C(_269_), .Y(_3879_) );
OAI21X1 OAI21X1_1227 ( .A(_3878_), .B(_3879_), .C(_4210__bF_buf0), .Y(_3880_) );
AOI21X1 AOI21X1_676 ( .A(micro_hash_ucr_pipe60_bF_buf3), .B(_2468_), .C(micro_hash_ucr_pipe61_bF_buf1), .Y(_3881_) );
AOI21X1 AOI21X1_677 ( .A(_3881_), .B(_3880_), .C(micro_hash_ucr_pipe62_bF_buf3), .Y(_3882_) );
OAI21X1 OAI21X1_1228 ( .A(_4207__bF_buf3), .B(micro_hash_ucr_b_3_bF_buf0_), .C(_4204_), .Y(_3883_) );
OAI21X1 OAI21X1_1229 ( .A(_3882_), .B(_3883_), .C(_278__bF_buf1), .Y(_3884_) );
AOI21X1 AOI21X1_678 ( .A(micro_hash_ucr_pipe64_bF_buf2), .B(_2468_), .C(micro_hash_ucr_pipe65_bF_buf0), .Y(_3885_) );
AOI21X1 AOI21X1_679 ( .A(_3885_), .B(_3884_), .C(micro_hash_ucr_pipe66_bF_buf2), .Y(_3886_) );
OAI21X1 OAI21X1_1230 ( .A(_1078__bF_buf2), .B(micro_hash_ucr_b_3_bF_buf3_), .C(_4201__bF_buf0), .Y(_3887_) );
OAI21X1 OAI21X1_1231 ( .A(_3886_), .B(_3887_), .C(_4199__bF_buf1), .Y(_3888_) );
OAI21X1 OAI21X1_1232 ( .A(_4199__bF_buf1), .B(micro_hash_ucr_b_3_bF_buf2_), .C(_3888_), .Y(_3889_) );
NOR2X1 NOR2X1_727 ( .A(_345_), .B(_3889_), .Y(_127__3_) );
NAND2X1 NAND2X1_545 ( .A(micro_hash_ucr_pipe63_bF_buf3), .B(micro_hash_ucr_c_0_bF_buf3_), .Y(_3890_) );
NAND2X1 NAND2X1_546 ( .A(micro_hash_ucr_pipe61_bF_buf0), .B(micro_hash_ucr_c_0_bF_buf2_), .Y(_3891_) );
INVX8 INVX8_92 ( .A(micro_hash_ucr_b_4_), .Y(_3892_) );
NAND2X1 NAND2X1_547 ( .A(micro_hash_ucr_pipe56_bF_buf2), .B(_3892__bF_buf2), .Y(_3893_) );
NAND2X1 NAND2X1_548 ( .A(micro_hash_ucr_pipe55), .B(micro_hash_ucr_c_0_bF_buf1_), .Y(_3894_) );
NOR2X1 NOR2X1_728 ( .A(_742__bF_buf1), .B(_3892__bF_buf2), .Y(_3895_) );
NAND2X1 NAND2X1_549 ( .A(micro_hash_ucr_pipe53_bF_buf0), .B(micro_hash_ucr_c_0_bF_buf0_), .Y(_3896_) );
NAND2X1 NAND2X1_550 ( .A(micro_hash_ucr_pipe52_bF_buf0), .B(micro_hash_ucr_b_4_), .Y(_3897_) );
NAND2X1 NAND2X1_551 ( .A(micro_hash_ucr_pipe36_bF_buf3), .B(_3892__bF_buf1), .Y(_3898_) );
NAND2X1 NAND2X1_552 ( .A(micro_hash_ucr_pipe35), .B(micro_hash_ucr_c_0_bF_buf3_), .Y(_3899_) );
NAND2X1 NAND2X1_553 ( .A(micro_hash_ucr_pipe34_bF_buf1), .B(_3892__bF_buf1), .Y(_3900_) );
NAND2X1 NAND2X1_554 ( .A(micro_hash_ucr_pipe33_bF_buf1), .B(micro_hash_ucr_c_0_bF_buf2_), .Y(_3901_) );
NAND2X1 NAND2X1_555 ( .A(micro_hash_ucr_b_4_), .B(micro_hash_ucr_pipe24_bF_buf0), .Y(_3902_) );
NAND2X1 NAND2X1_556 ( .A(micro_hash_ucr_pipe23), .B(_2391_), .Y(_3903_) );
NAND2X1 NAND2X1_557 ( .A(micro_hash_ucr_pipe19), .B(micro_hash_ucr_c_0_bF_buf1_), .Y(_3904_) );
NAND2X1 NAND2X1_558 ( .A(micro_hash_ucr_pipe18_bF_buf1), .B(_3892__bF_buf0), .Y(_3905_) );
NAND2X1 NAND2X1_559 ( .A(micro_hash_ucr_pipe17), .B(micro_hash_ucr_c_0_bF_buf0_), .Y(_3906_) );
NAND2X1 NAND2X1_560 ( .A(micro_hash_ucr_pipe16), .B(_3892__bF_buf0), .Y(_3907_) );
NAND2X1 NAND2X1_561 ( .A(micro_hash_ucr_pipe15), .B(micro_hash_ucr_c_0_bF_buf3_), .Y(_3908_) );
NOR2X1 NOR2X1_729 ( .A(_2391_), .B(_4279_), .Y(_3909_) );
NOR2X1 NOR2X1_730 ( .A(micro_hash_ucr_b_4_), .B(_4260_), .Y(_3910_) );
NAND2X1 NAND2X1_562 ( .A(micro_hash_ucr_b_4_), .B(_4246_), .Y(_3911_) );
OAI21X1 OAI21X1_1233 ( .A(_2925_), .B(micro_hash_ucr_pipe13), .C(_2391_), .Y(_3912_) );
NAND3X1 NAND3X1_214 ( .A(_4255_), .B(_2479_), .C(_2823_), .Y(_3913_) );
NAND2X1 NAND2X1_563 ( .A(_3913_), .B(_3912_), .Y(_3914_) );
AOI21X1 AOI21X1_680 ( .A(_3911_), .B(_3914_), .C(_3910_), .Y(_3915_) );
OAI21X1 OAI21X1_1234 ( .A(_3915_), .B(_3909_), .C(_4240_), .Y(_3916_) );
NAND3X1 NAND3X1_215 ( .A(_4239__bF_buf3), .B(_3908_), .C(_3916_), .Y(_3917_) );
NAND3X1 NAND3X1_216 ( .A(_4238__bF_buf2), .B(_3907_), .C(_3917_), .Y(_3918_) );
NAND3X1 NAND3X1_217 ( .A(_624__bF_buf1), .B(_3906_), .C(_3918_), .Y(_3919_) );
NAND3X1 NAND3X1_218 ( .A(_2816_), .B(_3905_), .C(_3919_), .Y(_3920_) );
AOI21X1 AOI21X1_681 ( .A(_3904_), .B(_3920_), .C(micro_hash_ucr_pipe20_bF_buf2), .Y(_3921_) );
OAI21X1 OAI21X1_1235 ( .A(_3892__bF_buf0), .B(_4237__bF_buf0), .C(_4236__bF_buf2), .Y(_3922_) );
AOI21X1 AOI21X1_682 ( .A(micro_hash_ucr_pipe21), .B(_2391_), .C(micro_hash_ucr_pipe22_bF_buf2), .Y(_3923_) );
OAI21X1 OAI21X1_1236 ( .A(_3921_), .B(_3922_), .C(_3923_), .Y(_3924_) );
NAND2X1 NAND2X1_564 ( .A(micro_hash_ucr_b_4_), .B(micro_hash_ucr_pipe22_bF_buf3), .Y(_3925_) );
NAND3X1 NAND3X1_219 ( .A(_4234__bF_buf3), .B(_3925_), .C(_3924_), .Y(_3926_) );
NAND3X1 NAND3X1_220 ( .A(_4233__bF_buf4), .B(_3903_), .C(_3926_), .Y(_3927_) );
AOI21X1 AOI21X1_683 ( .A(_3902_), .B(_3927_), .C(micro_hash_ucr_pipe25_bF_buf1), .Y(_3928_) );
OAI21X1 OAI21X1_1237 ( .A(_389__bF_buf3), .B(_2391_), .C(_4230__bF_buf4), .Y(_3929_) );
AOI21X1 AOI21X1_684 ( .A(micro_hash_ucr_pipe26_bF_buf2), .B(_3892__bF_buf3), .C(micro_hash_ucr_pipe27_bF_buf2), .Y(_3930_) );
OAI21X1 OAI21X1_1238 ( .A(_3928_), .B(_3929_), .C(_3930_), .Y(_3931_) );
AOI21X1 AOI21X1_685 ( .A(micro_hash_ucr_pipe27_bF_buf3), .B(micro_hash_ucr_c_0_bF_buf2_), .C(micro_hash_ucr_pipe28_bF_buf2), .Y(_3932_) );
AOI22X1 AOI22X1_30 ( .A(_3892__bF_buf3), .B(micro_hash_ucr_pipe28_bF_buf1), .C(_3931_), .D(_3932_), .Y(_3933_) );
OAI21X1 OAI21X1_1239 ( .A(_219_), .B(_2391_), .C(_4228__bF_buf0), .Y(_3934_) );
AOI21X1 AOI21X1_686 ( .A(_219_), .B(_3933_), .C(_3934_), .Y(_3935_) );
OAI21X1 OAI21X1_1240 ( .A(_4228__bF_buf0), .B(micro_hash_ucr_b_4_), .C(_317__bF_buf0), .Y(_3936_) );
AOI21X1 AOI21X1_687 ( .A(micro_hash_ucr_pipe31_bF_buf0), .B(micro_hash_ucr_c_0_bF_buf1_), .C(micro_hash_ucr_pipe32_bF_buf1), .Y(_3937_) );
OAI21X1 OAI21X1_1241 ( .A(_3935_), .B(_3936_), .C(_3937_), .Y(_3938_) );
NAND2X1 NAND2X1_565 ( .A(micro_hash_ucr_pipe32_bF_buf1), .B(_3892__bF_buf3), .Y(_3939_) );
NAND3X1 NAND3X1_221 ( .A(_318_), .B(_3939_), .C(_3938_), .Y(_3940_) );
NAND3X1 NAND3X1_222 ( .A(_4225__bF_buf1), .B(_3901_), .C(_3940_), .Y(_3941_) );
NAND3X1 NAND3X1_223 ( .A(_230__bF_buf1), .B(_3900_), .C(_3941_), .Y(_3942_) );
NAND3X1 NAND3X1_224 ( .A(_4224__bF_buf3), .B(_3899_), .C(_3942_), .Y(_3943_) );
NAND3X1 NAND3X1_225 ( .A(_2815_), .B(_3898_), .C(_3943_), .Y(_3944_) );
AOI21X1 AOI21X1_688 ( .A(micro_hash_ucr_pipe37_bF_buf3), .B(micro_hash_ucr_c_0_bF_buf0_), .C(micro_hash_ucr_pipe38_bF_buf0), .Y(_3945_) );
OAI21X1 OAI21X1_1242 ( .A(_701__bF_buf1), .B(micro_hash_ucr_b_4_), .C(_2813__bF_buf1), .Y(_3946_) );
AOI21X1 AOI21X1_689 ( .A(_3945_), .B(_3944_), .C(_3946_), .Y(_3947_) );
OAI21X1 OAI21X1_1243 ( .A(_2813__bF_buf1), .B(_2391_), .C(_296__bF_buf3), .Y(_3948_) );
NAND2X1 NAND2X1_566 ( .A(micro_hash_ucr_pipe40_bF_buf3), .B(_3892__bF_buf1), .Y(_3949_) );
OAI21X1 OAI21X1_1244 ( .A(_3947_), .B(_3948_), .C(_3949_), .Y(_3950_) );
NAND2X1 NAND2X1_567 ( .A(micro_hash_ucr_pipe41_bF_buf0), .B(micro_hash_ucr_c_0_bF_buf3_), .Y(_3951_) );
OAI21X1 OAI21X1_1245 ( .A(_3950_), .B(micro_hash_ucr_pipe41_bF_buf0), .C(_3951_), .Y(_3952_) );
AOI21X1 AOI21X1_690 ( .A(micro_hash_ucr_pipe42_bF_buf1), .B(_3892__bF_buf1), .C(micro_hash_ucr_pipe43), .Y(_3953_) );
OAI21X1 OAI21X1_1246 ( .A(_3952_), .B(micro_hash_ucr_pipe42_bF_buf1), .C(_3953_), .Y(_3954_) );
AOI21X1 AOI21X1_691 ( .A(micro_hash_ucr_pipe43), .B(micro_hash_ucr_c_0_bF_buf2_), .C(micro_hash_ucr_pipe44_bF_buf2), .Y(_3955_) );
AOI22X1 AOI22X1_31 ( .A(micro_hash_ucr_pipe44_bF_buf2), .B(_3892__bF_buf1), .C(_3954_), .D(_3955_), .Y(_3956_) );
NAND2X1 NAND2X1_568 ( .A(_336_), .B(_3956_), .Y(_3957_) );
OAI21X1 OAI21X1_1247 ( .A(_336_), .B(_2391_), .C(_3957_), .Y(_3958_) );
AOI21X1 AOI21X1_692 ( .A(micro_hash_ucr_pipe46_bF_buf4), .B(_3892__bF_buf2), .C(micro_hash_ucr_pipe47), .Y(_3959_) );
OAI21X1 OAI21X1_1248 ( .A(_3958_), .B(micro_hash_ucr_pipe46_bF_buf4), .C(_3959_), .Y(_3960_) );
OAI21X1 OAI21X1_1249 ( .A(_249__bF_buf3), .B(_2391_), .C(_3960_), .Y(_3961_) );
NAND2X1 NAND2X1_569 ( .A(_4217__bF_buf3), .B(_3961_), .Y(_3962_) );
OAI21X1 OAI21X1_1250 ( .A(_4217__bF_buf3), .B(_3892__bF_buf2), .C(_3962_), .Y(_3963_) );
NOR2X1 NOR2X1_731 ( .A(micro_hash_ucr_pipe49_bF_buf2), .B(_3963_), .Y(_3964_) );
OAI21X1 OAI21X1_1251 ( .A(_304_), .B(micro_hash_ucr_c_0_bF_buf1_), .C(_4215__bF_buf2), .Y(_3965_) );
OAI22X1 OAI22X1_47 ( .A(_4215__bF_buf1), .B(_3892__bF_buf2), .C(_3964_), .D(_3965_), .Y(_3966_) );
NAND2X1 NAND2X1_570 ( .A(micro_hash_ucr_pipe51), .B(_2391_), .Y(_3967_) );
OAI21X1 OAI21X1_1252 ( .A(_3966_), .B(micro_hash_ucr_pipe51), .C(_3967_), .Y(_3968_) );
OAI21X1 OAI21X1_1253 ( .A(_3968_), .B(micro_hash_ucr_pipe52_bF_buf0), .C(_3897_), .Y(_3969_) );
NAND2X1 NAND2X1_571 ( .A(_2812_), .B(_3969_), .Y(_3970_) );
AOI21X1 AOI21X1_693 ( .A(_3896_), .B(_3970_), .C(micro_hash_ucr_pipe54_bF_buf4), .Y(_3971_) );
OAI21X1 OAI21X1_1254 ( .A(_3971_), .B(_3895_), .C(_2811__bF_buf0), .Y(_3972_) );
NAND3X1 NAND3X1_226 ( .A(_832__bF_buf2), .B(_3894_), .C(_3972_), .Y(_3973_) );
NAND3X1 NAND3X1_227 ( .A(_4212_), .B(_3893_), .C(_3973_), .Y(_3974_) );
AOI21X1 AOI21X1_694 ( .A(micro_hash_ucr_pipe57_bF_buf1), .B(micro_hash_ucr_c_0_bF_buf0_), .C(micro_hash_ucr_pipe58_bF_buf3), .Y(_3975_) );
OAI21X1 OAI21X1_1255 ( .A(_4211__bF_buf0), .B(micro_hash_ucr_b_4_), .C(_269_), .Y(_3976_) );
AOI21X1 AOI21X1_695 ( .A(_3975_), .B(_3974_), .C(_3976_), .Y(_3977_) );
OAI21X1 OAI21X1_1256 ( .A(_269_), .B(_2391_), .C(_4210__bF_buf3), .Y(_3978_) );
OAI22X1 OAI22X1_48 ( .A(_4210__bF_buf3), .B(micro_hash_ucr_b_4_), .C(_3977_), .D(_3978_), .Y(_3979_) );
OAI21X1 OAI21X1_1257 ( .A(_3979_), .B(micro_hash_ucr_pipe61_bF_buf0), .C(_3891_), .Y(_3980_) );
NAND2X1 NAND2X1_572 ( .A(micro_hash_ucr_pipe62_bF_buf2), .B(_3892__bF_buf3), .Y(_3981_) );
OAI21X1 OAI21X1_1258 ( .A(_3980_), .B(micro_hash_ucr_pipe62_bF_buf2), .C(_3981_), .Y(_3982_) );
OAI21X1 OAI21X1_1259 ( .A(_3982_), .B(micro_hash_ucr_pipe63_bF_buf3), .C(_3890_), .Y(_3983_) );
NAND2X1 NAND2X1_573 ( .A(micro_hash_ucr_pipe64_bF_buf0), .B(_3892__bF_buf3), .Y(_3984_) );
OAI21X1 OAI21X1_1260 ( .A(_3983_), .B(micro_hash_ucr_pipe64_bF_buf1), .C(_3984_), .Y(_3985_) );
AOI21X1 AOI21X1_696 ( .A(micro_hash_ucr_pipe65_bF_buf4), .B(micro_hash_ucr_c_0_bF_buf3_), .C(micro_hash_ucr_pipe66_bF_buf0), .Y(_3986_) );
OAI21X1 OAI21X1_1261 ( .A(_3985_), .B(micro_hash_ucr_pipe65_bF_buf4), .C(_3986_), .Y(_3987_) );
AOI21X1 AOI21X1_697 ( .A(micro_hash_ucr_pipe66_bF_buf0), .B(_3892__bF_buf0), .C(micro_hash_ucr_pipe67), .Y(_3988_) );
OAI21X1 OAI21X1_1262 ( .A(_4201__bF_buf0), .B(_2391_), .C(_4199__bF_buf4), .Y(_3989_) );
AOI21X1 AOI21X1_698 ( .A(_3988_), .B(_3987_), .C(_3989_), .Y(_3990_) );
OAI21X1 OAI21X1_1263 ( .A(_4199__bF_buf0), .B(micro_hash_ucr_b_4_), .C(_344_), .Y(_3991_) );
OAI22X1 OAI22X1_49 ( .A(_2391_), .B(_2181_), .C(_3990_), .D(_3991_), .Y(_127__4_) );
NAND2X1 NAND2X1_574 ( .A(micro_hash_ucr_c_1_bF_buf0_), .B(_198_), .Y(_3992_) );
NAND2X1 NAND2X1_575 ( .A(micro_hash_ucr_pipe63_bF_buf2), .B(micro_hash_ucr_c_1_bF_buf3_), .Y(_3993_) );
NAND2X1 NAND2X1_576 ( .A(micro_hash_ucr_pipe62_bF_buf1), .B(_2487__bF_buf0), .Y(_3994_) );
NAND2X1 NAND2X1_577 ( .A(micro_hash_ucr_pipe61_bF_buf1), .B(micro_hash_ucr_c_1_bF_buf2_), .Y(_3995_) );
NAND2X1 NAND2X1_578 ( .A(micro_hash_ucr_pipe57_bF_buf3), .B(_591__bF_buf1), .Y(_3996_) );
NAND2X1 NAND2X1_579 ( .A(micro_hash_ucr_pipe52_bF_buf1), .B(_2487__bF_buf3), .Y(_3997_) );
NOR2X1 NOR2X1_732 ( .A(micro_hash_ucr_c_1_bF_buf1_), .B(_255__bF_buf2), .Y(_3998_) );
NAND2X1 NAND2X1_580 ( .A(micro_hash_ucr_pipe50_bF_buf1), .B(_2487__bF_buf3), .Y(_3999_) );
NOR2X1 NOR2X1_733 ( .A(micro_hash_ucr_c_1_bF_buf0_), .B(_304_), .Y(_4000_) );
NAND2X1 NAND2X1_581 ( .A(micro_hash_ucr_pipe37_bF_buf0), .B(micro_hash_ucr_c_1_bF_buf3_), .Y(_4001_) );
NAND2X1 NAND2X1_582 ( .A(micro_hash_ucr_b_5_bF_buf2_), .B(micro_hash_ucr_pipe32_bF_buf2), .Y(_4002_) );
NAND2X1 NAND2X1_583 ( .A(micro_hash_ucr_b_5_bF_buf1_), .B(micro_hash_ucr_pipe20_bF_buf2), .Y(_4003_) );
NAND2X1 NAND2X1_584 ( .A(micro_hash_ucr_b_5_bF_buf0_), .B(micro_hash_ucr_pipe14), .Y(_4004_) );
OAI21X1 OAI21X1_1264 ( .A(_4257_), .B(micro_hash_ucr_pipe12_bF_buf1), .C(_2487__bF_buf1), .Y(_4005_) );
NOR2X1 NOR2X1_734 ( .A(micro_hash_ucr_pipe13), .B(_3152_), .Y(_4006_) );
NAND2X1 NAND2X1_585 ( .A(_4242_), .B(_4272_), .Y(_4007_) );
NOR2X1 NOR2X1_735 ( .A(H_13_), .B(_4266_), .Y(_4008_) );
AOI22X1 AOI22X1_32 ( .A(_4253_), .B(_4008_), .C(_4007_), .D(_591__bF_buf3), .Y(_4009_) );
OAI21X1 OAI21X1_1265 ( .A(_4009_), .B(_4006_), .C(_4005_), .Y(_4010_) );
NOR2X1 NOR2X1_736 ( .A(micro_hash_ucr_pipe13), .B(_2487__bF_buf1), .Y(_4011_) );
AOI22X1 AOI22X1_33 ( .A(micro_hash_ucr_pipe12_bF_buf1), .B(_4011_), .C(_4278_), .D(micro_hash_ucr_c_1_bF_buf2_), .Y(_4012_) );
AND2X2 AND2X2_266 ( .A(_4010_), .B(_4012_), .Y(_4013_) );
OAI21X1 OAI21X1_1266 ( .A(_4013_), .B(micro_hash_ucr_pipe14), .C(_4004_), .Y(_4014_) );
NAND2X1 NAND2X1_586 ( .A(micro_hash_ucr_pipe15), .B(_591__bF_buf3), .Y(_4015_) );
OAI21X1 OAI21X1_1267 ( .A(_4014_), .B(micro_hash_ucr_pipe15), .C(_4015_), .Y(_4016_) );
OAI21X1 OAI21X1_1268 ( .A(_4239__bF_buf1), .B(micro_hash_ucr_b_5_bF_buf3_), .C(_4238__bF_buf0), .Y(_4017_) );
AOI21X1 AOI21X1_699 ( .A(_4239__bF_buf1), .B(_4016_), .C(_4017_), .Y(_4018_) );
OAI21X1 OAI21X1_1269 ( .A(_4238__bF_buf0), .B(_591__bF_buf2), .C(_624__bF_buf2), .Y(_4019_) );
OAI22X1 OAI22X1_50 ( .A(micro_hash_ucr_b_5_bF_buf2_), .B(_624__bF_buf2), .C(_4018_), .D(_4019_), .Y(_4020_) );
NAND2X1 NAND2X1_587 ( .A(_2816_), .B(_4020_), .Y(_4021_) );
OAI21X1 OAI21X1_1270 ( .A(_2816_), .B(micro_hash_ucr_c_1_bF_buf1_), .C(_4021_), .Y(_4022_) );
OAI21X1 OAI21X1_1271 ( .A(_4022_), .B(micro_hash_ucr_pipe20_bF_buf2), .C(_4003_), .Y(_4023_) );
NAND2X1 NAND2X1_588 ( .A(_4236__bF_buf3), .B(_4023_), .Y(_4024_) );
OAI21X1 OAI21X1_1272 ( .A(_4236__bF_buf3), .B(_591__bF_buf2), .C(_4024_), .Y(_4025_) );
AOI21X1 AOI21X1_700 ( .A(micro_hash_ucr_pipe22_bF_buf2), .B(_2487__bF_buf1), .C(micro_hash_ucr_pipe23), .Y(_4026_) );
OAI21X1 OAI21X1_1273 ( .A(_4025_), .B(micro_hash_ucr_pipe22_bF_buf2), .C(_4026_), .Y(_4027_) );
OAI21X1 OAI21X1_1274 ( .A(_4234__bF_buf1), .B(_591__bF_buf2), .C(_4027_), .Y(_4028_) );
NAND2X1 NAND2X1_589 ( .A(_4233__bF_buf2), .B(_4028_), .Y(_4029_) );
OAI21X1 OAI21X1_1275 ( .A(_2487__bF_buf2), .B(_4233__bF_buf2), .C(_4029_), .Y(_4030_) );
OAI21X1 OAI21X1_1276 ( .A(_389__bF_buf0), .B(_591__bF_buf2), .C(_4230__bF_buf0), .Y(_4031_) );
AOI21X1 AOI21X1_701 ( .A(_389__bF_buf0), .B(_4030_), .C(_4031_), .Y(_4032_) );
OAI21X1 OAI21X1_1277 ( .A(_4230__bF_buf2), .B(micro_hash_ucr_b_5_bF_buf1_), .C(_4229_), .Y(_4033_) );
OAI22X1 OAI22X1_51 ( .A(_4229_), .B(_591__bF_buf0), .C(_4032_), .D(_4033_), .Y(_4034_) );
OAI21X1 OAI21X1_1278 ( .A(_2487__bF_buf2), .B(_220__bF_buf4), .C(_219_), .Y(_4035_) );
AOI21X1 AOI21X1_702 ( .A(_220__bF_buf4), .B(_4034_), .C(_4035_), .Y(_4036_) );
OAI21X1 OAI21X1_1279 ( .A(_219_), .B(micro_hash_ucr_c_1_bF_buf0_), .C(_4228__bF_buf2), .Y(_4037_) );
OAI22X1 OAI22X1_52 ( .A(_2487__bF_buf2), .B(_4228__bF_buf2), .C(_4036_), .D(_4037_), .Y(_4038_) );
NAND2X1 NAND2X1_590 ( .A(micro_hash_ucr_pipe31_bF_buf3), .B(_591__bF_buf0), .Y(_4039_) );
OAI21X1 OAI21X1_1280 ( .A(_4038_), .B(micro_hash_ucr_pipe31_bF_buf1), .C(_4039_), .Y(_4040_) );
OAI21X1 OAI21X1_1281 ( .A(_4040_), .B(micro_hash_ucr_pipe32_bF_buf2), .C(_4002_), .Y(_4041_) );
OAI21X1 OAI21X1_1282 ( .A(_318_), .B(_591__bF_buf0), .C(_4225__bF_buf2), .Y(_4042_) );
AOI21X1 AOI21X1_703 ( .A(_318_), .B(_4041_), .C(_4042_), .Y(_4043_) );
OAI21X1 OAI21X1_1283 ( .A(_4225__bF_buf3), .B(micro_hash_ucr_b_5_bF_buf0_), .C(_230__bF_buf3), .Y(_4044_) );
AOI21X1 AOI21X1_704 ( .A(micro_hash_ucr_pipe35), .B(micro_hash_ucr_c_1_bF_buf3_), .C(micro_hash_ucr_pipe36_bF_buf2), .Y(_4045_) );
OAI21X1 OAI21X1_1284 ( .A(_4043_), .B(_4044_), .C(_4045_), .Y(_4046_) );
NAND2X1 NAND2X1_591 ( .A(micro_hash_ucr_pipe36_bF_buf2), .B(_2487__bF_buf0), .Y(_4047_) );
NAND3X1 NAND3X1_228 ( .A(_2815_), .B(_4047_), .C(_4046_), .Y(_4048_) );
AOI21X1 AOI21X1_705 ( .A(_4001_), .B(_4048_), .C(micro_hash_ucr_pipe38_bF_buf1), .Y(_4049_) );
OAI21X1 OAI21X1_1285 ( .A(_2487__bF_buf0), .B(_701__bF_buf3), .C(_2813__bF_buf3), .Y(_4050_) );
AOI21X1 AOI21X1_706 ( .A(micro_hash_ucr_pipe39), .B(_591__bF_buf1), .C(micro_hash_ucr_pipe40_bF_buf2), .Y(_4051_) );
OAI21X1 OAI21X1_1286 ( .A(_4049_), .B(_4050_), .C(_4051_), .Y(_4052_) );
NAND2X1 NAND2X1_592 ( .A(micro_hash_ucr_pipe40_bF_buf2), .B(micro_hash_ucr_b_5_bF_buf3_), .Y(_4053_) );
AOI21X1 AOI21X1_707 ( .A(_4053_), .B(_4052_), .C(micro_hash_ucr_pipe41_bF_buf1), .Y(_4054_) );
OAI21X1 OAI21X1_1287 ( .A(_2814_), .B(_591__bF_buf1), .C(_4220__bF_buf3), .Y(_4055_) );
AOI21X1 AOI21X1_708 ( .A(micro_hash_ucr_pipe42_bF_buf3), .B(_2487__bF_buf3), .C(micro_hash_ucr_pipe43), .Y(_4056_) );
OAI21X1 OAI21X1_1288 ( .A(_4054_), .B(_4055_), .C(_4056_), .Y(_4057_) );
AOI21X1 AOI21X1_709 ( .A(micro_hash_ucr_pipe43), .B(micro_hash_ucr_c_1_bF_buf2_), .C(micro_hash_ucr_pipe44_bF_buf3), .Y(_4058_) );
AOI22X1 AOI22X1_34 ( .A(micro_hash_ucr_pipe44_bF_buf3), .B(_2487__bF_buf3), .C(_4057_), .D(_4058_), .Y(_4059_) );
OAI21X1 OAI21X1_1289 ( .A(_336_), .B(_591__bF_buf1), .C(_4218__bF_buf0), .Y(_4060_) );
AOI21X1 AOI21X1_710 ( .A(_336_), .B(_4059_), .C(_4060_), .Y(_4061_) );
OAI21X1 OAI21X1_1290 ( .A(_4218__bF_buf0), .B(micro_hash_ucr_b_5_bF_buf2_), .C(_249__bF_buf0), .Y(_4062_) );
AOI21X1 AOI21X1_711 ( .A(micro_hash_ucr_pipe47), .B(micro_hash_ucr_c_1_bF_buf1_), .C(micro_hash_ucr_pipe48_bF_buf4), .Y(_4063_) );
OAI21X1 OAI21X1_1291 ( .A(_4061_), .B(_4062_), .C(_4063_), .Y(_4064_) );
NAND2X1 NAND2X1_593 ( .A(micro_hash_ucr_pipe48_bF_buf4), .B(_2487__bF_buf3), .Y(_4065_) );
AOI21X1 AOI21X1_712 ( .A(_4065_), .B(_4064_), .C(micro_hash_ucr_pipe49_bF_buf3), .Y(_4066_) );
OAI21X1 OAI21X1_1292 ( .A(_4066_), .B(_4000_), .C(_4215__bF_buf3), .Y(_4067_) );
AOI21X1 AOI21X1_713 ( .A(_3999_), .B(_4067_), .C(micro_hash_ucr_pipe51), .Y(_4068_) );
OAI21X1 OAI21X1_1293 ( .A(_4068_), .B(_3998_), .C(_4214__bF_buf4), .Y(_4069_) );
NAND3X1 NAND3X1_229 ( .A(_2812_), .B(_3997_), .C(_4069_), .Y(_4070_) );
AOI21X1 AOI21X1_714 ( .A(micro_hash_ucr_pipe53_bF_buf2), .B(micro_hash_ucr_c_1_bF_buf0_), .C(micro_hash_ucr_pipe54_bF_buf1), .Y(_4071_) );
OAI21X1 OAI21X1_1294 ( .A(_742__bF_buf2), .B(micro_hash_ucr_b_5_bF_buf1_), .C(_2811__bF_buf3), .Y(_4072_) );
AOI21X1 AOI21X1_715 ( .A(_4071_), .B(_4070_), .C(_4072_), .Y(_4073_) );
OAI21X1 OAI21X1_1295 ( .A(_2811__bF_buf3), .B(_591__bF_buf1), .C(_832__bF_buf1), .Y(_4074_) );
OAI22X1 OAI22X1_53 ( .A(_832__bF_buf1), .B(micro_hash_ucr_b_5_bF_buf0_), .C(_4073_), .D(_4074_), .Y(_4075_) );
NAND2X1 NAND2X1_594 ( .A(_4212_), .B(_4075_), .Y(_4076_) );
NAND3X1 NAND3X1_230 ( .A(_4211__bF_buf4), .B(_3996_), .C(_4076_), .Y(_4077_) );
AOI21X1 AOI21X1_716 ( .A(micro_hash_ucr_pipe58_bF_buf2), .B(micro_hash_ucr_b_5_bF_buf3_), .C(micro_hash_ucr_pipe59), .Y(_4078_) );
OAI21X1 OAI21X1_1296 ( .A(_269_), .B(micro_hash_ucr_c_1_bF_buf3_), .C(_4210__bF_buf0), .Y(_4079_) );
AOI21X1 AOI21X1_717 ( .A(_4078_), .B(_4077_), .C(_4079_), .Y(_4080_) );
NOR2X1 NOR2X1_737 ( .A(_4210__bF_buf0), .B(_2487__bF_buf0), .Y(_4081_) );
OAI21X1 OAI21X1_1297 ( .A(_4080_), .B(_4081_), .C(_4208_), .Y(_4082_) );
NAND3X1 NAND3X1_231 ( .A(_4207__bF_buf3), .B(_3995_), .C(_4082_), .Y(_4083_) );
NAND3X1 NAND3X1_232 ( .A(_4204_), .B(_3994_), .C(_4083_), .Y(_4084_) );
NAND3X1 NAND3X1_233 ( .A(_278__bF_buf1), .B(_3993_), .C(_4084_), .Y(_4085_) );
OAI21X1 OAI21X1_1298 ( .A(_278__bF_buf2), .B(micro_hash_ucr_b_5_bF_buf2_), .C(_4085_), .Y(_4086_) );
AOI21X1 AOI21X1_718 ( .A(micro_hash_ucr_pipe65_bF_buf3), .B(micro_hash_ucr_c_1_bF_buf2_), .C(micro_hash_ucr_pipe66_bF_buf2), .Y(_4087_) );
OAI21X1 OAI21X1_1299 ( .A(_4086_), .B(micro_hash_ucr_pipe65_bF_buf3), .C(_4087_), .Y(_4088_) );
AOI21X1 AOI21X1_719 ( .A(micro_hash_ucr_pipe66_bF_buf3), .B(_2487__bF_buf2), .C(micro_hash_ucr_pipe67), .Y(_4089_) );
OAI21X1 OAI21X1_1300 ( .A(_4201__bF_buf2), .B(_591__bF_buf2), .C(_4199__bF_buf4), .Y(_4090_) );
AOI21X1 AOI21X1_720 ( .A(_4089_), .B(_4088_), .C(_4090_), .Y(_4091_) );
OAI21X1 OAI21X1_1301 ( .A(_4199__bF_buf5), .B(micro_hash_ucr_b_5_bF_buf1_), .C(_344_), .Y(_4092_) );
OAI21X1 OAI21X1_1302 ( .A(_4091_), .B(_4092_), .C(_3992_), .Y(_127__5_) );
NAND2X1 NAND2X1_595 ( .A(micro_hash_ucr_pipe62_bF_buf2), .B(micro_hash_ucr_b_6_bF_buf3_), .Y(_4093_) );
NAND2X1 NAND2X1_596 ( .A(micro_hash_ucr_pipe61_bF_buf3), .B(_845__bF_buf3), .Y(_4094_) );
NAND2X1 NAND2X1_597 ( .A(micro_hash_ucr_pipe60_bF_buf3), .B(micro_hash_ucr_b_6_bF_buf2_), .Y(_4095_) );
NAND2X1 NAND2X1_598 ( .A(micro_hash_ucr_pipe59), .B(_845__bF_buf3), .Y(_4096_) );
NAND2X1 NAND2X1_599 ( .A(micro_hash_ucr_pipe58_bF_buf3), .B(micro_hash_ucr_b_6_bF_buf1_), .Y(_4097_) );
NAND2X1 NAND2X1_600 ( .A(micro_hash_ucr_pipe57_bF_buf2), .B(_845__bF_buf2), .Y(_4098_) );
NAND2X1 NAND2X1_601 ( .A(micro_hash_ucr_pipe56_bF_buf0), .B(micro_hash_ucr_b_6_bF_buf0_), .Y(_4099_) );
NAND2X1 NAND2X1_602 ( .A(micro_hash_ucr_pipe55), .B(_845__bF_buf2), .Y(_4100_) );
NAND2X1 NAND2X1_603 ( .A(micro_hash_ucr_pipe51), .B(micro_hash_ucr_c_2_bF_buf3_), .Y(_4101_) );
NAND2X1 NAND2X1_604 ( .A(micro_hash_ucr_pipe46_bF_buf3), .B(micro_hash_ucr_b_6_bF_buf3_), .Y(_4102_) );
NAND2X1 NAND2X1_605 ( .A(micro_hash_ucr_pipe45), .B(_845__bF_buf1), .Y(_4103_) );
NAND2X1 NAND2X1_606 ( .A(micro_hash_ucr_pipe44_bF_buf3), .B(micro_hash_ucr_b_6_bF_buf2_), .Y(_4104_) );
NAND2X1 NAND2X1_607 ( .A(micro_hash_ucr_pipe43), .B(_845__bF_buf1), .Y(_4105_) );
NAND2X1 NAND2X1_608 ( .A(micro_hash_ucr_pipe42_bF_buf3), .B(micro_hash_ucr_b_6_bF_buf1_), .Y(_4106_) );
NAND2X1 NAND2X1_609 ( .A(micro_hash_ucr_pipe41_bF_buf2), .B(_845__bF_buf1), .Y(_4107_) );
NAND2X1 NAND2X1_610 ( .A(micro_hash_ucr_pipe36_bF_buf2), .B(_399__bF_buf0), .Y(_4108_) );
NAND2X1 NAND2X1_611 ( .A(micro_hash_ucr_pipe35), .B(micro_hash_ucr_c_2_bF_buf2_), .Y(_4109_) );
NAND2X1 NAND2X1_612 ( .A(micro_hash_ucr_pipe34_bF_buf3), .B(_399__bF_buf1), .Y(_4110_) );
NAND2X1 NAND2X1_613 ( .A(micro_hash_ucr_pipe33_bF_buf1), .B(micro_hash_ucr_c_2_bF_buf1_), .Y(_4111_) );
NAND2X1 NAND2X1_614 ( .A(micro_hash_ucr_pipe32_bF_buf4), .B(_399__bF_buf1), .Y(_4112_) );
NAND2X1 NAND2X1_615 ( .A(micro_hash_ucr_pipe31_bF_buf0), .B(micro_hash_ucr_c_2_bF_buf0_), .Y(_4113_) );
NAND2X1 NAND2X1_616 ( .A(micro_hash_ucr_pipe30_bF_buf2), .B(_399__bF_buf1), .Y(_4114_) );
NAND2X1 NAND2X1_617 ( .A(micro_hash_ucr_pipe29), .B(micro_hash_ucr_c_2_bF_buf3_), .Y(_4115_) );
NAND2X1 NAND2X1_618 ( .A(micro_hash_ucr_pipe28_bF_buf1), .B(_399__bF_buf1), .Y(_4116_) );
NAND2X1 NAND2X1_619 ( .A(micro_hash_ucr_pipe27_bF_buf2), .B(micro_hash_ucr_c_2_bF_buf2_), .Y(_4117_) );
NAND2X1 NAND2X1_620 ( .A(micro_hash_ucr_pipe20_bF_buf3), .B(_399__bF_buf2), .Y(_4118_) );
NAND2X1 NAND2X1_621 ( .A(micro_hash_ucr_pipe19), .B(micro_hash_ucr_c_2_bF_buf1_), .Y(_4119_) );
NOR2X1 NOR2X1_738 ( .A(_399__bF_buf2), .B(_624__bF_buf3), .Y(_4120_) );
NAND2X1 NAND2X1_622 ( .A(micro_hash_ucr_pipe17), .B(micro_hash_ucr_c_2_bF_buf0_), .Y(_4121_) );
OAI21X1 OAI21X1_1303 ( .A(_4240_), .B(_845__bF_buf0), .C(_4239__bF_buf0), .Y(_4122_) );
OAI21X1 OAI21X1_1304 ( .A(_4257_), .B(micro_hash_ucr_pipe12_bF_buf1), .C(_399__bF_buf3), .Y(_4123_) );
NOR2X1 NOR2X1_739 ( .A(H_14_), .B(_4266_), .Y(_4124_) );
AOI22X1 AOI22X1_35 ( .A(_4253_), .B(_4124_), .C(_4007_), .D(_845__bF_buf0), .Y(_4125_) );
OAI21X1 OAI21X1_1305 ( .A(_4125_), .B(_4006_), .C(_4123_), .Y(_4126_) );
NOR2X1 NOR2X1_740 ( .A(micro_hash_ucr_pipe13), .B(_399__bF_buf3), .Y(_4127_) );
AOI22X1 AOI22X1_36 ( .A(micro_hash_ucr_pipe12_bF_buf1), .B(_4127_), .C(_4278_), .D(micro_hash_ucr_c_2_bF_buf3_), .Y(_4128_) );
AND2X2 AND2X2_267 ( .A(_4126_), .B(_4128_), .Y(_4129_) );
OAI21X1 OAI21X1_1306 ( .A(_4241__bF_buf0), .B(micro_hash_ucr_b_6_bF_buf0_), .C(_4240_), .Y(_4130_) );
AOI21X1 AOI21X1_721 ( .A(_4241__bF_buf0), .B(_4129_), .C(_4130_), .Y(_4131_) );
AOI21X1 AOI21X1_722 ( .A(micro_hash_ucr_pipe16), .B(_399__bF_buf3), .C(micro_hash_ucr_pipe17), .Y(_4132_) );
OAI21X1 OAI21X1_1307 ( .A(_4131_), .B(_4122_), .C(_4132_), .Y(_4133_) );
AOI21X1 AOI21X1_723 ( .A(_4121_), .B(_4133_), .C(micro_hash_ucr_pipe18_bF_buf0), .Y(_4134_) );
OAI21X1 OAI21X1_1308 ( .A(_4134_), .B(_4120_), .C(_2816_), .Y(_4135_) );
NAND3X1 NAND3X1_234 ( .A(_4237__bF_buf3), .B(_4119_), .C(_4135_), .Y(_4136_) );
NAND3X1 NAND3X1_235 ( .A(_4236__bF_buf0), .B(_4118_), .C(_4136_), .Y(_4137_) );
AOI21X1 AOI21X1_724 ( .A(micro_hash_ucr_pipe21), .B(micro_hash_ucr_c_2_bF_buf2_), .C(micro_hash_ucr_pipe22_bF_buf3), .Y(_4138_) );
OAI21X1 OAI21X1_1309 ( .A(_4262__bF_buf2), .B(micro_hash_ucr_b_6_bF_buf3_), .C(_4234__bF_buf3), .Y(_4139_) );
AOI21X1 AOI21X1_725 ( .A(_4138_), .B(_4137_), .C(_4139_), .Y(_4140_) );
OAI21X1 OAI21X1_1310 ( .A(_4234__bF_buf2), .B(_845__bF_buf0), .C(_4233__bF_buf3), .Y(_4141_) );
OAI22X1 OAI22X1_54 ( .A(micro_hash_ucr_b_6_bF_buf2_), .B(_4233__bF_buf3), .C(_4140_), .D(_4141_), .Y(_4142_) );
OAI21X1 OAI21X1_1311 ( .A(_389__bF_buf3), .B(micro_hash_ucr_c_2_bF_buf1_), .C(_4230__bF_buf1), .Y(_4143_) );
AOI21X1 AOI21X1_726 ( .A(_389__bF_buf1), .B(_4142_), .C(_4143_), .Y(_4144_) );
NOR2X1 NOR2X1_741 ( .A(_399__bF_buf2), .B(_4230__bF_buf1), .Y(_4145_) );
OAI21X1 OAI21X1_1312 ( .A(_4144_), .B(_4145_), .C(_4229_), .Y(_4146_) );
NAND3X1 NAND3X1_236 ( .A(_220__bF_buf2), .B(_4117_), .C(_4146_), .Y(_4147_) );
NAND3X1 NAND3X1_237 ( .A(_219_), .B(_4116_), .C(_4147_), .Y(_4148_) );
NAND3X1 NAND3X1_238 ( .A(_4228__bF_buf3), .B(_4115_), .C(_4148_), .Y(_4149_) );
NAND3X1 NAND3X1_239 ( .A(_317__bF_buf0), .B(_4114_), .C(_4149_), .Y(_4150_) );
NAND3X1 NAND3X1_240 ( .A(_4226__bF_buf2), .B(_4113_), .C(_4150_), .Y(_4151_) );
NAND3X1 NAND3X1_241 ( .A(_318_), .B(_4112_), .C(_4151_), .Y(_4152_) );
NAND3X1 NAND3X1_242 ( .A(_4225__bF_buf1), .B(_4111_), .C(_4152_), .Y(_4153_) );
NAND3X1 NAND3X1_243 ( .A(_230__bF_buf1), .B(_4110_), .C(_4153_), .Y(_4154_) );
NAND3X1 NAND3X1_244 ( .A(_4224__bF_buf0), .B(_4109_), .C(_4154_), .Y(_4155_) );
NAND3X1 NAND3X1_245 ( .A(_2815_), .B(_4108_), .C(_4155_), .Y(_4156_) );
AOI21X1 AOI21X1_727 ( .A(micro_hash_ucr_pipe37_bF_buf1), .B(micro_hash_ucr_c_2_bF_buf0_), .C(micro_hash_ucr_pipe38_bF_buf2), .Y(_4157_) );
OAI21X1 OAI21X1_1313 ( .A(_701__bF_buf1), .B(micro_hash_ucr_b_6_bF_buf1_), .C(_2813__bF_buf2), .Y(_4158_) );
AOI21X1 AOI21X1_728 ( .A(_4157_), .B(_4156_), .C(_4158_), .Y(_4159_) );
OAI21X1 OAI21X1_1314 ( .A(_2813__bF_buf3), .B(_845__bF_buf1), .C(_296__bF_buf0), .Y(_4160_) );
OAI22X1 OAI22X1_55 ( .A(_296__bF_buf0), .B(micro_hash_ucr_b_6_bF_buf0_), .C(_4159_), .D(_4160_), .Y(_4161_) );
NAND2X1 NAND2X1_623 ( .A(_2814_), .B(_4161_), .Y(_4162_) );
NAND3X1 NAND3X1_246 ( .A(_4220__bF_buf1), .B(_4107_), .C(_4162_), .Y(_4163_) );
NAND3X1 NAND3X1_247 ( .A(_242__bF_buf3), .B(_4106_), .C(_4163_), .Y(_4164_) );
NAND3X1 NAND3X1_248 ( .A(_4219__bF_buf4), .B(_4105_), .C(_4164_), .Y(_4165_) );
NAND3X1 NAND3X1_249 ( .A(_336_), .B(_4104_), .C(_4165_), .Y(_4166_) );
NAND3X1 NAND3X1_250 ( .A(_4218__bF_buf0), .B(_4103_), .C(_4166_), .Y(_4167_) );
AOI21X1 AOI21X1_729 ( .A(_4102_), .B(_4167_), .C(micro_hash_ucr_pipe47), .Y(_4168_) );
OAI21X1 OAI21X1_1315 ( .A(_249__bF_buf1), .B(_845__bF_buf2), .C(_4217__bF_buf0), .Y(_4169_) );
AOI21X1 AOI21X1_730 ( .A(micro_hash_ucr_pipe48_bF_buf3), .B(_399__bF_buf0), .C(micro_hash_ucr_pipe49_bF_buf0), .Y(_4170_) );
OAI21X1 OAI21X1_1316 ( .A(_4168_), .B(_4169_), .C(_4170_), .Y(_4171_) );
AOI21X1 AOI21X1_731 ( .A(micro_hash_ucr_pipe49_bF_buf0), .B(micro_hash_ucr_c_2_bF_buf3_), .C(micro_hash_ucr_pipe50_bF_buf1), .Y(_4172_) );
NAND2X1 NAND2X1_624 ( .A(_4172_), .B(_4171_), .Y(_4173_) );
NAND2X1 NAND2X1_625 ( .A(micro_hash_ucr_pipe50_bF_buf3), .B(_399__bF_buf0), .Y(_4174_) );
NAND3X1 NAND3X1_251 ( .A(_255__bF_buf2), .B(_4174_), .C(_4173_), .Y(_4175_) );
AOI21X1 AOI21X1_732 ( .A(_4101_), .B(_4175_), .C(micro_hash_ucr_pipe52_bF_buf0), .Y(_4176_) );
OAI21X1 OAI21X1_1317 ( .A(_4214__bF_buf2), .B(_399__bF_buf0), .C(_2812_), .Y(_4177_) );
AOI21X1 AOI21X1_733 ( .A(micro_hash_ucr_pipe53_bF_buf0), .B(_845__bF_buf2), .C(micro_hash_ucr_pipe54_bF_buf4), .Y(_4178_) );
OAI21X1 OAI21X1_1318 ( .A(_4176_), .B(_4177_), .C(_4178_), .Y(_4179_) );
NAND2X1 NAND2X1_626 ( .A(micro_hash_ucr_pipe54_bF_buf4), .B(micro_hash_ucr_b_6_bF_buf3_), .Y(_4180_) );
NAND3X1 NAND3X1_252 ( .A(_2811__bF_buf0), .B(_4180_), .C(_4179_), .Y(_4181_) );
NAND3X1 NAND3X1_253 ( .A(_832__bF_buf2), .B(_4100_), .C(_4181_), .Y(_4182_) );
NAND3X1 NAND3X1_254 ( .A(_4212_), .B(_4099_), .C(_4182_), .Y(_4183_) );
NAND3X1 NAND3X1_255 ( .A(_4211__bF_buf0), .B(_4098_), .C(_4183_), .Y(_4184_) );
NAND3X1 NAND3X1_256 ( .A(_269_), .B(_4097_), .C(_4184_), .Y(_4185_) );
NAND3X1 NAND3X1_257 ( .A(_4210__bF_buf3), .B(_4096_), .C(_4185_), .Y(_4186_) );
NAND3X1 NAND3X1_258 ( .A(_4208_), .B(_4095_), .C(_4186_), .Y(_4187_) );
NAND3X1 NAND3X1_259 ( .A(_4207__bF_buf2), .B(_4094_), .C(_4187_), .Y(_4188_) );
AOI21X1 AOI21X1_734 ( .A(_4093_), .B(_4188_), .C(micro_hash_ucr_pipe63_bF_buf2), .Y(_4189_) );
OAI21X1 OAI21X1_1319 ( .A(_4204_), .B(_845__bF_buf3), .C(_278__bF_buf0), .Y(_4190_) );
AOI21X1 AOI21X1_735 ( .A(micro_hash_ucr_pipe64_bF_buf1), .B(_399__bF_buf3), .C(micro_hash_ucr_pipe65_bF_buf4), .Y(_4191_) );
OAI21X1 OAI21X1_1320 ( .A(_4189_), .B(_4190_), .C(_4191_), .Y(_4192_) );
AOI21X1 AOI21X1_736 ( .A(micro_hash_ucr_pipe65_bF_buf4), .B(micro_hash_ucr_c_2_bF_buf2_), .C(micro_hash_ucr_pipe66_bF_buf0), .Y(_4193_) );
NOR2X1 NOR2X1_742 ( .A(micro_hash_ucr_b_6_bF_buf2_), .B(_1078__bF_buf1), .Y(_4194_) );
AOI21X1 AOI21X1_737 ( .A(_4193_), .B(_4192_), .C(_4194_), .Y(_4195_) );
OAI21X1 OAI21X1_1321 ( .A(_4201__bF_buf1), .B(_845__bF_buf3), .C(_4199__bF_buf0), .Y(_4196_) );
AOI21X1 AOI21X1_738 ( .A(_4201__bF_buf1), .B(_4195_), .C(_4196_), .Y(_4197_) );
OAI21X1 OAI21X1_1322 ( .A(_4199__bF_buf0), .B(micro_hash_ucr_b_6_bF_buf1_), .C(_344_), .Y(_4198_) );
OAI22X1 OAI22X1_56 ( .A(_845__bF_buf3), .B(_2181_), .C(_4197_), .D(_4198_), .Y(_127__6_) );
DFFPOSX1 DFFPOSX1_388 ( .CLK(clk_bF_buf75), .D(_129__0_), .Q(H_0_) );
DFFPOSX1 DFFPOSX1_389 ( .CLK(clk_bF_buf75), .D(_129__1_), .Q(H_1_) );
DFFPOSX1 DFFPOSX1_390 ( .CLK(clk_bF_buf24), .D(_129__2_), .Q(H_2_) );
DFFPOSX1 DFFPOSX1_391 ( .CLK(clk_bF_buf24), .D(_129__3_), .Q(H_3_) );
DFFPOSX1 DFFPOSX1_392 ( .CLK(clk_bF_buf24), .D(_129__4_), .Q(H_4_) );
DFFPOSX1 DFFPOSX1_393 ( .CLK(clk_bF_buf24), .D(_129__5_), .Q(H_5_) );
DFFPOSX1 DFFPOSX1_394 ( .CLK(clk_bF_buf18), .D(_129__6_), .Q(H_6_) );
DFFPOSX1 DFFPOSX1_395 ( .CLK(clk_bF_buf18), .D(_129__7_), .Q(H_7_) );
DFFPOSX1 DFFPOSX1_396 ( .CLK(clk_bF_buf24), .D(_129__8_), .Q(H_8_) );
DFFPOSX1 DFFPOSX1_397 ( .CLK(clk_bF_buf24), .D(_129__9_), .Q(H_9_) );
DFFPOSX1 DFFPOSX1_398 ( .CLK(clk_bF_buf24), .D(_129__10_), .Q(H_10_) );
DFFPOSX1 DFFPOSX1_399 ( .CLK(clk_bF_buf18), .D(_129__11_), .Q(H_11_) );
DFFPOSX1 DFFPOSX1_400 ( .CLK(clk_bF_buf18), .D(_129__12_), .Q(H_12_) );
DFFPOSX1 DFFPOSX1_401 ( .CLK(clk_bF_buf18), .D(_129__13_), .Q(H_13_) );
DFFPOSX1 DFFPOSX1_402 ( .CLK(clk_bF_buf18), .D(_129__14_), .Q(H_14_) );
DFFPOSX1 DFFPOSX1_403 ( .CLK(clk_bF_buf14), .D(_129__15_), .Q(H_15_) );
DFFPOSX1 DFFPOSX1_404 ( .CLK(clk_bF_buf24), .D(_129__16_), .Q(H_16_) );
DFFPOSX1 DFFPOSX1_405 ( .CLK(clk_bF_buf14), .D(_129__17_), .Q(H_17_) );
DFFPOSX1 DFFPOSX1_406 ( .CLK(clk_bF_buf14), .D(_129__18_), .Q(H_18_) );
DFFPOSX1 DFFPOSX1_407 ( .CLK(clk_bF_buf14), .D(_129__19_), .Q(H_19_) );
DFFPOSX1 DFFPOSX1_408 ( .CLK(clk_bF_buf51), .D(_129__20_), .Q(H_20_) );
DFFPOSX1 DFFPOSX1_409 ( .CLK(clk_bF_buf51), .D(_129__21_), .Q(H_21_) );
DFFPOSX1 DFFPOSX1_410 ( .CLK(clk_bF_buf51), .D(_129__22_), .Q(H_22_) );
DFFPOSX1 DFFPOSX1_411 ( .CLK(clk_bF_buf51), .D(_129__23_), .Q(H_23_) );
DFFPOSX1 DFFPOSX1_412 ( .CLK(clk_bF_buf14), .D(_203_), .Q(comparador_valid_hash) );
DFFPOSX1 DFFPOSX1_413 ( .CLK(clk_bF_buf5), .D(_128__0_), .Q(micro_hash_ucr_c_0_) );
DFFPOSX1 DFFPOSX1_414 ( .CLK(clk_bF_buf5), .D(_128__1_), .Q(micro_hash_ucr_c_1_) );
DFFPOSX1 DFFPOSX1_415 ( .CLK(clk_bF_buf31), .D(_128__2_), .Q(micro_hash_ucr_c_2_) );
DFFPOSX1 DFFPOSX1_416 ( .CLK(clk_bF_buf21), .D(_128__3_), .Q(micro_hash_ucr_c_3_) );
DFFPOSX1 DFFPOSX1_417 ( .CLK(clk_bF_buf48), .D(_128__4_), .Q(micro_hash_ucr_c_4_) );
DFFPOSX1 DFFPOSX1_418 ( .CLK(clk_bF_buf48), .D(_128__5_), .Q(micro_hash_ucr_c_5_) );
DFFPOSX1 DFFPOSX1_419 ( .CLK(clk_bF_buf46), .D(_128__6_), .Q(micro_hash_ucr_c_6_) );
DFFPOSX1 DFFPOSX1_420 ( .CLK(clk_bF_buf80), .D(_128__7_), .Q(micro_hash_ucr_c_7_) );
DFFPOSX1 DFFPOSX1_421 ( .CLK(clk_bF_buf1), .D(_204__0_), .Q(micro_hash_ucr_x_0_) );
DFFPOSX1 DFFPOSX1_422 ( .CLK(clk_bF_buf71), .D(_204__1_), .Q(micro_hash_ucr_x_1_) );
DFFPOSX1 DFFPOSX1_423 ( .CLK(clk_bF_buf1), .D(_204__2_), .Q(micro_hash_ucr_x_2_) );
DFFPOSX1 DFFPOSX1_424 ( .CLK(clk_bF_buf75), .D(_204__3_), .Q(micro_hash_ucr_x_3_) );
DFFPOSX1 DFFPOSX1_425 ( .CLK(clk_bF_buf46), .D(_204__4_), .Q(micro_hash_ucr_x_4_) );
DFFPOSX1 DFFPOSX1_426 ( .CLK(clk_bF_buf48), .D(_204__5_), .Q(micro_hash_ucr_x_5_) );
DFFPOSX1 DFFPOSX1_427 ( .CLK(clk_bF_buf80), .D(_204__6_), .Q(micro_hash_ucr_x_6_) );
DFFPOSX1 DFFPOSX1_428 ( .CLK(clk_bF_buf71), .D(_204__7_), .Q(micro_hash_ucr_x_7_) );
DFFPOSX1 DFFPOSX1_429 ( .CLK(clk_bF_buf21), .D(_130__0_), .Q(micro_hash_ucr_k_0_) );
DFFPOSX1 DFFPOSX1_430 ( .CLK(clk_bF_buf21), .D(_130__1_), .Q(micro_hash_ucr_k_1_) );
DFFPOSX1 DFFPOSX1_431 ( .CLK(clk_bF_buf11), .D(_130__2_), .Q(micro_hash_ucr_k_2_) );
DFFPOSX1 DFFPOSX1_432 ( .CLK(clk_bF_buf48), .D(_130__3_), .Q(micro_hash_ucr_k_3_) );
DFFPOSX1 DFFPOSX1_433 ( .CLK(clk_bF_buf80), .D(_130__4_), .Q(micro_hash_ucr_k_4_) );
DFFPOSX1 DFFPOSX1_434 ( .CLK(clk_bF_buf68), .D(_130__5_), .Q(micro_hash_ucr_k_5_) );
DFFPOSX1 DFFPOSX1_435 ( .CLK(clk_bF_buf46), .D(_130__6_), .Q(micro_hash_ucr_k_6_) );
DFFPOSX1 DFFPOSX1_436 ( .CLK(clk_bF_buf46), .D(_130__7_), .Q(micro_hash_ucr_k_7_) );
DFFPOSX1 DFFPOSX1_437 ( .CLK(clk_bF_buf8), .D(_125__0_), .Q(micro_hash_ucr_Wx_0_) );
DFFPOSX1 DFFPOSX1_438 ( .CLK(clk_bF_buf8), .D(_125__1_), .Q(micro_hash_ucr_Wx_1_) );
DFFPOSX1 DFFPOSX1_439 ( .CLK(clk_bF_buf64), .D(_125__2_), .Q(micro_hash_ucr_Wx_2_) );
DFFPOSX1 DFFPOSX1_440 ( .CLK(clk_bF_buf64), .D(_125__3_), .Q(micro_hash_ucr_Wx_3_) );
DFFPOSX1 DFFPOSX1_441 ( .CLK(clk_bF_buf82), .D(_125__4_), .Q(micro_hash_ucr_Wx_4_) );
DFFPOSX1 DFFPOSX1_442 ( .CLK(clk_bF_buf69), .D(_125__5_), .Q(micro_hash_ucr_Wx_5_) );
DFFPOSX1 DFFPOSX1_443 ( .CLK(clk_bF_buf12), .D(_125__6_), .Q(micro_hash_ucr_Wx_6_) );
DFFPOSX1 DFFPOSX1_444 ( .CLK(clk_bF_buf51), .D(_125__7_), .Q(micro_hash_ucr_Wx_7_) );
DFFPOSX1 DFFPOSX1_445 ( .CLK(clk_bF_buf7), .D(_125__8_), .Q(micro_hash_ucr_Wx_8_) );
DFFPOSX1 DFFPOSX1_446 ( .CLK(clk_bF_buf64), .D(_125__9_), .Q(micro_hash_ucr_Wx_9_) );
DFFPOSX1 DFFPOSX1_447 ( .CLK(clk_bF_buf47), .D(_125__10_), .Q(micro_hash_ucr_Wx_10_) );
DFFPOSX1 DFFPOSX1_448 ( .CLK(clk_bF_buf6), .D(_125__11_), .Q(micro_hash_ucr_Wx_11_) );
DFFPOSX1 DFFPOSX1_449 ( .CLK(clk_bF_buf82), .D(_125__12_), .Q(micro_hash_ucr_Wx_12_) );
DFFPOSX1 DFFPOSX1_450 ( .CLK(clk_bF_buf8), .D(_125__13_), .Q(micro_hash_ucr_Wx_13_) );
DFFPOSX1 DFFPOSX1_451 ( .CLK(clk_bF_buf2), .D(_125__14_), .Q(micro_hash_ucr_Wx_14_) );
DFFPOSX1 DFFPOSX1_452 ( .CLK(clk_bF_buf12), .D(_125__15_), .Q(micro_hash_ucr_Wx_15_) );
DFFPOSX1 DFFPOSX1_453 ( .CLK(clk_bF_buf8), .D(_125__16_), .Q(micro_hash_ucr_Wx_16_) );
DFFPOSX1 DFFPOSX1_454 ( .CLK(clk_bF_buf41), .D(_125__17_), .Q(micro_hash_ucr_Wx_17_) );
DFFPOSX1 DFFPOSX1_455 ( .CLK(clk_bF_buf64), .D(_125__18_), .Q(micro_hash_ucr_Wx_18_) );
DFFPOSX1 DFFPOSX1_456 ( .CLK(clk_bF_buf47), .D(_125__19_), .Q(micro_hash_ucr_Wx_19_) );
DFFPOSX1 DFFPOSX1_457 ( .CLK(clk_bF_buf8), .D(_125__20_), .Q(micro_hash_ucr_Wx_20_) );
DFFPOSX1 DFFPOSX1_458 ( .CLK(clk_bF_buf59), .D(_125__21_), .Q(micro_hash_ucr_Wx_21_) );
DFFPOSX1 DFFPOSX1_459 ( .CLK(clk_bF_buf59), .D(_125__22_), .Q(micro_hash_ucr_Wx_22_) );
DFFPOSX1 DFFPOSX1_460 ( .CLK(clk_bF_buf50), .D(_125__23_), .Q(micro_hash_ucr_Wx_23_) );
DFFPOSX1 DFFPOSX1_461 ( .CLK(clk_bF_buf69), .D(_125__24_), .Q(micro_hash_ucr_Wx_24_) );
DFFPOSX1 DFFPOSX1_462 ( .CLK(clk_bF_buf41), .D(_125__25_), .Q(micro_hash_ucr_Wx_25_) );
DFFPOSX1 DFFPOSX1_463 ( .CLK(clk_bF_buf16), .D(_125__26_), .Q(micro_hash_ucr_Wx_26_) );
DFFPOSX1 DFFPOSX1_464 ( .CLK(clk_bF_buf16), .D(_125__27_), .Q(micro_hash_ucr_Wx_27_) );
DFFPOSX1 DFFPOSX1_465 ( .CLK(clk_bF_buf2), .D(_125__28_), .Q(micro_hash_ucr_Wx_28_) );
DFFPOSX1 DFFPOSX1_466 ( .CLK(clk_bF_buf59), .D(_125__29_), .Q(micro_hash_ucr_Wx_29_) );
DFFPOSX1 DFFPOSX1_467 ( .CLK(clk_bF_buf59), .D(_125__30_), .Q(micro_hash_ucr_Wx_30_) );
DFFPOSX1 DFFPOSX1_468 ( .CLK(clk_bF_buf50), .D(_125__31_), .Q(micro_hash_ucr_Wx_31_) );
DFFPOSX1 DFFPOSX1_469 ( .CLK(clk_bF_buf76), .D(_125__32_), .Q(micro_hash_ucr_Wx_32_) );
DFFPOSX1 DFFPOSX1_470 ( .CLK(clk_bF_buf76), .D(_125__33_), .Q(micro_hash_ucr_Wx_33_) );
DFFPOSX1 DFFPOSX1_471 ( .CLK(clk_bF_buf30), .D(_125__34_), .Q(micro_hash_ucr_Wx_34_) );
DFFPOSX1 DFFPOSX1_472 ( .CLK(clk_bF_buf79), .D(_125__35_), .Q(micro_hash_ucr_Wx_35_) );
DFFPOSX1 DFFPOSX1_473 ( .CLK(clk_bF_buf54), .D(_125__36_), .Q(micro_hash_ucr_Wx_36_) );
DFFPOSX1 DFFPOSX1_474 ( .CLK(clk_bF_buf16), .D(_125__37_), .Q(micro_hash_ucr_Wx_37_) );
DFFPOSX1 DFFPOSX1_475 ( .CLK(clk_bF_buf64), .D(_125__38_), .Q(micro_hash_ucr_Wx_38_) );
DFFPOSX1 DFFPOSX1_476 ( .CLK(clk_bF_buf6), .D(_125__39_), .Q(micro_hash_ucr_Wx_39_) );
DFFPOSX1 DFFPOSX1_477 ( .CLK(clk_bF_buf55), .D(_125__40_), .Q(micro_hash_ucr_Wx_40_) );
DFFPOSX1 DFFPOSX1_478 ( .CLK(clk_bF_buf39), .D(_125__41_), .Q(micro_hash_ucr_Wx_41_) );
DFFPOSX1 DFFPOSX1_479 ( .CLK(clk_bF_buf60), .D(_125__42_), .Q(micro_hash_ucr_Wx_42_) );
DFFPOSX1 DFFPOSX1_480 ( .CLK(clk_bF_buf44), .D(_125__43_), .Q(micro_hash_ucr_Wx_43_) );
DFFPOSX1 DFFPOSX1_481 ( .CLK(clk_bF_buf60), .D(_125__44_), .Q(micro_hash_ucr_Wx_44_) );
DFFPOSX1 DFFPOSX1_482 ( .CLK(clk_bF_buf41), .D(_125__45_), .Q(micro_hash_ucr_Wx_45_) );
DFFPOSX1 DFFPOSX1_483 ( .CLK(clk_bF_buf41), .D(_125__46_), .Q(micro_hash_ucr_Wx_46_) );
DFFPOSX1 DFFPOSX1_484 ( .CLK(clk_bF_buf12), .D(_125__47_), .Q(micro_hash_ucr_Wx_47_) );
DFFPOSX1 DFFPOSX1_485 ( .CLK(clk_bF_buf55), .D(_125__48_), .Q(micro_hash_ucr_Wx_48_) );
DFFPOSX1 DFFPOSX1_486 ( .CLK(clk_bF_buf70), .D(_125__49_), .Q(micro_hash_ucr_Wx_49_) );
DFFPOSX1 DFFPOSX1_487 ( .CLK(clk_bF_buf60), .D(_125__50_), .Q(micro_hash_ucr_Wx_50_) );
DFFPOSX1 DFFPOSX1_488 ( .CLK(clk_bF_buf39), .D(_125__51_), .Q(micro_hash_ucr_Wx_51_) );
DFFPOSX1 DFFPOSX1_489 ( .CLK(clk_bF_buf60), .D(_125__52_), .Q(micro_hash_ucr_Wx_52_) );
DFFPOSX1 DFFPOSX1_490 ( .CLK(clk_bF_buf6), .D(_125__53_), .Q(micro_hash_ucr_Wx_53_) );
DFFPOSX1 DFFPOSX1_491 ( .CLK(clk_bF_buf2), .D(_125__54_), .Q(micro_hash_ucr_Wx_54_) );
DFFPOSX1 DFFPOSX1_492 ( .CLK(clk_bF_buf12), .D(_125__55_), .Q(micro_hash_ucr_Wx_55_) );
DFFPOSX1 DFFPOSX1_493 ( .CLK(clk_bF_buf19), .D(_125__56_), .Q(micro_hash_ucr_Wx_56_) );
DFFPOSX1 DFFPOSX1_494 ( .CLK(clk_bF_buf55), .D(_125__57_), .Q(micro_hash_ucr_Wx_57_) );
DFFPOSX1 DFFPOSX1_495 ( .CLK(clk_bF_buf27), .D(_125__58_), .Q(micro_hash_ucr_Wx_58_) );
DFFPOSX1 DFFPOSX1_496 ( .CLK(clk_bF_buf44), .D(_125__59_), .Q(micro_hash_ucr_Wx_59_) );
DFFPOSX1 DFFPOSX1_497 ( .CLK(clk_bF_buf54), .D(_125__60_), .Q(micro_hash_ucr_Wx_60_) );
DFFPOSX1 DFFPOSX1_498 ( .CLK(clk_bF_buf41), .D(_125__61_), .Q(micro_hash_ucr_Wx_61_) );
DFFPOSX1 DFFPOSX1_499 ( .CLK(clk_bF_buf6), .D(_125__62_), .Q(micro_hash_ucr_Wx_62_) );
DFFPOSX1 DFFPOSX1_500 ( .CLK(clk_bF_buf12), .D(_125__63_), .Q(micro_hash_ucr_Wx_63_) );
DFFPOSX1 DFFPOSX1_501 ( .CLK(clk_bF_buf39), .D(_125__64_), .Q(micro_hash_ucr_Wx_64_) );
DFFPOSX1 DFFPOSX1_502 ( .CLK(clk_bF_buf55), .D(_125__65_), .Q(micro_hash_ucr_Wx_65_) );
DFFPOSX1 DFFPOSX1_503 ( .CLK(clk_bF_buf0), .D(_125__66_), .Q(micro_hash_ucr_Wx_66_) );
DFFPOSX1 DFFPOSX1_504 ( .CLK(clk_bF_buf55), .D(_125__67_), .Q(micro_hash_ucr_Wx_67_) );
DFFPOSX1 DFFPOSX1_505 ( .CLK(clk_bF_buf54), .D(_125__68_), .Q(micro_hash_ucr_Wx_68_) );
DFFPOSX1 DFFPOSX1_506 ( .CLK(clk_bF_buf16), .D(_125__69_), .Q(micro_hash_ucr_Wx_69_) );
DFFPOSX1 DFFPOSX1_507 ( .CLK(clk_bF_buf69), .D(_125__70_), .Q(micro_hash_ucr_Wx_70_) );
DFFPOSX1 DFFPOSX1_508 ( .CLK(clk_bF_buf50), .D(_125__71_), .Q(micro_hash_ucr_Wx_71_) );
DFFPOSX1 DFFPOSX1_509 ( .CLK(clk_bF_buf76), .D(_125__72_), .Q(micro_hash_ucr_Wx_72_) );
DFFPOSX1 DFFPOSX1_510 ( .CLK(clk_bF_buf23), .D(_125__73_), .Q(micro_hash_ucr_Wx_73_) );
DFFPOSX1 DFFPOSX1_511 ( .CLK(clk_bF_buf23), .D(_125__74_), .Q(micro_hash_ucr_Wx_74_) );
DFFPOSX1 DFFPOSX1_512 ( .CLK(clk_bF_buf79), .D(_125__75_), .Q(micro_hash_ucr_Wx_75_) );
DFFPOSX1 DFFPOSX1_513 ( .CLK(clk_bF_buf54), .D(_125__76_), .Q(micro_hash_ucr_Wx_76_) );
DFFPOSX1 DFFPOSX1_514 ( .CLK(clk_bF_buf16), .D(_125__77_), .Q(micro_hash_ucr_Wx_77_) );
DFFPOSX1 DFFPOSX1_515 ( .CLK(clk_bF_buf8), .D(_125__78_), .Q(micro_hash_ucr_Wx_78_) );
DFFPOSX1 DFFPOSX1_516 ( .CLK(clk_bF_buf2), .D(_125__79_), .Q(micro_hash_ucr_Wx_79_) );
DFFPOSX1 DFFPOSX1_517 ( .CLK(clk_bF_buf76), .D(_125__80_), .Q(micro_hash_ucr_Wx_80_) );
DFFPOSX1 DFFPOSX1_518 ( .CLK(clk_bF_buf55), .D(_125__81_), .Q(micro_hash_ucr_Wx_81_) );
DFFPOSX1 DFFPOSX1_519 ( .CLK(clk_bF_buf0), .D(_125__82_), .Q(micro_hash_ucr_Wx_82_) );
DFFPOSX1 DFFPOSX1_520 ( .CLK(clk_bF_buf44), .D(_125__83_), .Q(micro_hash_ucr_Wx_83_) );
DFFPOSX1 DFFPOSX1_521 ( .CLK(clk_bF_buf64), .D(_125__84_), .Q(micro_hash_ucr_Wx_84_) );
DFFPOSX1 DFFPOSX1_522 ( .CLK(clk_bF_buf54), .D(_125__85_), .Q(micro_hash_ucr_Wx_85_) );
DFFPOSX1 DFFPOSX1_523 ( .CLK(clk_bF_buf41), .D(_125__86_), .Q(micro_hash_ucr_Wx_86_) );
DFFPOSX1 DFFPOSX1_524 ( .CLK(clk_bF_buf12), .D(_125__87_), .Q(micro_hash_ucr_Wx_87_) );
DFFPOSX1 DFFPOSX1_525 ( .CLK(clk_bF_buf11), .D(_125__88_), .Q(micro_hash_ucr_Wx_88_) );
DFFPOSX1 DFFPOSX1_526 ( .CLK(clk_bF_buf0), .D(_125__89_), .Q(micro_hash_ucr_Wx_89_) );
DFFPOSX1 DFFPOSX1_527 ( .CLK(clk_bF_buf0), .D(_125__90_), .Q(micro_hash_ucr_Wx_90_) );
DFFPOSX1 DFFPOSX1_528 ( .CLK(clk_bF_buf13), .D(_125__91_), .Q(micro_hash_ucr_Wx_91_) );
DFFPOSX1 DFFPOSX1_529 ( .CLK(clk_bF_buf60), .D(_125__92_), .Q(micro_hash_ucr_Wx_92_) );
DFFPOSX1 DFFPOSX1_530 ( .CLK(clk_bF_buf41), .D(_125__93_), .Q(micro_hash_ucr_Wx_93_) );
DFFPOSX1 DFFPOSX1_531 ( .CLK(clk_bF_buf8), .D(_125__94_), .Q(micro_hash_ucr_Wx_94_) );
DFFPOSX1 DFFPOSX1_532 ( .CLK(clk_bF_buf12), .D(_125__95_), .Q(micro_hash_ucr_Wx_95_) );
DFFPOSX1 DFFPOSX1_533 ( .CLK(clk_bF_buf23), .D(_125__96_), .Q(micro_hash_ucr_Wx_96_) );
DFFPOSX1 DFFPOSX1_534 ( .CLK(clk_bF_buf16), .D(_125__97_), .Q(micro_hash_ucr_Wx_97_) );
DFFPOSX1 DFFPOSX1_535 ( .CLK(clk_bF_buf23), .D(_125__98_), .Q(micro_hash_ucr_Wx_98_) );
DFFPOSX1 DFFPOSX1_536 ( .CLK(clk_bF_buf34), .D(_125__99_), .Q(micro_hash_ucr_Wx_99_) );
DFFPOSX1 DFFPOSX1_537 ( .CLK(clk_bF_buf16), .D(_125__100_), .Q(micro_hash_ucr_Wx_100_) );
DFFPOSX1 DFFPOSX1_538 ( .CLK(clk_bF_buf19), .D(_125__101_), .Q(micro_hash_ucr_Wx_101_) );
DFFPOSX1 DFFPOSX1_539 ( .CLK(clk_bF_buf64), .D(_125__102_), .Q(micro_hash_ucr_Wx_102_) );
DFFPOSX1 DFFPOSX1_540 ( .CLK(clk_bF_buf59), .D(_125__103_), .Q(micro_hash_ucr_Wx_103_) );
DFFPOSX1 DFFPOSX1_541 ( .CLK(clk_bF_buf23), .D(_125__104_), .Q(micro_hash_ucr_Wx_104_) );
DFFPOSX1 DFFPOSX1_542 ( .CLK(clk_bF_buf60), .D(_125__105_), .Q(micro_hash_ucr_Wx_105_) );
DFFPOSX1 DFFPOSX1_543 ( .CLK(clk_bF_buf0), .D(_125__106_), .Q(micro_hash_ucr_Wx_106_) );
DFFPOSX1 DFFPOSX1_544 ( .CLK(clk_bF_buf44), .D(_125__107_), .Q(micro_hash_ucr_Wx_107_) );
DFFPOSX1 DFFPOSX1_545 ( .CLK(clk_bF_buf41), .D(_125__108_), .Q(micro_hash_ucr_Wx_108_) );
DFFPOSX1 DFFPOSX1_546 ( .CLK(clk_bF_buf41), .D(_125__109_), .Q(micro_hash_ucr_Wx_109_) );
DFFPOSX1 DFFPOSX1_547 ( .CLK(clk_bF_buf2), .D(_125__110_), .Q(micro_hash_ucr_Wx_110_) );
DFFPOSX1 DFFPOSX1_548 ( .CLK(clk_bF_buf7), .D(_125__111_), .Q(micro_hash_ucr_Wx_111_) );
DFFPOSX1 DFFPOSX1_549 ( .CLK(clk_bF_buf11), .D(_125__112_), .Q(micro_hash_ucr_Wx_112_) );
DFFPOSX1 DFFPOSX1_550 ( .CLK(clk_bF_buf54), .D(_125__113_), .Q(micro_hash_ucr_Wx_113_) );
DFFPOSX1 DFFPOSX1_551 ( .CLK(clk_bF_buf27), .D(_125__114_), .Q(micro_hash_ucr_Wx_114_) );
DFFPOSX1 DFFPOSX1_552 ( .CLK(clk_bF_buf79), .D(_125__115_), .Q(micro_hash_ucr_Wx_115_) );
DFFPOSX1 DFFPOSX1_553 ( .CLK(clk_bF_buf60), .D(_125__116_), .Q(micro_hash_ucr_Wx_116_) );
DFFPOSX1 DFFPOSX1_554 ( .CLK(clk_bF_buf47), .D(_125__117_), .Q(micro_hash_ucr_Wx_117_) );
DFFPOSX1 DFFPOSX1_555 ( .CLK(clk_bF_buf82), .D(_125__118_), .Q(micro_hash_ucr_Wx_118_) );
DFFPOSX1 DFFPOSX1_556 ( .CLK(clk_bF_buf12), .D(_125__119_), .Q(micro_hash_ucr_Wx_119_) );
DFFPOSX1 DFFPOSX1_557 ( .CLK(clk_bF_buf21), .D(_125__120_), .Q(micro_hash_ucr_Wx_120_) );
DFFPOSX1 DFFPOSX1_558 ( .CLK(clk_bF_buf27), .D(_125__121_), .Q(micro_hash_ucr_Wx_121_) );
DFFPOSX1 DFFPOSX1_559 ( .CLK(clk_bF_buf0), .D(_125__122_), .Q(micro_hash_ucr_Wx_122_) );
DFFPOSX1 DFFPOSX1_560 ( .CLK(clk_bF_buf79), .D(_125__123_), .Q(micro_hash_ucr_Wx_123_) );
DFFPOSX1 DFFPOSX1_561 ( .CLK(clk_bF_buf64), .D(_125__124_), .Q(micro_hash_ucr_Wx_124_) );
DFFPOSX1 DFFPOSX1_562 ( .CLK(clk_bF_buf54), .D(_125__125_), .Q(micro_hash_ucr_Wx_125_) );
DFFPOSX1 DFFPOSX1_563 ( .CLK(clk_bF_buf8), .D(_125__126_), .Q(micro_hash_ucr_Wx_126_) );
DFFPOSX1 DFFPOSX1_564 ( .CLK(clk_bF_buf2), .D(_125__127_), .Q(micro_hash_ucr_Wx_127_) );
DFFPOSX1 DFFPOSX1_565 ( .CLK(clk_bF_buf21), .D(_125__128_), .Q(micro_hash_ucr_Wx_128_) );
DFFPOSX1 DFFPOSX1_566 ( .CLK(clk_bF_buf9), .D(_125__129_), .Q(micro_hash_ucr_Wx_129_) );
DFFPOSX1 DFFPOSX1_567 ( .CLK(clk_bF_buf63), .D(_125__130_), .Q(micro_hash_ucr_Wx_130_) );
DFFPOSX1 DFFPOSX1_568 ( .CLK(clk_bF_buf70), .D(_125__131_), .Q(micro_hash_ucr_Wx_131_) );
DFFPOSX1 DFFPOSX1_569 ( .CLK(clk_bF_buf19), .D(_125__132_), .Q(micro_hash_ucr_Wx_132_) );
DFFPOSX1 DFFPOSX1_570 ( .CLK(clk_bF_buf19), .D(_125__133_), .Q(micro_hash_ucr_Wx_133_) );
DFFPOSX1 DFFPOSX1_571 ( .CLK(clk_bF_buf68), .D(_125__134_), .Q(micro_hash_ucr_Wx_134_) );
DFFPOSX1 DFFPOSX1_572 ( .CLK(clk_bF_buf81), .D(_125__135_), .Q(micro_hash_ucr_Wx_135_) );
DFFPOSX1 DFFPOSX1_573 ( .CLK(clk_bF_buf62), .D(_125__136_), .Q(micro_hash_ucr_Wx_136_) );
DFFPOSX1 DFFPOSX1_574 ( .CLK(clk_bF_buf11), .D(_125__137_), .Q(micro_hash_ucr_Wx_137_) );
DFFPOSX1 DFFPOSX1_575 ( .CLK(clk_bF_buf63), .D(_125__138_), .Q(micro_hash_ucr_Wx_138_) );
DFFPOSX1 DFFPOSX1_576 ( .CLK(clk_bF_buf55), .D(_125__139_), .Q(micro_hash_ucr_Wx_139_) );
DFFPOSX1 DFFPOSX1_577 ( .CLK(clk_bF_buf76), .D(_125__140_), .Q(micro_hash_ucr_Wx_140_) );
DFFPOSX1 DFFPOSX1_578 ( .CLK(clk_bF_buf25), .D(_125__141_), .Q(micro_hash_ucr_Wx_141_) );
DFFPOSX1 DFFPOSX1_579 ( .CLK(clk_bF_buf68), .D(_125__142_), .Q(micro_hash_ucr_Wx_142_) );
DFFPOSX1 DFFPOSX1_580 ( .CLK(clk_bF_buf59), .D(_125__143_), .Q(micro_hash_ucr_Wx_143_) );
DFFPOSX1 DFFPOSX1_581 ( .CLK(clk_bF_buf21), .D(_125__144_), .Q(micro_hash_ucr_Wx_144_) );
DFFPOSX1 DFFPOSX1_582 ( .CLK(clk_bF_buf43), .D(_125__145_), .Q(micro_hash_ucr_Wx_145_) );
DFFPOSX1 DFFPOSX1_583 ( .CLK(clk_bF_buf63), .D(_125__146_), .Q(micro_hash_ucr_Wx_146_) );
DFFPOSX1 DFFPOSX1_584 ( .CLK(clk_bF_buf44), .D(_125__147_), .Q(micro_hash_ucr_Wx_147_) );
DFFPOSX1 DFFPOSX1_585 ( .CLK(clk_bF_buf76), .D(_125__148_), .Q(micro_hash_ucr_Wx_148_) );
DFFPOSX1 DFFPOSX1_586 ( .CLK(clk_bF_buf76), .D(_125__149_), .Q(micro_hash_ucr_Wx_149_) );
DFFPOSX1 DFFPOSX1_587 ( .CLK(clk_bF_buf2), .D(_125__150_), .Q(micro_hash_ucr_Wx_150_) );
DFFPOSX1 DFFPOSX1_588 ( .CLK(clk_bF_buf2), .D(_125__151_), .Q(micro_hash_ucr_Wx_151_) );
DFFPOSX1 DFFPOSX1_589 ( .CLK(clk_bF_buf21), .D(_125__152_), .Q(micro_hash_ucr_Wx_152_) );
DFFPOSX1 DFFPOSX1_590 ( .CLK(clk_bF_buf11), .D(_125__153_), .Q(micro_hash_ucr_Wx_153_) );
DFFPOSX1 DFFPOSX1_591 ( .CLK(clk_bF_buf0), .D(_125__154_), .Q(micro_hash_ucr_Wx_154_) );
DFFPOSX1 DFFPOSX1_592 ( .CLK(clk_bF_buf70), .D(_125__155_), .Q(micro_hash_ucr_Wx_155_) );
DFFPOSX1 DFFPOSX1_593 ( .CLK(clk_bF_buf76), .D(_125__156_), .Q(micro_hash_ucr_Wx_156_) );
DFFPOSX1 DFFPOSX1_594 ( .CLK(clk_bF_buf19), .D(_125__157_), .Q(micro_hash_ucr_Wx_157_) );
DFFPOSX1 DFFPOSX1_595 ( .CLK(clk_bF_buf25), .D(_125__158_), .Q(micro_hash_ucr_Wx_158_) );
DFFPOSX1 DFFPOSX1_596 ( .CLK(clk_bF_buf81), .D(_125__159_), .Q(micro_hash_ucr_Wx_159_) );
DFFPOSX1 DFFPOSX1_597 ( .CLK(clk_bF_buf21), .D(_125__160_), .Q(micro_hash_ucr_Wx_160_) );
DFFPOSX1 DFFPOSX1_598 ( .CLK(clk_bF_buf43), .D(_125__161_), .Q(micro_hash_ucr_Wx_161_) );
DFFPOSX1 DFFPOSX1_599 ( .CLK(clk_bF_buf63), .D(_125__162_), .Q(micro_hash_ucr_Wx_162_) );
DFFPOSX1 DFFPOSX1_600 ( .CLK(clk_bF_buf70), .D(_125__163_), .Q(micro_hash_ucr_Wx_163_) );
DFFPOSX1 DFFPOSX1_601 ( .CLK(clk_bF_buf29), .D(_125__164_), .Q(micro_hash_ucr_Wx_164_) );
DFFPOSX1 DFFPOSX1_602 ( .CLK(clk_bF_buf19), .D(_125__165_), .Q(micro_hash_ucr_Wx_165_) );
DFFPOSX1 DFFPOSX1_603 ( .CLK(clk_bF_buf68), .D(_125__166_), .Q(micro_hash_ucr_Wx_166_) );
DFFPOSX1 DFFPOSX1_604 ( .CLK(clk_bF_buf2), .D(_125__167_), .Q(micro_hash_ucr_Wx_167_) );
DFFPOSX1 DFFPOSX1_605 ( .CLK(clk_bF_buf62), .D(_125__168_), .Q(micro_hash_ucr_Wx_168_) );
DFFPOSX1 DFFPOSX1_606 ( .CLK(clk_bF_buf9), .D(_125__169_), .Q(micro_hash_ucr_Wx_169_) );
DFFPOSX1 DFFPOSX1_607 ( .CLK(clk_bF_buf63), .D(_125__170_), .Q(micro_hash_ucr_Wx_170_) );
DFFPOSX1 DFFPOSX1_608 ( .CLK(clk_bF_buf11), .D(_125__171_), .Q(micro_hash_ucr_Wx_171_) );
DFFPOSX1 DFFPOSX1_609 ( .CLK(clk_bF_buf76), .D(_125__172_), .Q(micro_hash_ucr_Wx_172_) );
DFFPOSX1 DFFPOSX1_610 ( .CLK(clk_bF_buf25), .D(_125__173_), .Q(micro_hash_ucr_Wx_173_) );
DFFPOSX1 DFFPOSX1_611 ( .CLK(clk_bF_buf68), .D(_125__174_), .Q(micro_hash_ucr_Wx_174_) );
DFFPOSX1 DFFPOSX1_612 ( .CLK(clk_bF_buf59), .D(_125__175_), .Q(micro_hash_ucr_Wx_175_) );
DFFPOSX1 DFFPOSX1_613 ( .CLK(clk_bF_buf21), .D(_125__176_), .Q(micro_hash_ucr_Wx_176_) );
DFFPOSX1 DFFPOSX1_614 ( .CLK(clk_bF_buf43), .D(_125__177_), .Q(micro_hash_ucr_Wx_177_) );
DFFPOSX1 DFFPOSX1_615 ( .CLK(clk_bF_buf63), .D(_125__178_), .Q(micro_hash_ucr_Wx_178_) );
DFFPOSX1 DFFPOSX1_616 ( .CLK(clk_bF_buf44), .D(_125__179_), .Q(micro_hash_ucr_Wx_179_) );
DFFPOSX1 DFFPOSX1_617 ( .CLK(clk_bF_buf29), .D(_125__180_), .Q(micro_hash_ucr_Wx_180_) );
DFFPOSX1 DFFPOSX1_618 ( .CLK(clk_bF_buf19), .D(_125__181_), .Q(micro_hash_ucr_Wx_181_) );
DFFPOSX1 DFFPOSX1_619 ( .CLK(clk_bF_buf68), .D(_125__182_), .Q(micro_hash_ucr_Wx_182_) );
DFFPOSX1 DFFPOSX1_620 ( .CLK(clk_bF_buf81), .D(_125__183_), .Q(micro_hash_ucr_Wx_183_) );
DFFPOSX1 DFFPOSX1_621 ( .CLK(clk_bF_buf62), .D(_125__184_), .Q(micro_hash_ucr_Wx_184_) );
DFFPOSX1 DFFPOSX1_622 ( .CLK(clk_bF_buf43), .D(_125__185_), .Q(micro_hash_ucr_Wx_185_) );
DFFPOSX1 DFFPOSX1_623 ( .CLK(clk_bF_buf9), .D(_125__186_), .Q(micro_hash_ucr_Wx_186_) );
DFFPOSX1 DFFPOSX1_624 ( .CLK(clk_bF_buf11), .D(_125__187_), .Q(micro_hash_ucr_Wx_187_) );
DFFPOSX1 DFFPOSX1_625 ( .CLK(clk_bF_buf29), .D(_125__188_), .Q(micro_hash_ucr_Wx_188_) );
DFFPOSX1 DFFPOSX1_626 ( .CLK(clk_bF_buf19), .D(_125__189_), .Q(micro_hash_ucr_Wx_189_) );
DFFPOSX1 DFFPOSX1_627 ( .CLK(clk_bF_buf68), .D(_125__190_), .Q(micro_hash_ucr_Wx_190_) );
DFFPOSX1 DFFPOSX1_628 ( .CLK(clk_bF_buf81), .D(_125__191_), .Q(micro_hash_ucr_Wx_191_) );
DFFPOSX1 DFFPOSX1_629 ( .CLK(clk_bF_buf62), .D(_125__192_), .Q(micro_hash_ucr_Wx_192_) );
DFFPOSX1 DFFPOSX1_630 ( .CLK(clk_bF_buf43), .D(_125__193_), .Q(micro_hash_ucr_Wx_193_) );
DFFPOSX1 DFFPOSX1_631 ( .CLK(clk_bF_buf63), .D(_125__194_), .Q(micro_hash_ucr_Wx_194_) );
DFFPOSX1 DFFPOSX1_632 ( .CLK(clk_bF_buf70), .D(_125__195_), .Q(micro_hash_ucr_Wx_195_) );
DFFPOSX1 DFFPOSX1_633 ( .CLK(clk_bF_buf76), .D(_125__196_), .Q(micro_hash_ucr_Wx_196_) );
DFFPOSX1 DFFPOSX1_634 ( .CLK(clk_bF_buf29), .D(_125__197_), .Q(micro_hash_ucr_Wx_197_) );
DFFPOSX1 DFFPOSX1_635 ( .CLK(clk_bF_buf48), .D(_125__198_), .Q(micro_hash_ucr_Wx_198_) );
DFFPOSX1 DFFPOSX1_636 ( .CLK(clk_bF_buf81), .D(_125__199_), .Q(micro_hash_ucr_Wx_199_) );
DFFPOSX1 DFFPOSX1_637 ( .CLK(clk_bF_buf62), .D(_125__200_), .Q(micro_hash_ucr_Wx_200_) );
DFFPOSX1 DFFPOSX1_638 ( .CLK(clk_bF_buf9), .D(_125__201_), .Q(micro_hash_ucr_Wx_201_) );
DFFPOSX1 DFFPOSX1_639 ( .CLK(clk_bF_buf0), .D(_125__202_), .Q(micro_hash_ucr_Wx_202_) );
DFFPOSX1 DFFPOSX1_640 ( .CLK(clk_bF_buf70), .D(_125__203_), .Q(micro_hash_ucr_Wx_203_) );
DFFPOSX1 DFFPOSX1_641 ( .CLK(clk_bF_buf29), .D(_125__204_), .Q(micro_hash_ucr_Wx_204_) );
DFFPOSX1 DFFPOSX1_642 ( .CLK(clk_bF_buf25), .D(_125__205_), .Q(micro_hash_ucr_Wx_205_) );
DFFPOSX1 DFFPOSX1_643 ( .CLK(clk_bF_buf68), .D(_125__206_), .Q(micro_hash_ucr_Wx_206_) );
DFFPOSX1 DFFPOSX1_644 ( .CLK(clk_bF_buf81), .D(_125__207_), .Q(micro_hash_ucr_Wx_207_) );
DFFPOSX1 DFFPOSX1_645 ( .CLK(clk_bF_buf5), .D(_125__208_), .Q(micro_hash_ucr_Wx_208_) );
DFFPOSX1 DFFPOSX1_646 ( .CLK(clk_bF_buf9), .D(_125__209_), .Q(micro_hash_ucr_Wx_209_) );
DFFPOSX1 DFFPOSX1_647 ( .CLK(clk_bF_buf63), .D(_125__210_), .Q(micro_hash_ucr_Wx_210_) );
DFFPOSX1 DFFPOSX1_648 ( .CLK(clk_bF_buf23), .D(_125__211_), .Q(micro_hash_ucr_Wx_211_) );
DFFPOSX1 DFFPOSX1_649 ( .CLK(clk_bF_buf29), .D(_125__212_), .Q(micro_hash_ucr_Wx_212_) );
DFFPOSX1 DFFPOSX1_650 ( .CLK(clk_bF_buf25), .D(_125__213_), .Q(micro_hash_ucr_Wx_213_) );
DFFPOSX1 DFFPOSX1_651 ( .CLK(clk_bF_buf46), .D(_125__214_), .Q(micro_hash_ucr_Wx_214_) );
DFFPOSX1 DFFPOSX1_652 ( .CLK(clk_bF_buf81), .D(_125__215_), .Q(micro_hash_ucr_Wx_215_) );
DFFPOSX1 DFFPOSX1_653 ( .CLK(clk_bF_buf62), .D(_125__216_), .Q(micro_hash_ucr_Wx_216_) );
DFFPOSX1 DFFPOSX1_654 ( .CLK(clk_bF_buf43), .D(_125__217_), .Q(micro_hash_ucr_Wx_217_) );
DFFPOSX1 DFFPOSX1_655 ( .CLK(clk_bF_buf63), .D(_125__218_), .Q(micro_hash_ucr_Wx_218_) );
DFFPOSX1 DFFPOSX1_656 ( .CLK(clk_bF_buf44), .D(_125__219_), .Q(micro_hash_ucr_Wx_219_) );
DFFPOSX1 DFFPOSX1_657 ( .CLK(clk_bF_buf29), .D(_125__220_), .Q(micro_hash_ucr_Wx_220_) );
DFFPOSX1 DFFPOSX1_658 ( .CLK(clk_bF_buf25), .D(_125__221_), .Q(micro_hash_ucr_Wx_221_) );
DFFPOSX1 DFFPOSX1_659 ( .CLK(clk_bF_buf46), .D(_125__222_), .Q(micro_hash_ucr_Wx_222_) );
DFFPOSX1 DFFPOSX1_660 ( .CLK(clk_bF_buf81), .D(_125__223_), .Q(micro_hash_ucr_Wx_223_) );
DFFPOSX1 DFFPOSX1_661 ( .CLK(clk_bF_buf5), .D(_125__224_), .Q(micro_hash_ucr_Wx_224_) );
DFFPOSX1 DFFPOSX1_662 ( .CLK(clk_bF_buf9), .D(_125__225_), .Q(micro_hash_ucr_Wx_225_) );
DFFPOSX1 DFFPOSX1_663 ( .CLK(clk_bF_buf63), .D(_125__226_), .Q(micro_hash_ucr_Wx_226_) );
DFFPOSX1 DFFPOSX1_664 ( .CLK(clk_bF_buf70), .D(_125__227_), .Q(micro_hash_ucr_Wx_227_) );
DFFPOSX1 DFFPOSX1_665 ( .CLK(clk_bF_buf29), .D(_125__228_), .Q(micro_hash_ucr_Wx_228_) );
DFFPOSX1 DFFPOSX1_666 ( .CLK(clk_bF_buf25), .D(_125__229_), .Q(micro_hash_ucr_Wx_229_) );
DFFPOSX1 DFFPOSX1_667 ( .CLK(clk_bF_buf46), .D(_125__230_), .Q(micro_hash_ucr_Wx_230_) );
DFFPOSX1 DFFPOSX1_668 ( .CLK(clk_bF_buf81), .D(_125__231_), .Q(micro_hash_ucr_Wx_231_) );
DFFPOSX1 DFFPOSX1_669 ( .CLK(clk_bF_buf5), .D(_125__232_), .Q(micro_hash_ucr_Wx_232_) );
DFFPOSX1 DFFPOSX1_670 ( .CLK(clk_bF_buf9), .D(_125__233_), .Q(micro_hash_ucr_Wx_233_) );
DFFPOSX1 DFFPOSX1_671 ( .CLK(clk_bF_buf43), .D(_125__234_), .Q(micro_hash_ucr_Wx_234_) );
DFFPOSX1 DFFPOSX1_672 ( .CLK(clk_bF_buf23), .D(_125__235_), .Q(micro_hash_ucr_Wx_235_) );
DFFPOSX1 DFFPOSX1_673 ( .CLK(clk_bF_buf11), .D(_125__236_), .Q(micro_hash_ucr_Wx_236_) );
DFFPOSX1 DFFPOSX1_674 ( .CLK(clk_bF_buf25), .D(_125__237_), .Q(micro_hash_ucr_Wx_237_) );
DFFPOSX1 DFFPOSX1_675 ( .CLK(clk_bF_buf46), .D(_125__238_), .Q(micro_hash_ucr_Wx_238_) );
DFFPOSX1 DFFPOSX1_676 ( .CLK(clk_bF_buf81), .D(_125__239_), .Q(micro_hash_ucr_Wx_239_) );
DFFPOSX1 DFFPOSX1_677 ( .CLK(clk_bF_buf5), .D(_125__240_), .Q(micro_hash_ucr_Wx_240_) );
DFFPOSX1 DFFPOSX1_678 ( .CLK(clk_bF_buf9), .D(_125__241_), .Q(micro_hash_ucr_Wx_241_) );
DFFPOSX1 DFFPOSX1_679 ( .CLK(clk_bF_buf43), .D(_125__242_), .Q(micro_hash_ucr_Wx_242_) );
DFFPOSX1 DFFPOSX1_680 ( .CLK(clk_bF_buf23), .D(_125__243_), .Q(micro_hash_ucr_Wx_243_) );
DFFPOSX1 DFFPOSX1_681 ( .CLK(clk_bF_buf29), .D(_125__244_), .Q(micro_hash_ucr_Wx_244_) );
DFFPOSX1 DFFPOSX1_682 ( .CLK(clk_bF_buf25), .D(_125__245_), .Q(micro_hash_ucr_Wx_245_) );
DFFPOSX1 DFFPOSX1_683 ( .CLK(clk_bF_buf68), .D(_125__246_), .Q(micro_hash_ucr_Wx_246_) );
DFFPOSX1 DFFPOSX1_684 ( .CLK(clk_bF_buf68), .D(_125__247_), .Q(micro_hash_ucr_Wx_247_) );
DFFPOSX1 DFFPOSX1_685 ( .CLK(clk_bF_buf5), .D(_125__248_), .Q(micro_hash_ucr_Wx_248_) );
DFFPOSX1 DFFPOSX1_686 ( .CLK(clk_bF_buf9), .D(_125__249_), .Q(micro_hash_ucr_Wx_249_) );
DFFPOSX1 DFFPOSX1_687 ( .CLK(clk_bF_buf43), .D(_125__250_), .Q(micro_hash_ucr_Wx_250_) );
DFFPOSX1 DFFPOSX1_688 ( .CLK(clk_bF_buf23), .D(_125__251_), .Q(micro_hash_ucr_Wx_251_) );
DFFPOSX1 DFFPOSX1_689 ( .CLK(clk_bF_buf11), .D(_125__252_), .Q(micro_hash_ucr_Wx_252_) );
DFFPOSX1 DFFPOSX1_690 ( .CLK(clk_bF_buf19), .D(_125__253_), .Q(micro_hash_ucr_Wx_253_) );
DFFPOSX1 DFFPOSX1_691 ( .CLK(clk_bF_buf46), .D(_125__254_), .Q(micro_hash_ucr_Wx_254_) );
DFFPOSX1 DFFPOSX1_692 ( .CLK(clk_bF_buf51), .D(_125__255_), .Q(micro_hash_ucr_Wx_255_) );
DFFPOSX1 DFFPOSX1_693 ( .CLK(clk_bF_buf71), .D(_127__0_), .Q(micro_hash_ucr_b_0_) );
DFFPOSX1 DFFPOSX1_694 ( .CLK(clk_bF_buf71), .D(_127__1_), .Q(micro_hash_ucr_b_1_) );
DFFPOSX1 DFFPOSX1_695 ( .CLK(clk_bF_buf71), .D(_127__2_), .Q(micro_hash_ucr_b_2_) );
DFFPOSX1 DFFPOSX1_696 ( .CLK(clk_bF_buf71), .D(_127__3_), .Q(micro_hash_ucr_b_3_) );
DFFPOSX1 DFFPOSX1_697 ( .CLK(clk_bF_buf83), .D(_127__4_), .Q(micro_hash_ucr_b_4_) );
DFFPOSX1 DFFPOSX1_698 ( .CLK(clk_bF_buf83), .D(_127__5_), .Q(micro_hash_ucr_b_5_) );
DFFPOSX1 DFFPOSX1_699 ( .CLK(clk_bF_buf83), .D(_127__6_), .Q(micro_hash_ucr_b_6_) );
DFFPOSX1 DFFPOSX1_700 ( .CLK(clk_bF_buf71), .D(_127__7_), .Q(micro_hash_ucr_b_7_) );
DFFPOSX1 DFFPOSX1_701 ( .CLK(clk_bF_buf14), .D(_131__bF_buf6), .Q(micro_hash_ucr_pipe0) );
DFFPOSX1 DFFPOSX1_702 ( .CLK(clk_bF_buf83), .D(_126__0_), .Q(micro_hash_ucr_a_0_) );
DFFPOSX1 DFFPOSX1_703 ( .CLK(clk_bF_buf83), .D(_126__1_), .Q(micro_hash_ucr_a_1_) );
DFFPOSX1 DFFPOSX1_704 ( .CLK(clk_bF_buf83), .D(_126__2_), .Q(micro_hash_ucr_a_2_) );
DFFPOSX1 DFFPOSX1_705 ( .CLK(clk_bF_buf75), .D(_126__3_), .Q(micro_hash_ucr_a_3_) );
DFFPOSX1 DFFPOSX1_706 ( .CLK(clk_bF_buf83), .D(_126__4_), .Q(micro_hash_ucr_a_4_) );
DFFPOSX1 DFFPOSX1_707 ( .CLK(clk_bF_buf33), .D(_126__5_), .Q(micro_hash_ucr_a_5_) );
DFFPOSX1 DFFPOSX1_708 ( .CLK(clk_bF_buf71), .D(_126__6_), .Q(micro_hash_ucr_a_6_) );
DFFPOSX1 DFFPOSX1_709 ( .CLK(clk_bF_buf83), .D(_126__7_), .Q(micro_hash_ucr_a_7_) );
DFFPOSX1 DFFPOSX1_710 ( .CLK(clk_bF_buf51), .D(_142_), .Q(micro_hash_ucr_pipe1) );
DFFPOSX1 DFFPOSX1_711 ( .CLK(clk_bF_buf14), .D(_153_), .Q(micro_hash_ucr_pipe2) );
DFFPOSX1 DFFPOSX1_712 ( .CLK(clk_bF_buf15), .D(_164_), .Q(micro_hash_ucr_pipe3) );
DFFPOSX1 DFFPOSX1_713 ( .CLK(clk_bF_buf15), .D(_175_), .Q(micro_hash_ucr_pipe4) );
DFFPOSX1 DFFPOSX1_714 ( .CLK(clk_bF_buf14), .D(_186_), .Q(micro_hash_ucr_pipe5) );
DFFPOSX1 DFFPOSX1_715 ( .CLK(clk_bF_buf18), .D(_197_), .Q(micro_hash_ucr_pipe6) );
DFFPOSX1 DFFPOSX1_716 ( .CLK(clk_bF_buf80), .D(_200_), .Q(micro_hash_ucr_pipe7) );
DFFPOSX1 DFFPOSX1_717 ( .CLK(clk_bF_buf51), .D(_201_), .Q(micro_hash_ucr_pipe8) );
DFFPOSX1 DFFPOSX1_718 ( .CLK(clk_bF_buf80), .D(_202_), .Q(micro_hash_ucr_pipe9) );
DFFPOSX1 DFFPOSX1_719 ( .CLK(clk_bF_buf51), .D(_132_), .Q(micro_hash_ucr_pipe10) );
DFFPOSX1 DFFPOSX1_720 ( .CLK(clk_bF_buf75), .D(_133_), .Q(micro_hash_ucr_pipe11) );
DFFPOSX1 DFFPOSX1_721 ( .CLK(clk_bF_buf24), .D(_134_), .Q(micro_hash_ucr_pipe12) );
DFFPOSX1 DFFPOSX1_722 ( .CLK(clk_bF_buf18), .D(_135_), .Q(micro_hash_ucr_pipe13) );
DFFPOSX1 DFFPOSX1_723 ( .CLK(clk_bF_buf75), .D(_136_), .Q(micro_hash_ucr_pipe14) );
DFFPOSX1 DFFPOSX1_724 ( .CLK(clk_bF_buf75), .D(_137_), .Q(micro_hash_ucr_pipe15) );
DFFPOSX1 DFFPOSX1_725 ( .CLK(clk_bF_buf75), .D(_138_), .Q(micro_hash_ucr_pipe16) );
DFFPOSX1 DFFPOSX1_726 ( .CLK(clk_bF_buf75), .D(_139_), .Q(micro_hash_ucr_pipe17) );
DFFPOSX1 DFFPOSX1_727 ( .CLK(clk_bF_buf80), .D(_140_), .Q(micro_hash_ucr_pipe18) );
DFFPOSX1 DFFPOSX1_728 ( .CLK(clk_bF_buf80), .D(_141_), .Q(micro_hash_ucr_pipe19) );
DFFPOSX1 DFFPOSX1_729 ( .CLK(clk_bF_buf80), .D(_143_), .Q(micro_hash_ucr_pipe20) );
DFFPOSX1 DFFPOSX1_730 ( .CLK(clk_bF_buf75), .D(_144_), .Q(micro_hash_ucr_pipe21) );
DFFPOSX1 DFFPOSX1_731 ( .CLK(clk_bF_buf80), .D(_145_), .Q(micro_hash_ucr_pipe22) );
DFFPOSX1 DFFPOSX1_732 ( .CLK(clk_bF_buf80), .D(_146_), .Q(micro_hash_ucr_pipe23) );
DFFPOSX1 DFFPOSX1_733 ( .CLK(clk_bF_buf48), .D(_147_), .Q(micro_hash_ucr_pipe24) );
DFFPOSX1 DFFPOSX1_734 ( .CLK(clk_bF_buf48), .D(_148_), .Q(micro_hash_ucr_pipe25) );
DFFPOSX1 DFFPOSX1_735 ( .CLK(clk_bF_buf48), .D(_149_), .Q(micro_hash_ucr_pipe26) );
DFFPOSX1 DFFPOSX1_736 ( .CLK(clk_bF_buf48), .D(_150_), .Q(micro_hash_ucr_pipe27) );
DFFPOSX1 DFFPOSX1_737 ( .CLK(clk_bF_buf1), .D(_151_), .Q(micro_hash_ucr_pipe28) );
DFFPOSX1 DFFPOSX1_738 ( .CLK(clk_bF_buf1), .D(_152_), .Q(micro_hash_ucr_pipe29) );
DFFPOSX1 DFFPOSX1_739 ( .CLK(clk_bF_buf1), .D(_154_), .Q(micro_hash_ucr_pipe30) );
DFFPOSX1 DFFPOSX1_740 ( .CLK(clk_bF_buf1), .D(_155_), .Q(micro_hash_ucr_pipe31) );
DFFPOSX1 DFFPOSX1_741 ( .CLK(clk_bF_buf1), .D(_156_), .Q(micro_hash_ucr_pipe32) );
DFFPOSX1 DFFPOSX1_742 ( .CLK(clk_bF_buf1), .D(_157_), .Q(micro_hash_ucr_pipe33) );
DFFPOSX1 DFFPOSX1_743 ( .CLK(clk_bF_buf1), .D(_158_), .Q(micro_hash_ucr_pipe34) );
DFFPOSX1 DFFPOSX1_744 ( .CLK(clk_bF_buf71), .D(_159_), .Q(micro_hash_ucr_pipe35) );
DFFPOSX1 DFFPOSX1_745 ( .CLK(clk_bF_buf62), .D(_160_), .Q(micro_hash_ucr_pipe36) );
DFFPOSX1 DFFPOSX1_746 ( .CLK(clk_bF_buf62), .D(_161_), .Q(micro_hash_ucr_pipe37) );
DFFPOSX1 DFFPOSX1_747 ( .CLK(clk_bF_buf62), .D(_162_), .Q(micro_hash_ucr_pipe38) );
DFFPOSX1 DFFPOSX1_748 ( .CLK(clk_bF_buf62), .D(_163_), .Q(micro_hash_ucr_pipe39) );
DFFPOSX1 DFFPOSX1_749 ( .CLK(clk_bF_buf5), .D(_165_), .Q(micro_hash_ucr_pipe40) );
DFFPOSX1 DFFPOSX1_750 ( .CLK(clk_bF_buf31), .D(_166_), .Q(micro_hash_ucr_pipe41) );
DFFPOSX1 DFFPOSX1_751 ( .CLK(clk_bF_buf31), .D(_167_), .Q(micro_hash_ucr_pipe42) );
DFFPOSX1 DFFPOSX1_752 ( .CLK(clk_bF_buf31), .D(_168_), .Q(micro_hash_ucr_pipe43) );
DFFPOSX1 DFFPOSX1_753 ( .CLK(clk_bF_buf31), .D(_169_), .Q(micro_hash_ucr_pipe44) );
DFFPOSX1 DFFPOSX1_754 ( .CLK(clk_bF_buf3), .D(_170_), .Q(micro_hash_ucr_pipe45) );
DFFPOSX1 DFFPOSX1_755 ( .CLK(clk_bF_buf31), .D(_171_), .Q(micro_hash_ucr_pipe46) );
DFFPOSX1 DFFPOSX1_756 ( .CLK(clk_bF_buf31), .D(_172_), .Q(micro_hash_ucr_pipe47) );
DFFPOSX1 DFFPOSX1_757 ( .CLK(clk_bF_buf31), .D(_173_), .Q(micro_hash_ucr_pipe48) );
DFFPOSX1 DFFPOSX1_758 ( .CLK(clk_bF_buf3), .D(_174_), .Q(micro_hash_ucr_pipe49) );
DFFPOSX1 DFFPOSX1_759 ( .CLK(clk_bF_buf31), .D(_176_), .Q(micro_hash_ucr_pipe50) );
DFFPOSX1 DFFPOSX1_760 ( .CLK(clk_bF_buf3), .D(_177_), .Q(micro_hash_ucr_pipe51) );
DFFPOSX1 DFFPOSX1_761 ( .CLK(clk_bF_buf3), .D(_178_), .Q(micro_hash_ucr_pipe52) );
DFFPOSX1 DFFPOSX1_762 ( .CLK(clk_bF_buf3), .D(_179_), .Q(micro_hash_ucr_pipe53) );
DFFPOSX1 DFFPOSX1_763 ( .CLK(clk_bF_buf3), .D(_180_), .Q(micro_hash_ucr_pipe54) );
DFFPOSX1 DFFPOSX1_764 ( .CLK(clk_bF_buf3), .D(_181_), .Q(micro_hash_ucr_pipe55) );
DFFPOSX1 DFFPOSX1_765 ( .CLK(clk_bF_buf3), .D(_182_), .Q(micro_hash_ucr_pipe56) );
DFFPOSX1 DFFPOSX1_766 ( .CLK(clk_bF_buf33), .D(_183_), .Q(micro_hash_ucr_pipe57) );
DFFPOSX1 DFFPOSX1_767 ( .CLK(clk_bF_buf3), .D(_184_), .Q(micro_hash_ucr_pipe58) );
DFFPOSX1 DFFPOSX1_768 ( .CLK(clk_bF_buf33), .D(_185_), .Q(micro_hash_ucr_pipe59) );
DFFPOSX1 DFFPOSX1_769 ( .CLK(clk_bF_buf33), .D(_187_), .Q(micro_hash_ucr_pipe60) );
DFFPOSX1 DFFPOSX1_770 ( .CLK(clk_bF_buf33), .D(_188_), .Q(micro_hash_ucr_pipe61) );
DFFPOSX1 DFFPOSX1_771 ( .CLK(clk_bF_buf33), .D(_189_), .Q(micro_hash_ucr_pipe62) );
DFFPOSX1 DFFPOSX1_772 ( .CLK(clk_bF_buf33), .D(_190_), .Q(micro_hash_ucr_pipe63) );
DFFPOSX1 DFFPOSX1_773 ( .CLK(clk_bF_buf33), .D(_191_), .Q(micro_hash_ucr_pipe64) );
DFFPOSX1 DFFPOSX1_774 ( .CLK(clk_bF_buf33), .D(_192_), .Q(micro_hash_ucr_pipe65) );
DFFPOSX1 DFFPOSX1_775 ( .CLK(clk_bF_buf83), .D(_193_), .Q(micro_hash_ucr_pipe66) );
DFFPOSX1 DFFPOSX1_776 ( .CLK(clk_bF_buf71), .D(_194_), .Q(micro_hash_ucr_pipe67) );
DFFPOSX1 DFFPOSX1_777 ( .CLK(clk_bF_buf83), .D(_195_), .Q(micro_hash_ucr_pipe68) );
DFFPOSX1 DFFPOSX1_778 ( .CLK(clk_bF_buf5), .D(_196_), .Q(micro_hash_ucr_pipe69) );
DFFPOSX1 DFFPOSX1_779 ( .CLK(clk_bF_buf18), .D(_198_), .Q(micro_hash_ucr_pipe70) );
DFFPOSX1 DFFPOSX1_780 ( .CLK(clk_bF_buf14), .D(_199_), .Q(micro_hash_ucr_pipe71) );
INVX8 INVX8_93 ( .A(reset_bF_buf5), .Y(_4283_) );
NAND2X1 NAND2X1_627 ( .A(next_b_data_in_prev_0_), .B(_4283__bF_buf28), .Y(_4284_) );
MUX2X1 MUX2X1_52 ( .A(data_in[0]), .B(next_b_data_in_prev_0_), .S(_0__bF_buf3), .Y(_4285_) );
OAI21X1 OAI21X1_1323 ( .A(_4285_), .B(_4283__bF_buf28), .C(_4284_), .Y(_4281__0_) );
NAND2X1 NAND2X1_628 ( .A(next_b_data_in_prev_1_), .B(_4283__bF_buf19), .Y(_4286_) );
MUX2X1 MUX2X1_53 ( .A(data_in[1]), .B(next_b_data_in_prev_1_), .S(_0__bF_buf0), .Y(_4287_) );
OAI21X1 OAI21X1_1324 ( .A(_4287_), .B(_4283__bF_buf19), .C(_4286_), .Y(_4281__1_) );
NAND2X1 NAND2X1_629 ( .A(next_b_data_in_prev_2_), .B(_4283__bF_buf6), .Y(_4288_) );
MUX2X1 MUX2X1_54 ( .A(data_in[2]), .B(next_b_data_in_prev_2_), .S(_0__bF_buf3), .Y(_4289_) );
OAI21X1 OAI21X1_1325 ( .A(_4289_), .B(_4283__bF_buf6), .C(_4288_), .Y(_4281__2_) );
NAND2X1 NAND2X1_630 ( .A(next_b_data_in_prev_3_), .B(_4283__bF_buf25), .Y(_4290_) );
MUX2X1 MUX2X1_55 ( .A(data_in[3]), .B(next_b_data_in_prev_3_), .S(_0__bF_buf1), .Y(_4291_) );
OAI21X1 OAI21X1_1326 ( .A(_4291_), .B(_4283__bF_buf25), .C(_4290_), .Y(_4281__3_) );
NAND2X1 NAND2X1_631 ( .A(next_b_data_in_prev_4_), .B(_4283__bF_buf18), .Y(_4292_) );
MUX2X1 MUX2X1_56 ( .A(data_in[4]), .B(next_b_data_in_prev_4_), .S(_0__bF_buf3), .Y(_4293_) );
OAI21X1 OAI21X1_1327 ( .A(_4293_), .B(_4283__bF_buf18), .C(_4292_), .Y(_4281__4_) );
NAND2X1 NAND2X1_632 ( .A(next_b_data_in_prev_5_), .B(_4283__bF_buf33), .Y(_4294_) );
MUX2X1 MUX2X1_57 ( .A(data_in[5]), .B(next_b_data_in_prev_5_), .S(_0__bF_buf4), .Y(_4295_) );
OAI21X1 OAI21X1_1328 ( .A(_4295_), .B(_4283__bF_buf33), .C(_4294_), .Y(_4281__5_) );
NAND2X1 NAND2X1_633 ( .A(next_b_data_in_prev_6_), .B(_4283__bF_buf26), .Y(_4296_) );
MUX2X1 MUX2X1_58 ( .A(data_in[6]), .B(next_b_data_in_prev_6_), .S(_0__bF_buf7), .Y(_4297_) );
OAI21X1 OAI21X1_1329 ( .A(_4297_), .B(_4283__bF_buf26), .C(_4296_), .Y(_4281__6_) );
NAND2X1 NAND2X1_634 ( .A(next_b_data_in_prev_7_), .B(_4283__bF_buf8), .Y(_4298_) );
MUX2X1 MUX2X1_59 ( .A(data_in[7]), .B(next_b_data_in_prev_7_), .S(_0__bF_buf7), .Y(_4299_) );
OAI21X1 OAI21X1_1330 ( .A(_4299_), .B(_4283__bF_buf8), .C(_4298_), .Y(_4281__7_) );
NAND2X1 NAND2X1_635 ( .A(next_b_data_in_prev_8_), .B(_4283__bF_buf21), .Y(_4300_) );
MUX2X1 MUX2X1_60 ( .A(data_in[8]), .B(next_b_data_in_prev_8_), .S(_0__bF_buf0), .Y(_4301_) );
OAI21X1 OAI21X1_1331 ( .A(_4301_), .B(_4283__bF_buf21), .C(_4300_), .Y(_4281__8_) );
NAND2X1 NAND2X1_636 ( .A(next_b_data_in_prev_9_), .B(_4283__bF_buf28), .Y(_4302_) );
MUX2X1 MUX2X1_61 ( .A(data_in[9]), .B(next_b_data_in_prev_9_), .S(_0__bF_buf3), .Y(_4303_) );
OAI21X1 OAI21X1_1332 ( .A(_4303_), .B(_4283__bF_buf28), .C(_4302_), .Y(_4281__9_) );
NAND2X1 NAND2X1_637 ( .A(next_b_data_in_prev_10_), .B(_4283__bF_buf9), .Y(_4304_) );
MUX2X1 MUX2X1_62 ( .A(data_in[10]), .B(next_b_data_in_prev_10_), .S(_0__bF_buf1), .Y(_4305_) );
OAI21X1 OAI21X1_1333 ( .A(_4305_), .B(_4283__bF_buf7), .C(_4304_), .Y(_4281__10_) );
NAND2X1 NAND2X1_638 ( .A(next_b_data_in_prev_11_), .B(_4283__bF_buf34), .Y(_4306_) );
MUX2X1 MUX2X1_63 ( .A(data_in[11]), .B(next_b_data_in_prev_11_), .S(_0__bF_buf3), .Y(_4307_) );
OAI21X1 OAI21X1_1334 ( .A(_4307_), .B(_4283__bF_buf34), .C(_4306_), .Y(_4281__11_) );
NAND2X1 NAND2X1_639 ( .A(next_b_data_in_prev_12_), .B(_4283__bF_buf21), .Y(_4308_) );
MUX2X1 MUX2X1_64 ( .A(data_in[12]), .B(next_b_data_in_prev_12_), .S(_0__bF_buf0), .Y(_4309_) );
OAI21X1 OAI21X1_1335 ( .A(_4309_), .B(_4283__bF_buf21), .C(_4308_), .Y(_4281__12_) );
NAND2X1 NAND2X1_640 ( .A(next_b_data_in_prev_13_), .B(_4283__bF_buf39), .Y(_4310_) );
MUX2X1 MUX2X1_65 ( .A(data_in[13]), .B(next_b_data_in_prev_13_), .S(_0__bF_buf6), .Y(_4311_) );
OAI21X1 OAI21X1_1336 ( .A(_4311_), .B(_4283__bF_buf39), .C(_4310_), .Y(_4281__13_) );
NAND2X1 NAND2X1_641 ( .A(next_b_data_in_prev_14_), .B(_4283__bF_buf39), .Y(_4312_) );
MUX2X1 MUX2X1_66 ( .A(data_in[14]), .B(next_b_data_in_prev_14_), .S(_0__bF_buf6), .Y(_4313_) );
OAI21X1 OAI21X1_1337 ( .A(_4313_), .B(_4283__bF_buf39), .C(_4312_), .Y(_4281__14_) );
NAND2X1 NAND2X1_642 ( .A(next_b_data_in_prev_15_), .B(_4283__bF_buf27), .Y(_4314_) );
MUX2X1 MUX2X1_67 ( .A(data_in[15]), .B(next_b_data_in_prev_15_), .S(_0__bF_buf5), .Y(_4315_) );
OAI21X1 OAI21X1_1338 ( .A(_4315_), .B(_4283__bF_buf27), .C(_4314_), .Y(_4281__15_) );
NAND2X1 NAND2X1_643 ( .A(next_b_data_in_prev_16_), .B(_4283__bF_buf8), .Y(_4316_) );
MUX2X1 MUX2X1_68 ( .A(data_in[16]), .B(next_b_data_in_prev_16_), .S(_0__bF_buf7), .Y(_4317_) );
OAI21X1 OAI21X1_1339 ( .A(_4317_), .B(_4283__bF_buf8), .C(_4316_), .Y(_4281__16_) );
NAND2X1 NAND2X1_644 ( .A(next_b_data_in_prev_17_), .B(_4283__bF_buf42), .Y(_4318_) );
MUX2X1 MUX2X1_69 ( .A(data_in[17]), .B(next_b_data_in_prev_17_), .S(_0__bF_buf8), .Y(_4319_) );
OAI21X1 OAI21X1_1340 ( .A(_4319_), .B(_4283__bF_buf42), .C(_4318_), .Y(_4281__17_) );
NAND2X1 NAND2X1_645 ( .A(next_b_data_in_prev_18_), .B(_4283__bF_buf11), .Y(_4320_) );
MUX2X1 MUX2X1_70 ( .A(data_in[18]), .B(next_b_data_in_prev_18_), .S(_0__bF_buf7), .Y(_4321_) );
OAI21X1 OAI21X1_1341 ( .A(_4321_), .B(_4283__bF_buf30), .C(_4320_), .Y(_4281__18_) );
NAND2X1 NAND2X1_646 ( .A(next_b_data_in_prev_19_), .B(_4283__bF_buf20), .Y(_4322_) );
MUX2X1 MUX2X1_71 ( .A(data_in[19]), .B(next_b_data_in_prev_19_), .S(_0__bF_buf3), .Y(_4323_) );
OAI21X1 OAI21X1_1342 ( .A(_4323_), .B(_4283__bF_buf20), .C(_4322_), .Y(_4281__19_) );
NAND2X1 NAND2X1_647 ( .A(next_b_data_in_prev_20_), .B(_4283__bF_buf8), .Y(_4324_) );
MUX2X1 MUX2X1_72 ( .A(data_in[20]), .B(next_b_data_in_prev_20_), .S(_0__bF_buf7), .Y(_4325_) );
OAI21X1 OAI21X1_1343 ( .A(_4325_), .B(_4283__bF_buf8), .C(_4324_), .Y(_4281__20_) );
NAND2X1 NAND2X1_648 ( .A(next_b_data_in_prev_21_), .B(_4283__bF_buf32), .Y(_4326_) );
MUX2X1 MUX2X1_73 ( .A(data_in[21]), .B(next_b_data_in_prev_21_), .S(_0__bF_buf6), .Y(_4327_) );
OAI21X1 OAI21X1_1344 ( .A(_4327_), .B(_4283__bF_buf32), .C(_4326_), .Y(_4281__21_) );
NAND2X1 NAND2X1_649 ( .A(next_b_data_in_prev_22_), .B(_4283__bF_buf39), .Y(_4328_) );
MUX2X1 MUX2X1_74 ( .A(data_in[22]), .B(next_b_data_in_prev_22_), .S(_0__bF_buf0), .Y(_4329_) );
OAI21X1 OAI21X1_1345 ( .A(_4329_), .B(_4283__bF_buf39), .C(_4328_), .Y(_4281__22_) );
NAND2X1 NAND2X1_650 ( .A(next_b_data_in_prev_23_), .B(_4283__bF_buf29), .Y(_4330_) );
MUX2X1 MUX2X1_75 ( .A(data_in[23]), .B(next_b_data_in_prev_23_), .S(_0__bF_buf6), .Y(_4331_) );
OAI21X1 OAI21X1_1346 ( .A(_4331_), .B(_4283__bF_buf29), .C(_4330_), .Y(_4281__23_) );
NAND2X1 NAND2X1_651 ( .A(next_b_data_in_prev_24_), .B(_4283__bF_buf13), .Y(_4332_) );
MUX2X1 MUX2X1_76 ( .A(data_in[24]), .B(next_b_data_in_prev_24_), .S(_0__bF_buf4), .Y(_4333_) );
OAI21X1 OAI21X1_1347 ( .A(_4333_), .B(_4283__bF_buf33), .C(_4332_), .Y(_4281__24_) );
NAND2X1 NAND2X1_652 ( .A(next_b_data_in_prev_25_), .B(_4283__bF_buf22), .Y(_4334_) );
MUX2X1 MUX2X1_77 ( .A(data_in[25]), .B(next_b_data_in_prev_25_), .S(_0__bF_buf2), .Y(_4335_) );
OAI21X1 OAI21X1_1348 ( .A(_4335_), .B(_4283__bF_buf22), .C(_4334_), .Y(_4281__25_) );
NAND2X1 NAND2X1_653 ( .A(next_b_data_in_prev_26_), .B(_4283__bF_buf12), .Y(_4336_) );
MUX2X1 MUX2X1_78 ( .A(data_in[26]), .B(next_b_data_in_prev_26_), .S(_0__bF_buf8), .Y(_4337_) );
OAI21X1 OAI21X1_1349 ( .A(_4337_), .B(_4283__bF_buf12), .C(_4336_), .Y(_4281__26_) );
NAND2X1 NAND2X1_654 ( .A(next_b_data_in_prev_27_), .B(_4283__bF_buf41), .Y(_4338_) );
MUX2X1 MUX2X1_79 ( .A(data_in[27]), .B(next_b_data_in_prev_27_), .S(_0__bF_buf8), .Y(_4339_) );
OAI21X1 OAI21X1_1350 ( .A(_4339_), .B(_4283__bF_buf41), .C(_4338_), .Y(_4281__27_) );
NAND2X1 NAND2X1_655 ( .A(next_b_data_in_prev_28_), .B(_4283__bF_buf13), .Y(_4340_) );
MUX2X1 MUX2X1_80 ( .A(data_in[28]), .B(next_b_data_in_prev_28_), .S(_0__bF_buf4), .Y(_4341_) );
OAI21X1 OAI21X1_1351 ( .A(_4341_), .B(_4283__bF_buf13), .C(_4340_), .Y(_4281__28_) );
NAND2X1 NAND2X1_656 ( .A(next_b_data_in_prev_29_), .B(_4283__bF_buf1), .Y(_4342_) );
MUX2X1 MUX2X1_81 ( .A(data_in[29]), .B(next_b_data_in_prev_29_), .S(_0__bF_buf5), .Y(_4343_) );
OAI21X1 OAI21X1_1352 ( .A(_4343_), .B(_4283__bF_buf1), .C(_4342_), .Y(_4281__29_) );
NAND2X1 NAND2X1_657 ( .A(next_b_data_in_prev_30_), .B(_4283__bF_buf19), .Y(_4344_) );
MUX2X1 MUX2X1_82 ( .A(data_in[30]), .B(next_b_data_in_prev_30_), .S(_0__bF_buf0), .Y(_4345_) );
OAI21X1 OAI21X1_1353 ( .A(_4345_), .B(_4283__bF_buf19), .C(_4344_), .Y(_4281__30_) );
NAND2X1 NAND2X1_658 ( .A(next_b_data_in_prev_31_), .B(_4283__bF_buf2), .Y(_4346_) );
MUX2X1 MUX2X1_83 ( .A(data_in[31]), .B(next_b_data_in_prev_31_), .S(_0__bF_buf5), .Y(_4347_) );
OAI21X1 OAI21X1_1354 ( .A(_4347_), .B(_4283__bF_buf2), .C(_4346_), .Y(_4281__31_) );
NAND2X1 NAND2X1_659 ( .A(next_b_data_in_prev_32_), .B(_4283__bF_buf36), .Y(_4348_) );
MUX2X1 MUX2X1_84 ( .A(data_in[32]), .B(next_b_data_in_prev_32_), .S(_0__bF_buf4), .Y(_4349_) );
OAI21X1 OAI21X1_1355 ( .A(_4349_), .B(_4283__bF_buf36), .C(_4348_), .Y(_4281__32_) );
NAND2X1 NAND2X1_660 ( .A(next_b_data_in_prev_33_), .B(_4283__bF_buf6), .Y(_4350_) );
MUX2X1 MUX2X1_85 ( .A(data_in[33]), .B(next_b_data_in_prev_33_), .S(_0__bF_buf8), .Y(_4351_) );
OAI21X1 OAI21X1_1356 ( .A(_4351_), .B(_4283__bF_buf6), .C(_4350_), .Y(_4281__33_) );
NAND2X1 NAND2X1_661 ( .A(next_b_data_in_prev_34_), .B(_4283__bF_buf36), .Y(_4352_) );
MUX2X1 MUX2X1_86 ( .A(data_in[34]), .B(next_b_data_in_prev_34_), .S(_0__bF_buf4), .Y(_4353_) );
OAI21X1 OAI21X1_1357 ( .A(_4353_), .B(_4283__bF_buf13), .C(_4352_), .Y(_4281__34_) );
NAND2X1 NAND2X1_662 ( .A(next_b_data_in_prev_35_), .B(_4283__bF_buf5), .Y(_4354_) );
MUX2X1 MUX2X1_87 ( .A(data_in[35]), .B(next_b_data_in_prev_35_), .S(_0__bF_buf2), .Y(_4355_) );
OAI21X1 OAI21X1_1358 ( .A(_4355_), .B(_4283__bF_buf5), .C(_4354_), .Y(_4281__35_) );
NAND2X1 NAND2X1_663 ( .A(next_b_data_in_prev_36_), .B(_4283__bF_buf17), .Y(_4356_) );
MUX2X1 MUX2X1_88 ( .A(data_in[36]), .B(next_b_data_in_prev_36_), .S(_0__bF_buf4), .Y(_4357_) );
OAI21X1 OAI21X1_1359 ( .A(_4357_), .B(_4283__bF_buf17), .C(_4356_), .Y(_4281__36_) );
NAND2X1 NAND2X1_664 ( .A(next_b_data_in_prev_37_), .B(_4283__bF_buf32), .Y(_4358_) );
MUX2X1 MUX2X1_89 ( .A(data_in[37]), .B(next_b_data_in_prev_37_), .S(_0__bF_buf0), .Y(_4359_) );
OAI21X1 OAI21X1_1360 ( .A(_4359_), .B(_4283__bF_buf32), .C(_4358_), .Y(_4281__37_) );
NAND2X1 NAND2X1_665 ( .A(next_b_data_in_prev_38_), .B(_4283__bF_buf2), .Y(_4360_) );
MUX2X1 MUX2X1_90 ( .A(data_in[38]), .B(next_b_data_in_prev_38_), .S(_0__bF_buf5), .Y(_4361_) );
OAI21X1 OAI21X1_1361 ( .A(_4361_), .B(_4283__bF_buf27), .C(_4360_), .Y(_4281__38_) );
NAND2X1 NAND2X1_666 ( .A(next_b_data_in_prev_39_), .B(_4283__bF_buf27), .Y(_4362_) );
MUX2X1 MUX2X1_91 ( .A(data_in[39]), .B(next_b_data_in_prev_39_), .S(_0__bF_buf5), .Y(_4363_) );
OAI21X1 OAI21X1_1362 ( .A(_4363_), .B(_4283__bF_buf27), .C(_4362_), .Y(_4281__39_) );
NAND2X1 NAND2X1_667 ( .A(next_b_data_in_prev_40_), .B(_4283__bF_buf40), .Y(_4364_) );
MUX2X1 MUX2X1_92 ( .A(data_in[40]), .B(next_b_data_in_prev_40_), .S(_0__bF_buf1), .Y(_4365_) );
OAI21X1 OAI21X1_1363 ( .A(_4365_), .B(_4283__bF_buf9), .C(_4364_), .Y(_4281__40_) );
NAND2X1 NAND2X1_668 ( .A(next_b_data_in_prev_41_), .B(_4283__bF_buf23), .Y(_4366_) );
MUX2X1 MUX2X1_93 ( .A(data_in[41]), .B(next_b_data_in_prev_41_), .S(_0__bF_buf4), .Y(_4367_) );
OAI21X1 OAI21X1_1364 ( .A(_4367_), .B(_4283__bF_buf23), .C(_4366_), .Y(_4281__41_) );
NAND2X1 NAND2X1_669 ( .A(next_b_data_in_prev_42_), .B(_4283__bF_buf34), .Y(_4368_) );
MUX2X1 MUX2X1_94 ( .A(data_in[42]), .B(next_b_data_in_prev_42_), .S(_0__bF_buf3), .Y(_4369_) );
OAI21X1 OAI21X1_1365 ( .A(_4369_), .B(_4283__bF_buf34), .C(_4368_), .Y(_4281__42_) );
NAND2X1 NAND2X1_670 ( .A(next_b_data_in_prev_43_), .B(_4283__bF_buf26), .Y(_4370_) );
MUX2X1 MUX2X1_95 ( .A(data_in[43]), .B(next_b_data_in_prev_43_), .S(_0__bF_buf7), .Y(_4371_) );
OAI21X1 OAI21X1_1366 ( .A(_4371_), .B(_4283__bF_buf26), .C(_4370_), .Y(_4281__43_) );
NAND2X1 NAND2X1_671 ( .A(next_b_data_in_prev_44_), .B(_4283__bF_buf9), .Y(_4372_) );
MUX2X1 MUX2X1_96 ( .A(data_in[44]), .B(next_b_data_in_prev_44_), .S(_0__bF_buf2), .Y(_4373_) );
OAI21X1 OAI21X1_1367 ( .A(_4373_), .B(_4283__bF_buf9), .C(_4372_), .Y(_4281__44_) );
NAND2X1 NAND2X1_672 ( .A(next_b_data_in_prev_45_), .B(_4283__bF_buf31), .Y(_4374_) );
MUX2X1 MUX2X1_97 ( .A(data_in[45]), .B(next_b_data_in_prev_45_), .S(_0__bF_buf2), .Y(_4375_) );
OAI21X1 OAI21X1_1368 ( .A(_4375_), .B(_4283__bF_buf31), .C(_4374_), .Y(_4281__45_) );
NAND2X1 NAND2X1_673 ( .A(next_b_data_in_prev_46_), .B(_4283__bF_buf29), .Y(_4376_) );
MUX2X1 MUX2X1_98 ( .A(data_in[46]), .B(next_b_data_in_prev_46_), .S(_0__bF_buf6), .Y(_4377_) );
OAI21X1 OAI21X1_1369 ( .A(_4377_), .B(_4283__bF_buf29), .C(_4376_), .Y(_4281__46_) );
NAND2X1 NAND2X1_674 ( .A(next_b_data_in_prev_47_), .B(_4283__bF_buf29), .Y(_4378_) );
MUX2X1 MUX2X1_99 ( .A(data_in[47]), .B(next_b_data_in_prev_47_), .S(_0__bF_buf6), .Y(_4379_) );
OAI21X1 OAI21X1_1370 ( .A(_4379_), .B(_4283__bF_buf29), .C(_4378_), .Y(_4281__47_) );
NAND2X1 NAND2X1_675 ( .A(next_b_data_in_prev_48_), .B(_4283__bF_buf7), .Y(_4380_) );
MUX2X1 MUX2X1_100 ( .A(data_in[48]), .B(next_b_data_in_prev_48_), .S(_0__bF_buf1), .Y(_4381_) );
OAI21X1 OAI21X1_1371 ( .A(_4381_), .B(_4283__bF_buf0), .C(_4380_), .Y(_4281__48_) );
NAND2X1 NAND2X1_676 ( .A(next_b_data_in_prev_49_), .B(_4283__bF_buf22), .Y(_4382_) );
MUX2X1 MUX2X1_101 ( .A(data_in[49]), .B(next_b_data_in_prev_49_), .S(_0__bF_buf3), .Y(_4383_) );
OAI21X1 OAI21X1_1372 ( .A(_4383_), .B(_4283__bF_buf34), .C(_4382_), .Y(_4281__49_) );
NAND2X1 NAND2X1_677 ( .A(next_b_data_in_prev_50_), .B(_4283__bF_buf42), .Y(_4384_) );
MUX2X1 MUX2X1_102 ( .A(data_in[50]), .B(next_b_data_in_prev_50_), .S(_0__bF_buf8), .Y(_4385_) );
OAI21X1 OAI21X1_1373 ( .A(_4385_), .B(_4283__bF_buf42), .C(_4384_), .Y(_4281__50_) );
NAND2X1 NAND2X1_678 ( .A(next_b_data_in_prev_51_), .B(_4283__bF_buf30), .Y(_4386_) );
MUX2X1 MUX2X1_103 ( .A(data_in[51]), .B(next_b_data_in_prev_51_), .S(_0__bF_buf7), .Y(_4387_) );
OAI21X1 OAI21X1_1374 ( .A(_4387_), .B(_4283__bF_buf30), .C(_4386_), .Y(_4281__51_) );
NAND2X1 NAND2X1_679 ( .A(next_b_data_in_prev_52_), .B(_4283__bF_buf13), .Y(_4388_) );
MUX2X1 MUX2X1_104 ( .A(data_in[52]), .B(next_b_data_in_prev_52_), .S(_0__bF_buf4), .Y(_4389_) );
OAI21X1 OAI21X1_1375 ( .A(_4389_), .B(_4283__bF_buf13), .C(_4388_), .Y(_4281__52_) );
NAND2X1 NAND2X1_680 ( .A(next_b_data_in_prev_53_), .B(_4283__bF_buf15), .Y(_4390_) );
MUX2X1 MUX2X1_105 ( .A(data_in[53]), .B(next_b_data_in_prev_53_), .S(_0__bF_buf8), .Y(_4391_) );
OAI21X1 OAI21X1_1376 ( .A(_4391_), .B(_4283__bF_buf15), .C(_4390_), .Y(_4281__53_) );
NAND2X1 NAND2X1_681 ( .A(next_b_data_in_prev_54_), .B(_4283__bF_buf23), .Y(_4392_) );
MUX2X1 MUX2X1_106 ( .A(data_in[54]), .B(next_b_data_in_prev_54_), .S(_0__bF_buf4), .Y(_4393_) );
OAI21X1 OAI21X1_1377 ( .A(_4393_), .B(_4283__bF_buf23), .C(_4392_), .Y(_4281__54_) );
NAND2X1 NAND2X1_682 ( .A(next_b_data_in_prev_55_), .B(_4283__bF_buf23), .Y(_4394_) );
MUX2X1 MUX2X1_107 ( .A(data_in[55]), .B(next_b_data_in_prev_55_), .S(_0__bF_buf4), .Y(_4395_) );
OAI21X1 OAI21X1_1378 ( .A(_4395_), .B(_4283__bF_buf23), .C(_4394_), .Y(_4281__55_) );
NAND2X1 NAND2X1_683 ( .A(next_b_data_in_prev_56_), .B(_4283__bF_buf24), .Y(_4396_) );
MUX2X1 MUX2X1_108 ( .A(data_in[56]), .B(next_b_data_in_prev_56_), .S(_0__bF_buf6), .Y(_4397_) );
OAI21X1 OAI21X1_1379 ( .A(_4397_), .B(_4283__bF_buf24), .C(_4396_), .Y(_4281__56_) );
NAND2X1 NAND2X1_684 ( .A(next_b_data_in_prev_57_), .B(_4283__bF_buf37), .Y(_4398_) );
MUX2X1 MUX2X1_109 ( .A(data_in[57]), .B(next_b_data_in_prev_57_), .S(_0__bF_buf8), .Y(_4399_) );
OAI21X1 OAI21X1_1380 ( .A(_4399_), .B(_4283__bF_buf37), .C(_4398_), .Y(_4281__57_) );
NAND2X1 NAND2X1_685 ( .A(next_b_data_in_prev_58_), .B(_4283__bF_buf22), .Y(_4400_) );
MUX2X1 MUX2X1_110 ( .A(data_in[58]), .B(next_b_data_in_prev_58_), .S(_0__bF_buf3), .Y(_4401_) );
OAI21X1 OAI21X1_1381 ( .A(_4401_), .B(_4283__bF_buf22), .C(_4400_), .Y(_4281__58_) );
NAND2X1 NAND2X1_686 ( .A(next_b_data_in_prev_59_), .B(_4283__bF_buf22), .Y(_4402_) );
MUX2X1 MUX2X1_111 ( .A(data_in[59]), .B(next_b_data_in_prev_59_), .S(_0__bF_buf2), .Y(_4403_) );
OAI21X1 OAI21X1_1382 ( .A(_4403_), .B(_4283__bF_buf22), .C(_4402_), .Y(_4281__59_) );
NAND2X1 NAND2X1_687 ( .A(next_b_data_in_prev_60_), .B(_4283__bF_buf9), .Y(_4404_) );
MUX2X1 MUX2X1_112 ( .A(data_in[60]), .B(next_b_data_in_prev_60_), .S(_0__bF_buf2), .Y(_4405_) );
OAI21X1 OAI21X1_1383 ( .A(_4405_), .B(_4283__bF_buf9), .C(_4404_), .Y(_4281__60_) );
NAND2X1 NAND2X1_688 ( .A(next_b_data_in_prev_61_), .B(_4283__bF_buf25), .Y(_4406_) );
MUX2X1 MUX2X1_113 ( .A(data_in[61]), .B(next_b_data_in_prev_61_), .S(_0__bF_buf1), .Y(_4407_) );
OAI21X1 OAI21X1_1384 ( .A(_4407_), .B(_4283__bF_buf25), .C(_4406_), .Y(_4281__61_) );
NAND2X1 NAND2X1_689 ( .A(next_b_data_in_prev_62_), .B(_4283__bF_buf32), .Y(_4408_) );
MUX2X1 MUX2X1_114 ( .A(data_in[62]), .B(next_b_data_in_prev_62_), .S(_0__bF_buf6), .Y(_4409_) );
endmodule
