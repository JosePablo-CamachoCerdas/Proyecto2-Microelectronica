module sistemacompletodes ( gnd, vdd, clk, reset, data_in, target, finished, nonce_out);

input gnd, vdd;
input clk;
input reset;
output finished;
input [95:0] data_in;
input [7:0] target;
output [31:0] nonce_out;

BUFX4 BUFX4_1 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf11) );
BUFX4 BUFX4_2 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf10) );
BUFX4 BUFX4_3 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf9) );
BUFX4 BUFX4_4 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf8) );
BUFX4 BUFX4_5 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf7) );
BUFX4 BUFX4_6 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf6) );
BUFX4 BUFX4_7 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf5) );
BUFX4 BUFX4_8 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf4) );
BUFX4 BUFX4_9 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf3) );
BUFX4 BUFX4_10 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf2) );
BUFX4 BUFX4_11 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf1) );
BUFX4 BUFX4_12 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf0) );
BUFX4 BUFX4_13 ( .gnd(gnd), .vdd(vdd), .A(_12916_), .Y(_12916__hier0_bF_buf5) );
BUFX4 BUFX4_14 ( .gnd(gnd), .vdd(vdd), .A(_12916_), .Y(_12916__hier0_bF_buf4) );
BUFX4 BUFX4_15 ( .gnd(gnd), .vdd(vdd), .A(_12916_), .Y(_12916__hier0_bF_buf3) );
BUFX4 BUFX4_16 ( .gnd(gnd), .vdd(vdd), .A(_12916_), .Y(_12916__hier0_bF_buf2) );
BUFX4 BUFX4_17 ( .gnd(gnd), .vdd(vdd), .A(_12916_), .Y(_12916__hier0_bF_buf1) );
BUFX4 BUFX4_18 ( .gnd(gnd), .vdd(vdd), .A(_12916_), .Y(_12916__hier0_bF_buf0) );
BUFX4 BUFX4_19 ( .gnd(gnd), .vdd(vdd), .A(_4608_), .Y(_4608__bF_buf3) );
BUFX4 BUFX4_20 ( .gnd(gnd), .vdd(vdd), .A(_4608_), .Y(_4608__bF_buf2) );
BUFX4 BUFX4_21 ( .gnd(gnd), .vdd(vdd), .A(_4608_), .Y(_4608__bF_buf1) );
BUFX4 BUFX4_22 ( .gnd(gnd), .vdd(vdd), .A(_4608_), .Y(_4608__bF_buf0) );
BUFX4 BUFX4_23 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_6_), .Y(micro_hash_ucr_3_a_6_bF_buf3_) );
BUFX4 BUFX4_24 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_6_), .Y(micro_hash_ucr_3_a_6_bF_buf2_) );
BUFX4 BUFX4_25 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_6_), .Y(micro_hash_ucr_3_a_6_bF_buf1_) );
BUFX4 BUFX4_26 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_6_), .Y(micro_hash_ucr_3_a_6_bF_buf0_) );
BUFX4 BUFX4_27 ( .gnd(gnd), .vdd(vdd), .A(_10387_), .Y(_10387__bF_buf3) );
BUFX4 BUFX4_28 ( .gnd(gnd), .vdd(vdd), .A(_10387_), .Y(_10387__bF_buf2) );
BUFX4 BUFX4_29 ( .gnd(gnd), .vdd(vdd), .A(_10387_), .Y(_10387__bF_buf1) );
BUFX4 BUFX4_30 ( .gnd(gnd), .vdd(vdd), .A(_10387_), .Y(_10387__bF_buf0) );
BUFX4 BUFX4_31 ( .gnd(gnd), .vdd(vdd), .A(_13356_), .Y(_13356__bF_buf4) );
BUFX4 BUFX4_32 ( .gnd(gnd), .vdd(vdd), .A(_13356_), .Y(_13356__bF_buf3) );
BUFX4 BUFX4_33 ( .gnd(gnd), .vdd(vdd), .A(_13356_), .Y(_13356__bF_buf2) );
BUFX4 BUFX4_34 ( .gnd(gnd), .vdd(vdd), .A(_13356_), .Y(_13356__bF_buf1) );
BUFX4 BUFX4_35 ( .gnd(gnd), .vdd(vdd), .A(_13356_), .Y(_13356__bF_buf0) );
BUFX4 BUFX4_36 ( .gnd(gnd), .vdd(vdd), .A(_5087_), .Y(_5087__bF_buf4) );
BUFX4 BUFX4_37 ( .gnd(gnd), .vdd(vdd), .A(_5087_), .Y(_5087__bF_buf3) );
BUFX4 BUFX4_38 ( .gnd(gnd), .vdd(vdd), .A(_5087_), .Y(_5087__bF_buf2) );
BUFX4 BUFX4_39 ( .gnd(gnd), .vdd(vdd), .A(_5087_), .Y(_5087__bF_buf1) );
BUFX4 BUFX4_40 ( .gnd(gnd), .vdd(vdd), .A(_5087_), .Y(_5087__bF_buf0) );
BUFX4 BUFX4_41 ( .gnd(gnd), .vdd(vdd), .A(_9299_), .Y(_9299__bF_buf3) );
BUFX4 BUFX4_42 ( .gnd(gnd), .vdd(vdd), .A(_9299_), .Y(_9299__bF_buf2) );
BUFX4 BUFX4_43 ( .gnd(gnd), .vdd(vdd), .A(_9299_), .Y(_9299__bF_buf1) );
BUFX4 BUFX4_44 ( .gnd(gnd), .vdd(vdd), .A(_9299_), .Y(_9299__bF_buf0) );
BUFX4 BUFX4_45 ( .gnd(gnd), .vdd(vdd), .A(_3094_), .Y(_3094__bF_buf3) );
BUFX4 BUFX4_46 ( .gnd(gnd), .vdd(vdd), .A(_3094_), .Y(_3094__bF_buf2) );
BUFX4 BUFX4_47 ( .gnd(gnd), .vdd(vdd), .A(_3094_), .Y(_3094__bF_buf1) );
BUFX4 BUFX4_48 ( .gnd(gnd), .vdd(vdd), .A(_3094_), .Y(_3094__bF_buf0) );
BUFX4 BUFX4_49 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_0_), .Y(micro_hash_ucr_3_b_0_bF_buf3_) );
BUFX4 BUFX4_50 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_0_), .Y(micro_hash_ucr_3_b_0_bF_buf2_) );
BUFX4 BUFX4_51 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_0_), .Y(micro_hash_ucr_3_b_0_bF_buf1_) );
BUFX4 BUFX4_52 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_0_), .Y(micro_hash_ucr_3_b_0_bF_buf0_) );
BUFX4 BUFX4_53 ( .gnd(gnd), .vdd(vdd), .A(_5105_), .Y(_5105__bF_buf4) );
BUFX4 BUFX4_54 ( .gnd(gnd), .vdd(vdd), .A(_5105_), .Y(_5105__bF_buf3) );
BUFX4 BUFX4_55 ( .gnd(gnd), .vdd(vdd), .A(_5105_), .Y(_5105__bF_buf2) );
BUFX4 BUFX4_56 ( .gnd(gnd), .vdd(vdd), .A(_5105_), .Y(_5105__bF_buf1) );
BUFX4 BUFX4_57 ( .gnd(gnd), .vdd(vdd), .A(_5105_), .Y(_5105__bF_buf0) );
BUFX4 BUFX4_58 ( .gnd(gnd), .vdd(vdd), .A(_9317_), .Y(_9317__bF_buf4) );
BUFX4 BUFX4_59 ( .gnd(gnd), .vdd(vdd), .A(_9317_), .Y(_9317__bF_buf3) );
BUFX4 BUFX4_60 ( .gnd(gnd), .vdd(vdd), .A(_9317_), .Y(_9317__bF_buf2) );
BUFX4 BUFX4_61 ( .gnd(gnd), .vdd(vdd), .A(_9317_), .Y(_9317__bF_buf1) );
BUFX4 BUFX4_62 ( .gnd(gnd), .vdd(vdd), .A(_9317_), .Y(_9317__bF_buf0) );
BUFX4 BUFX4_63 ( .gnd(gnd), .vdd(vdd), .A(_5084_), .Y(_5084__bF_buf3) );
BUFX4 BUFX4_64 ( .gnd(gnd), .vdd(vdd), .A(_5084_), .Y(_5084__bF_buf2) );
BUFX4 BUFX4_65 ( .gnd(gnd), .vdd(vdd), .A(_5084_), .Y(_5084__bF_buf1) );
BUFX4 BUFX4_66 ( .gnd(gnd), .vdd(vdd), .A(_5084_), .Y(_5084__bF_buf0) );
BUFX4 BUFX4_67 ( .gnd(gnd), .vdd(vdd), .A(_5598_), .Y(_5598__bF_buf3) );
BUFX4 BUFX4_68 ( .gnd(gnd), .vdd(vdd), .A(_5598_), .Y(_5598__bF_buf2) );
BUFX4 BUFX4_69 ( .gnd(gnd), .vdd(vdd), .A(_5598_), .Y(_5598__bF_buf1) );
BUFX4 BUFX4_70 ( .gnd(gnd), .vdd(vdd), .A(_5598_), .Y(_5598__bF_buf0) );
BUFX4 BUFX4_71 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe50), .Y(micro_hash_ucr_pipe50_bF_buf3) );
BUFX4 BUFX4_72 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe50), .Y(micro_hash_ucr_pipe50_bF_buf2) );
BUFX4 BUFX4_73 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe50), .Y(micro_hash_ucr_pipe50_bF_buf1) );
BUFX4 BUFX4_74 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe50), .Y(micro_hash_ucr_pipe50_bF_buf0) );
BUFX4 BUFX4_75 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe52), .Y(micro_hash_ucr_pipe52_bF_buf4) );
BUFX4 BUFX4_76 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe52), .Y(micro_hash_ucr_pipe52_bF_buf3) );
BUFX4 BUFX4_77 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe52), .Y(micro_hash_ucr_pipe52_bF_buf2) );
BUFX4 BUFX4_78 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe52), .Y(micro_hash_ucr_pipe52_bF_buf1) );
BUFX4 BUFX4_79 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe52), .Y(micro_hash_ucr_pipe52_bF_buf0) );
BUFX4 BUFX4_80 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe53), .Y(micro_hash_ucr_pipe53_bF_buf3) );
BUFX4 BUFX4_81 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe53), .Y(micro_hash_ucr_pipe53_bF_buf2) );
BUFX4 BUFX4_82 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe53), .Y(micro_hash_ucr_pipe53_bF_buf1) );
BUFX4 BUFX4_83 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe53), .Y(micro_hash_ucr_pipe53_bF_buf0) );
BUFX4 BUFX4_84 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe54), .Y(micro_hash_ucr_pipe54_bF_buf3) );
BUFX4 BUFX4_85 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe54), .Y(micro_hash_ucr_pipe54_bF_buf2) );
BUFX4 BUFX4_86 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe54), .Y(micro_hash_ucr_pipe54_bF_buf1) );
BUFX4 BUFX4_87 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe54), .Y(micro_hash_ucr_pipe54_bF_buf0) );
BUFX4 BUFX4_88 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe56), .Y(micro_hash_ucr_pipe56_bF_buf3) );
BUFX4 BUFX4_89 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe56), .Y(micro_hash_ucr_pipe56_bF_buf2) );
BUFX4 BUFX4_90 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe56), .Y(micro_hash_ucr_pipe56_bF_buf1) );
BUFX4 BUFX4_91 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe56), .Y(micro_hash_ucr_pipe56_bF_buf0) );
BUFX4 BUFX4_92 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe57), .Y(micro_hash_ucr_pipe57_bF_buf3) );
BUFX4 BUFX4_93 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe57), .Y(micro_hash_ucr_pipe57_bF_buf2) );
BUFX4 BUFX4_94 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe57), .Y(micro_hash_ucr_pipe57_bF_buf1) );
BUFX4 BUFX4_95 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe57), .Y(micro_hash_ucr_pipe57_bF_buf0) );
BUFX4 BUFX4_96 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe58), .Y(micro_hash_ucr_pipe58_bF_buf4) );
BUFX4 BUFX4_97 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe58), .Y(micro_hash_ucr_pipe58_bF_buf3) );
BUFX4 BUFX4_98 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe58), .Y(micro_hash_ucr_pipe58_bF_buf2) );
BUFX4 BUFX4_99 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe58), .Y(micro_hash_ucr_pipe58_bF_buf1) );
BUFX4 BUFX4_100 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe58), .Y(micro_hash_ucr_pipe58_bF_buf0) );
BUFX4 BUFX4_101 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_3_), .Y(micro_hash_ucr_c_3_bF_buf4_) );
BUFX4 BUFX4_102 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_3_), .Y(micro_hash_ucr_c_3_bF_buf3_) );
BUFX4 BUFX4_103 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_3_), .Y(micro_hash_ucr_c_3_bF_buf2_) );
BUFX4 BUFX4_104 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_3_), .Y(micro_hash_ucr_c_3_bF_buf1_) );
BUFX4 BUFX4_105 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_3_), .Y(micro_hash_ucr_c_3_bF_buf0_) );
BUFX4 BUFX4_106 ( .gnd(gnd), .vdd(vdd), .A(_926_), .Y(_926__bF_buf4) );
BUFX4 BUFX4_107 ( .gnd(gnd), .vdd(vdd), .A(_926_), .Y(_926__bF_buf3) );
BUFX4 BUFX4_108 ( .gnd(gnd), .vdd(vdd), .A(_926_), .Y(_926__bF_buf2) );
BUFX4 BUFX4_109 ( .gnd(gnd), .vdd(vdd), .A(_926_), .Y(_926__bF_buf1) );
BUFX4 BUFX4_110 ( .gnd(gnd), .vdd(vdd), .A(_926_), .Y(_926__bF_buf0) );
BUFX4 BUFX4_111 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_6_), .Y(micro_hash_ucr_b_6_bF_buf3_) );
BUFX4 BUFX4_112 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_6_), .Y(micro_hash_ucr_b_6_bF_buf2_) );
BUFX4 BUFX4_113 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_6_), .Y(micro_hash_ucr_b_6_bF_buf1_) );
BUFX4 BUFX4_114 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_6_), .Y(micro_hash_ucr_b_6_bF_buf0_) );
BUFX4 BUFX4_115 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_0_), .Y(micro_hash_ucr_3_a_0_bF_buf3_) );
BUFX4 BUFX4_116 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_0_), .Y(micro_hash_ucr_3_a_0_bF_buf2_) );
BUFX4 BUFX4_117 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_0_), .Y(micro_hash_ucr_3_a_0_bF_buf1_) );
BUFX4 BUFX4_118 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_0_), .Y(micro_hash_ucr_3_a_0_bF_buf0_) );
BUFX4 BUFX4_119 ( .gnd(gnd), .vdd(vdd), .A(_1956_), .Y(_1956__bF_buf5) );
BUFX4 BUFX4_120 ( .gnd(gnd), .vdd(vdd), .A(_1956_), .Y(_1956__bF_buf4) );
BUFX4 BUFX4_121 ( .gnd(gnd), .vdd(vdd), .A(_1956_), .Y(_1956__bF_buf3) );
BUFX4 BUFX4_122 ( .gnd(gnd), .vdd(vdd), .A(_1956_), .Y(_1956__bF_buf2) );
BUFX4 BUFX4_123 ( .gnd(gnd), .vdd(vdd), .A(_1956_), .Y(_1956__bF_buf1) );
BUFX4 BUFX4_124 ( .gnd(gnd), .vdd(vdd), .A(_1956_), .Y(_1956__bF_buf0) );
BUFX4 BUFX4_125 ( .gnd(gnd), .vdd(vdd), .A(_6154_), .Y(_6154__bF_buf3) );
BUFX4 BUFX4_126 ( .gnd(gnd), .vdd(vdd), .A(_6154_), .Y(_6154__bF_buf2) );
BUFX4 BUFX4_127 ( .gnd(gnd), .vdd(vdd), .A(_6154_), .Y(_6154__bF_buf1) );
BUFX4 BUFX4_128 ( .gnd(gnd), .vdd(vdd), .A(_6154_), .Y(_6154__bF_buf0) );
BUFX4 BUFX4_129 ( .gnd(gnd), .vdd(vdd), .A(_8814_), .Y(_8814__bF_buf3) );
BUFX4 BUFX4_130 ( .gnd(gnd), .vdd(vdd), .A(_8814_), .Y(_8814__bF_buf2) );
BUFX4 BUFX4_131 ( .gnd(gnd), .vdd(vdd), .A(_8814_), .Y(_8814__bF_buf1) );
BUFX4 BUFX4_132 ( .gnd(gnd), .vdd(vdd), .A(_8814_), .Y(_8814__bF_buf0) );
BUFX4 BUFX4_133 ( .gnd(gnd), .vdd(vdd), .A(_5081_), .Y(_5081__bF_buf3) );
BUFX4 BUFX4_134 ( .gnd(gnd), .vdd(vdd), .A(_5081_), .Y(_5081__bF_buf2) );
BUFX4 BUFX4_135 ( .gnd(gnd), .vdd(vdd), .A(_5081_), .Y(_5081__bF_buf1) );
BUFX4 BUFX4_136 ( .gnd(gnd), .vdd(vdd), .A(_5081_), .Y(_5081__bF_buf0) );
BUFX4 BUFX4_137 ( .gnd(gnd), .vdd(vdd), .A(_10798_), .Y(_10798__bF_buf5) );
BUFX4 BUFX4_138 ( .gnd(gnd), .vdd(vdd), .A(_10798_), .Y(_10798__bF_buf4) );
BUFX4 BUFX4_139 ( .gnd(gnd), .vdd(vdd), .A(_10798_), .Y(_10798__bF_buf3) );
BUFX4 BUFX4_140 ( .gnd(gnd), .vdd(vdd), .A(_10798_), .Y(_10798__bF_buf2) );
BUFX4 BUFX4_141 ( .gnd(gnd), .vdd(vdd), .A(_10798_), .Y(_10798__bF_buf1) );
BUFX4 BUFX4_142 ( .gnd(gnd), .vdd(vdd), .A(_10798_), .Y(_10798__bF_buf0) );
BUFX4 BUFX4_143 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe20), .Y(micro_hash_ucr_pipe20_bF_buf4) );
BUFX4 BUFX4_144 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe20), .Y(micro_hash_ucr_pipe20_bF_buf3) );
BUFX4 BUFX4_145 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe20), .Y(micro_hash_ucr_pipe20_bF_buf2) );
BUFX4 BUFX4_146 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe20), .Y(micro_hash_ucr_pipe20_bF_buf1) );
BUFX4 BUFX4_147 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe20), .Y(micro_hash_ucr_pipe20_bF_buf0) );
BUFX4 BUFX4_148 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe21), .Y(micro_hash_ucr_pipe21_bF_buf3) );
BUFX4 BUFX4_149 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe21), .Y(micro_hash_ucr_pipe21_bF_buf2) );
BUFX4 BUFX4_150 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe21), .Y(micro_hash_ucr_pipe21_bF_buf1) );
BUFX4 BUFX4_151 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe21), .Y(micro_hash_ucr_pipe21_bF_buf0) );
BUFX4 BUFX4_152 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe22), .Y(micro_hash_ucr_pipe22_bF_buf4) );
BUFX4 BUFX4_153 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe22), .Y(micro_hash_ucr_pipe22_bF_buf3) );
BUFX4 BUFX4_154 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe22), .Y(micro_hash_ucr_pipe22_bF_buf2) );
BUFX4 BUFX4_155 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe22), .Y(micro_hash_ucr_pipe22_bF_buf1) );
BUFX4 BUFX4_156 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe22), .Y(micro_hash_ucr_pipe22_bF_buf0) );
BUFX4 BUFX4_157 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe23), .Y(micro_hash_ucr_pipe23_bF_buf3) );
BUFX4 BUFX4_158 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe23), .Y(micro_hash_ucr_pipe23_bF_buf2) );
BUFX4 BUFX4_159 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe23), .Y(micro_hash_ucr_pipe23_bF_buf1) );
BUFX4 BUFX4_160 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe23), .Y(micro_hash_ucr_pipe23_bF_buf0) );
BUFX4 BUFX4_161 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe24), .Y(micro_hash_ucr_pipe24_bF_buf4) );
BUFX4 BUFX4_162 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe24), .Y(micro_hash_ucr_pipe24_bF_buf3) );
BUFX4 BUFX4_163 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe24), .Y(micro_hash_ucr_pipe24_bF_buf2) );
BUFX4 BUFX4_164 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe24), .Y(micro_hash_ucr_pipe24_bF_buf1) );
BUFX4 BUFX4_165 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe24), .Y(micro_hash_ucr_pipe24_bF_buf0) );
BUFX4 BUFX4_166 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe26), .Y(micro_hash_ucr_pipe26_bF_buf3) );
BUFX4 BUFX4_167 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe26), .Y(micro_hash_ucr_pipe26_bF_buf2) );
BUFX4 BUFX4_168 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe26), .Y(micro_hash_ucr_pipe26_bF_buf1) );
BUFX4 BUFX4_169 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe26), .Y(micro_hash_ucr_pipe26_bF_buf0) );
BUFX4 BUFX4_170 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe28), .Y(micro_hash_ucr_pipe28_bF_buf3) );
BUFX4 BUFX4_171 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe28), .Y(micro_hash_ucr_pipe28_bF_buf2) );
BUFX4 BUFX4_172 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe28), .Y(micro_hash_ucr_pipe28_bF_buf1) );
BUFX4 BUFX4_173 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe28), .Y(micro_hash_ucr_pipe28_bF_buf0) );
BUFX4 BUFX4_174 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe29), .Y(micro_hash_ucr_pipe29_bF_buf3) );
BUFX4 BUFX4_175 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe29), .Y(micro_hash_ucr_pipe29_bF_buf2) );
BUFX4 BUFX4_176 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe29), .Y(micro_hash_ucr_pipe29_bF_buf1) );
BUFX4 BUFX4_177 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe29), .Y(micro_hash_ucr_pipe29_bF_buf0) );
BUFX4 BUFX4_178 ( .gnd(gnd), .vdd(vdd), .A(_9293_), .Y(_9293__bF_buf3) );
BUFX4 BUFX4_179 ( .gnd(gnd), .vdd(vdd), .A(_9293_), .Y(_9293__bF_buf2) );
BUFX4 BUFX4_180 ( .gnd(gnd), .vdd(vdd), .A(_9293_), .Y(_9293__bF_buf1) );
BUFX4 BUFX4_181 ( .gnd(gnd), .vdd(vdd), .A(_9293_), .Y(_9293__bF_buf0) );
BUFX4 BUFX4_182 ( .gnd(gnd), .vdd(vdd), .A(_3106_), .Y(_3106__bF_buf5) );
BUFX4 BUFX4_183 ( .gnd(gnd), .vdd(vdd), .A(_3106_), .Y(_3106__bF_buf4) );
BUFX4 BUFX4_184 ( .gnd(gnd), .vdd(vdd), .A(_3106_), .Y(_3106__bF_buf3) );
BUFX4 BUFX4_185 ( .gnd(gnd), .vdd(vdd), .A(_3106_), .Y(_3106__bF_buf2) );
BUFX4 BUFX4_186 ( .gnd(gnd), .vdd(vdd), .A(_3106_), .Y(_3106__bF_buf1) );
BUFX4 BUFX4_187 ( .gnd(gnd), .vdd(vdd), .A(_3106_), .Y(_3106__bF_buf0) );
BUFX4 BUFX4_188 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_0_), .Y(micro_hash_ucr_c_0_bF_buf3_) );
BUFX4 BUFX4_189 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_0_), .Y(micro_hash_ucr_c_0_bF_buf2_) );
BUFX4 BUFX4_190 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_0_), .Y(micro_hash_ucr_c_0_bF_buf1_) );
BUFX4 BUFX4_191 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_0_), .Y(micro_hash_ucr_c_0_bF_buf0_) );
BUFX4 BUFX4_192 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_3_), .Y(micro_hash_ucr_b_3_bF_buf3_) );
BUFX4 BUFX4_193 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_3_), .Y(micro_hash_ucr_b_3_bF_buf2_) );
BUFX4 BUFX4_194 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_3_), .Y(micro_hash_ucr_b_3_bF_buf1_) );
BUFX4 BUFX4_195 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_3_), .Y(micro_hash_ucr_b_3_bF_buf0_) );
BUFX4 BUFX4_196 ( .gnd(gnd), .vdd(vdd), .A(_7776_), .Y(_7776__bF_buf4) );
BUFX4 BUFX4_197 ( .gnd(gnd), .vdd(vdd), .A(_7776_), .Y(_7776__bF_buf3) );
BUFX4 BUFX4_198 ( .gnd(gnd), .vdd(vdd), .A(_7776_), .Y(_7776__bF_buf2) );
BUFX4 BUFX4_199 ( .gnd(gnd), .vdd(vdd), .A(_7776_), .Y(_7776__bF_buf1) );
BUFX4 BUFX4_200 ( .gnd(gnd), .vdd(vdd), .A(_7776_), .Y(_7776__bF_buf0) );
BUFX4 BUFX4_201 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_6_), .Y(micro_hash_ucr_a_6_bF_buf3_) );
BUFX4 BUFX4_202 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_6_), .Y(micro_hash_ucr_a_6_bF_buf2_) );
BUFX4 BUFX4_203 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_6_), .Y(micro_hash_ucr_a_6_bF_buf1_) );
BUFX4 BUFX4_204 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_6_), .Y(micro_hash_ucr_a_6_bF_buf0_) );
BUFX4 BUFX4_205 ( .gnd(gnd), .vdd(vdd), .A(_9311_), .Y(_9311__bF_buf4) );
BUFX4 BUFX4_206 ( .gnd(gnd), .vdd(vdd), .A(_9311_), .Y(_9311__bF_buf3) );
BUFX4 BUFX4_207 ( .gnd(gnd), .vdd(vdd), .A(_9311_), .Y(_9311__bF_buf2) );
BUFX4 BUFX4_208 ( .gnd(gnd), .vdd(vdd), .A(_9311_), .Y(_9311__bF_buf1) );
BUFX4 BUFX4_209 ( .gnd(gnd), .vdd(vdd), .A(_9311_), .Y(_9311__bF_buf0) );
BUFX4 BUFX4_210 ( .gnd(gnd), .vdd(vdd), .A(_899_), .Y(_899__bF_buf3) );
BUFX4 BUFX4_211 ( .gnd(gnd), .vdd(vdd), .A(_899_), .Y(_899__bF_buf2) );
BUFX4 BUFX4_212 ( .gnd(gnd), .vdd(vdd), .A(_899_), .Y(_899__bF_buf1) );
BUFX4 BUFX4_213 ( .gnd(gnd), .vdd(vdd), .A(_899_), .Y(_899__bF_buf0) );
BUFX4 BUFX4_214 ( .gnd(gnd), .vdd(vdd), .A(_9290_), .Y(_9290__bF_buf3) );
BUFX4 BUFX4_215 ( .gnd(gnd), .vdd(vdd), .A(_9290_), .Y(_9290__bF_buf2) );
BUFX4 BUFX4_216 ( .gnd(gnd), .vdd(vdd), .A(_9290_), .Y(_9290__bF_buf1) );
BUFX4 BUFX4_217 ( .gnd(gnd), .vdd(vdd), .A(_9290_), .Y(_9290__bF_buf0) );
BUFX4 BUFX4_218 ( .gnd(gnd), .vdd(vdd), .A(_920_), .Y(_920__bF_buf4) );
BUFX4 BUFX4_219 ( .gnd(gnd), .vdd(vdd), .A(_920_), .Y(_920__bF_buf3) );
BUFX4 BUFX4_220 ( .gnd(gnd), .vdd(vdd), .A(_920_), .Y(_920__bF_buf2) );
BUFX4 BUFX4_221 ( .gnd(gnd), .vdd(vdd), .A(_920_), .Y(_920__bF_buf1) );
BUFX4 BUFX4_222 ( .gnd(gnd), .vdd(vdd), .A(_920_), .Y(_920__bF_buf0) );
BUFX4 BUFX4_223 ( .gnd(gnd), .vdd(vdd), .A(_5075_), .Y(_5075__bF_buf4) );
BUFX4 BUFX4_224 ( .gnd(gnd), .vdd(vdd), .A(_5075_), .Y(_5075__bF_buf3) );
BUFX4 BUFX4_225 ( .gnd(gnd), .vdd(vdd), .A(_5075_), .Y(_5075__bF_buf2) );
BUFX4 BUFX4_226 ( .gnd(gnd), .vdd(vdd), .A(_5075_), .Y(_5075__bF_buf1) );
BUFX4 BUFX4_227 ( .gnd(gnd), .vdd(vdd), .A(_5075_), .Y(_5075__bF_buf0) );
BUFX4 BUFX4_228 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_0_), .Y(micro_hash_ucr_b_0_bF_buf3_) );
BUFX4 BUFX4_229 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_0_), .Y(micro_hash_ucr_b_0_bF_buf2_) );
BUFX4 BUFX4_230 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_0_), .Y(micro_hash_ucr_b_0_bF_buf1_) );
BUFX4 BUFX4_231 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_0_), .Y(micro_hash_ucr_b_0_bF_buf0_) );
BUFX4 BUFX4_232 ( .gnd(gnd), .vdd(vdd), .A(_7315_), .Y(_7315__bF_buf5) );
BUFX4 BUFX4_233 ( .gnd(gnd), .vdd(vdd), .A(_7315_), .Y(_7315__bF_buf4) );
BUFX4 BUFX4_234 ( .gnd(gnd), .vdd(vdd), .A(_7315_), .Y(_7315__bF_buf3) );
BUFX4 BUFX4_235 ( .gnd(gnd), .vdd(vdd), .A(_7315_), .Y(_7315__bF_buf2) );
BUFX4 BUFX4_236 ( .gnd(gnd), .vdd(vdd), .A(_7315_), .Y(_7315__bF_buf1) );
BUFX4 BUFX4_237 ( .gnd(gnd), .vdd(vdd), .A(_7315_), .Y(_7315__bF_buf0) );
BUFX4 BUFX4_238 ( .gnd(gnd), .vdd(vdd), .A(_1721_), .Y(_1721__bF_buf4) );
BUFX4 BUFX4_239 ( .gnd(gnd), .vdd(vdd), .A(_1721_), .Y(_1721__bF_buf3) );
BUFX4 BUFX4_240 ( .gnd(gnd), .vdd(vdd), .A(_1721_), .Y(_1721__bF_buf2) );
BUFX4 BUFX4_241 ( .gnd(gnd), .vdd(vdd), .A(_1721_), .Y(_1721__bF_buf1) );
BUFX4 BUFX4_242 ( .gnd(gnd), .vdd(vdd), .A(_1721_), .Y(_1721__bF_buf0) );
BUFX4 BUFX4_243 ( .gnd(gnd), .vdd(vdd), .A(_9287_), .Y(_9287__bF_buf4) );
BUFX4 BUFX4_244 ( .gnd(gnd), .vdd(vdd), .A(_9287_), .Y(_9287__bF_buf3) );
BUFX4 BUFX4_245 ( .gnd(gnd), .vdd(vdd), .A(_9287_), .Y(_9287__bF_buf2) );
BUFX4 BUFX4_246 ( .gnd(gnd), .vdd(vdd), .A(_9287_), .Y(_9287__bF_buf1) );
BUFX4 BUFX4_247 ( .gnd(gnd), .vdd(vdd), .A(_9287_), .Y(_9287__bF_buf0) );
BUFX4 BUFX4_248 ( .gnd(gnd), .vdd(vdd), .A(_12900_), .Y(_12900__bF_buf3) );
BUFX4 BUFX4_249 ( .gnd(gnd), .vdd(vdd), .A(_12900_), .Y(_12900__bF_buf2) );
BUFX4 BUFX4_250 ( .gnd(gnd), .vdd(vdd), .A(_12900_), .Y(_12900__bF_buf1) );
BUFX4 BUFX4_251 ( .gnd(gnd), .vdd(vdd), .A(_12900_), .Y(_12900__bF_buf0) );
BUFX4 BUFX4_252 ( .gnd(gnd), .vdd(vdd), .A(_9305_), .Y(_9305__bF_buf4) );
BUFX4 BUFX4_253 ( .gnd(gnd), .vdd(vdd), .A(_9305_), .Y(_9305__bF_buf3) );
BUFX4 BUFX4_254 ( .gnd(gnd), .vdd(vdd), .A(_9305_), .Y(_9305__bF_buf2) );
BUFX4 BUFX4_255 ( .gnd(gnd), .vdd(vdd), .A(_9305_), .Y(_9305__bF_buf1) );
BUFX4 BUFX4_256 ( .gnd(gnd), .vdd(vdd), .A(_9305_), .Y(_9305__bF_buf0) );
BUFX4 BUFX4_257 ( .gnd(gnd), .vdd(vdd), .A(_896_), .Y(_896__bF_buf4) );
BUFX4 BUFX4_258 ( .gnd(gnd), .vdd(vdd), .A(_896_), .Y(_896__bF_buf3) );
BUFX4 BUFX4_259 ( .gnd(gnd), .vdd(vdd), .A(_896_), .Y(_896__bF_buf2) );
BUFX4 BUFX4_260 ( .gnd(gnd), .vdd(vdd), .A(_896_), .Y(_896__bF_buf1) );
BUFX4 BUFX4_261 ( .gnd(gnd), .vdd(vdd), .A(_896_), .Y(_896__bF_buf0) );
BUFX4 BUFX4_262 ( .gnd(gnd), .vdd(vdd), .A(_12001_), .Y(_12001__bF_buf4) );
BUFX4 BUFX4_263 ( .gnd(gnd), .vdd(vdd), .A(_12001_), .Y(_12001__bF_buf3) );
BUFX4 BUFX4_264 ( .gnd(gnd), .vdd(vdd), .A(_12001_), .Y(_12001__bF_buf2) );
BUFX4 BUFX4_265 ( .gnd(gnd), .vdd(vdd), .A(_12001_), .Y(_12001__bF_buf1) );
BUFX4 BUFX4_266 ( .gnd(gnd), .vdd(vdd), .A(_12001_), .Y(_12001__bF_buf0) );
BUFX4 BUFX4_267 ( .gnd(gnd), .vdd(vdd), .A(_400_), .Y(_400__bF_buf12) );
BUFX4 BUFX4_268 ( .gnd(gnd), .vdd(vdd), .A(_400_), .Y(_400__bF_buf11) );
BUFX4 BUFX4_269 ( .gnd(gnd), .vdd(vdd), .A(_400_), .Y(_400__bF_buf10) );
BUFX4 BUFX4_270 ( .gnd(gnd), .vdd(vdd), .A(_400_), .Y(_400__bF_buf9) );
BUFX4 BUFX4_271 ( .gnd(gnd), .vdd(vdd), .A(_400_), .Y(_400__bF_buf8) );
BUFX4 BUFX4_272 ( .gnd(gnd), .vdd(vdd), .A(_400_), .Y(_400__bF_buf7) );
BUFX4 BUFX4_273 ( .gnd(gnd), .vdd(vdd), .A(_400_), .Y(_400__bF_buf6) );
BUFX4 BUFX4_274 ( .gnd(gnd), .vdd(vdd), .A(_400_), .Y(_400__bF_buf5) );
BUFX4 BUFX4_275 ( .gnd(gnd), .vdd(vdd), .A(_400_), .Y(_400__bF_buf4) );
BUFX4 BUFX4_276 ( .gnd(gnd), .vdd(vdd), .A(_400_), .Y(_400__bF_buf3) );
BUFX4 BUFX4_277 ( .gnd(gnd), .vdd(vdd), .A(_400_), .Y(_400__bF_buf2) );
BUFX4 BUFX4_278 ( .gnd(gnd), .vdd(vdd), .A(_400_), .Y(_400__bF_buf1) );
BUFX4 BUFX4_279 ( .gnd(gnd), .vdd(vdd), .A(_400_), .Y(_400__bF_buf0) );
BUFX4 BUFX4_280 ( .gnd(gnd), .vdd(vdd), .A(_914_), .Y(_914__bF_buf4) );
BUFX4 BUFX4_281 ( .gnd(gnd), .vdd(vdd), .A(_914_), .Y(_914__bF_buf3) );
BUFX4 BUFX4_282 ( .gnd(gnd), .vdd(vdd), .A(_914_), .Y(_914__bF_buf2) );
BUFX4 BUFX4_283 ( .gnd(gnd), .vdd(vdd), .A(_914_), .Y(_914__bF_buf1) );
BUFX4 BUFX4_284 ( .gnd(gnd), .vdd(vdd), .A(_914_), .Y(_914__bF_buf0) );
BUFX4 BUFX4_285 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_0_), .Y(micro_hash_ucr_a_0_bF_buf3_) );
BUFX4 BUFX4_286 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_0_), .Y(micro_hash_ucr_a_0_bF_buf2_) );
BUFX4 BUFX4_287 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_0_), .Y(micro_hash_ucr_a_0_bF_buf1_) );
BUFX4 BUFX4_288 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_0_), .Y(micro_hash_ucr_a_0_bF_buf0_) );
CLKBUF1 CLKBUF1_1 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf11), .Y(clk_bF_buf157) );
CLKBUF1 CLKBUF1_2 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf10), .Y(clk_bF_buf156) );
CLKBUF1 CLKBUF1_3 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf155) );
CLKBUF1 CLKBUF1_4 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf154) );
CLKBUF1 CLKBUF1_5 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf153) );
CLKBUF1 CLKBUF1_6 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf152) );
CLKBUF1 CLKBUF1_7 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf151) );
CLKBUF1 CLKBUF1_8 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf150) );
CLKBUF1 CLKBUF1_9 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf149) );
CLKBUF1 CLKBUF1_10 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf148) );
CLKBUF1 CLKBUF1_11 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf147) );
CLKBUF1 CLKBUF1_12 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf146) );
CLKBUF1 CLKBUF1_13 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf11), .Y(clk_bF_buf145) );
CLKBUF1 CLKBUF1_14 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf10), .Y(clk_bF_buf144) );
CLKBUF1 CLKBUF1_15 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf143) );
CLKBUF1 CLKBUF1_16 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf142) );
CLKBUF1 CLKBUF1_17 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf141) );
CLKBUF1 CLKBUF1_18 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf140) );
CLKBUF1 CLKBUF1_19 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf139) );
CLKBUF1 CLKBUF1_20 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf138) );
CLKBUF1 CLKBUF1_21 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf137) );
CLKBUF1 CLKBUF1_22 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf136) );
CLKBUF1 CLKBUF1_23 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf135) );
CLKBUF1 CLKBUF1_24 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf134) );
CLKBUF1 CLKBUF1_25 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf11), .Y(clk_bF_buf133) );
CLKBUF1 CLKBUF1_26 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf10), .Y(clk_bF_buf132) );
CLKBUF1 CLKBUF1_27 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf131) );
CLKBUF1 CLKBUF1_28 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf130) );
CLKBUF1 CLKBUF1_29 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf129) );
CLKBUF1 CLKBUF1_30 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf128) );
CLKBUF1 CLKBUF1_31 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf127) );
CLKBUF1 CLKBUF1_32 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf126) );
CLKBUF1 CLKBUF1_33 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf125) );
CLKBUF1 CLKBUF1_34 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf124) );
CLKBUF1 CLKBUF1_35 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf123) );
CLKBUF1 CLKBUF1_36 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf122) );
CLKBUF1 CLKBUF1_37 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf11), .Y(clk_bF_buf121) );
CLKBUF1 CLKBUF1_38 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf10), .Y(clk_bF_buf120) );
CLKBUF1 CLKBUF1_39 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf119) );
CLKBUF1 CLKBUF1_40 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf118) );
CLKBUF1 CLKBUF1_41 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf117) );
CLKBUF1 CLKBUF1_42 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf116) );
CLKBUF1 CLKBUF1_43 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf115) );
CLKBUF1 CLKBUF1_44 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf114) );
CLKBUF1 CLKBUF1_45 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf113) );
CLKBUF1 CLKBUF1_46 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf112) );
CLKBUF1 CLKBUF1_47 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf111) );
CLKBUF1 CLKBUF1_48 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf110) );
CLKBUF1 CLKBUF1_49 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf11), .Y(clk_bF_buf109) );
CLKBUF1 CLKBUF1_50 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf10), .Y(clk_bF_buf108) );
CLKBUF1 CLKBUF1_51 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf107) );
CLKBUF1 CLKBUF1_52 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf106) );
CLKBUF1 CLKBUF1_53 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf105) );
CLKBUF1 CLKBUF1_54 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf104) );
CLKBUF1 CLKBUF1_55 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf103) );
CLKBUF1 CLKBUF1_56 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf102) );
CLKBUF1 CLKBUF1_57 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf101) );
CLKBUF1 CLKBUF1_58 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf100) );
CLKBUF1 CLKBUF1_59 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf99) );
CLKBUF1 CLKBUF1_60 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf98) );
CLKBUF1 CLKBUF1_61 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf11), .Y(clk_bF_buf97) );
CLKBUF1 CLKBUF1_62 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf10), .Y(clk_bF_buf96) );
CLKBUF1 CLKBUF1_63 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf95) );
CLKBUF1 CLKBUF1_64 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf94) );
CLKBUF1 CLKBUF1_65 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf93) );
CLKBUF1 CLKBUF1_66 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf92) );
CLKBUF1 CLKBUF1_67 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf91) );
CLKBUF1 CLKBUF1_68 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf90) );
CLKBUF1 CLKBUF1_69 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf89) );
CLKBUF1 CLKBUF1_70 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf88) );
CLKBUF1 CLKBUF1_71 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf87) );
CLKBUF1 CLKBUF1_72 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf86) );
CLKBUF1 CLKBUF1_73 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf11), .Y(clk_bF_buf85) );
CLKBUF1 CLKBUF1_74 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf10), .Y(clk_bF_buf84) );
CLKBUF1 CLKBUF1_75 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf83) );
CLKBUF1 CLKBUF1_76 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf82) );
CLKBUF1 CLKBUF1_77 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf81) );
CLKBUF1 CLKBUF1_78 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf80) );
CLKBUF1 CLKBUF1_79 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf79) );
CLKBUF1 CLKBUF1_80 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf78) );
CLKBUF1 CLKBUF1_81 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf77) );
CLKBUF1 CLKBUF1_82 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf76) );
CLKBUF1 CLKBUF1_83 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf75) );
CLKBUF1 CLKBUF1_84 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf74) );
CLKBUF1 CLKBUF1_85 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf11), .Y(clk_bF_buf73) );
CLKBUF1 CLKBUF1_86 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf10), .Y(clk_bF_buf72) );
CLKBUF1 CLKBUF1_87 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf71) );
CLKBUF1 CLKBUF1_88 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf70) );
CLKBUF1 CLKBUF1_89 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf69) );
CLKBUF1 CLKBUF1_90 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf68) );
CLKBUF1 CLKBUF1_91 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf67) );
CLKBUF1 CLKBUF1_92 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf66) );
CLKBUF1 CLKBUF1_93 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf65) );
CLKBUF1 CLKBUF1_94 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf64) );
CLKBUF1 CLKBUF1_95 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf63) );
CLKBUF1 CLKBUF1_96 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf62) );
CLKBUF1 CLKBUF1_97 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf11), .Y(clk_bF_buf61) );
CLKBUF1 CLKBUF1_98 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf10), .Y(clk_bF_buf60) );
CLKBUF1 CLKBUF1_99 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf59) );
CLKBUF1 CLKBUF1_100 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf58) );
CLKBUF1 CLKBUF1_101 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf57) );
CLKBUF1 CLKBUF1_102 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf56) );
CLKBUF1 CLKBUF1_103 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf55) );
CLKBUF1 CLKBUF1_104 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf54) );
CLKBUF1 CLKBUF1_105 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf53) );
CLKBUF1 CLKBUF1_106 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf52) );
CLKBUF1 CLKBUF1_107 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf51) );
CLKBUF1 CLKBUF1_108 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf50) );
CLKBUF1 CLKBUF1_109 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf11), .Y(clk_bF_buf49) );
CLKBUF1 CLKBUF1_110 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf10), .Y(clk_bF_buf48) );
CLKBUF1 CLKBUF1_111 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf47) );
CLKBUF1 CLKBUF1_112 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf46) );
CLKBUF1 CLKBUF1_113 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf45) );
CLKBUF1 CLKBUF1_114 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf44) );
CLKBUF1 CLKBUF1_115 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf43) );
CLKBUF1 CLKBUF1_116 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf42) );
CLKBUF1 CLKBUF1_117 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf41) );
CLKBUF1 CLKBUF1_118 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf40) );
CLKBUF1 CLKBUF1_119 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf39) );
CLKBUF1 CLKBUF1_120 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf38) );
CLKBUF1 CLKBUF1_121 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf11), .Y(clk_bF_buf37) );
CLKBUF1 CLKBUF1_122 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf10), .Y(clk_bF_buf36) );
CLKBUF1 CLKBUF1_123 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf35) );
CLKBUF1 CLKBUF1_124 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf34) );
CLKBUF1 CLKBUF1_125 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf33) );
CLKBUF1 CLKBUF1_126 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf32) );
CLKBUF1 CLKBUF1_127 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf31) );
CLKBUF1 CLKBUF1_128 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf30) );
CLKBUF1 CLKBUF1_129 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf29) );
CLKBUF1 CLKBUF1_130 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf28) );
CLKBUF1 CLKBUF1_131 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf27) );
CLKBUF1 CLKBUF1_132 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf26) );
CLKBUF1 CLKBUF1_133 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf11), .Y(clk_bF_buf25) );
CLKBUF1 CLKBUF1_134 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf10), .Y(clk_bF_buf24) );
CLKBUF1 CLKBUF1_135 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf23) );
CLKBUF1 CLKBUF1_136 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf22) );
CLKBUF1 CLKBUF1_137 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf21) );
CLKBUF1 CLKBUF1_138 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf20) );
CLKBUF1 CLKBUF1_139 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf19) );
CLKBUF1 CLKBUF1_140 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf18) );
CLKBUF1 CLKBUF1_141 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf17) );
CLKBUF1 CLKBUF1_142 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf16) );
CLKBUF1 CLKBUF1_143 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf15) );
CLKBUF1 CLKBUF1_144 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf14) );
CLKBUF1 CLKBUF1_145 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf11), .Y(clk_bF_buf13) );
CLKBUF1 CLKBUF1_146 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf10), .Y(clk_bF_buf12) );
CLKBUF1 CLKBUF1_147 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf11) );
CLKBUF1 CLKBUF1_148 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf10) );
CLKBUF1 CLKBUF1_149 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf9) );
CLKBUF1 CLKBUF1_150 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf8) );
CLKBUF1 CLKBUF1_151 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf7) );
CLKBUF1 CLKBUF1_152 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf6) );
CLKBUF1 CLKBUF1_153 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf5) );
CLKBUF1 CLKBUF1_154 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf4) );
CLKBUF1 CLKBUF1_155 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf3) );
CLKBUF1 CLKBUF1_156 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf2) );
CLKBUF1 CLKBUF1_157 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf11), .Y(clk_bF_buf1) );
CLKBUF1 CLKBUF1_158 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf10), .Y(clk_bF_buf0) );
BUFX4 BUFX4_289 ( .gnd(gnd), .vdd(vdd), .A(_10522_), .Y(_10522__bF_buf4) );
BUFX4 BUFX4_290 ( .gnd(gnd), .vdd(vdd), .A(_10522_), .Y(_10522__bF_buf3) );
BUFX4 BUFX4_291 ( .gnd(gnd), .vdd(vdd), .A(_10522_), .Y(_10522__bF_buf2) );
BUFX4 BUFX4_292 ( .gnd(gnd), .vdd(vdd), .A(_10522_), .Y(_10522__bF_buf1) );
BUFX4 BUFX4_293 ( .gnd(gnd), .vdd(vdd), .A(_10522_), .Y(_10522__bF_buf0) );
BUFX4 BUFX4_294 ( .gnd(gnd), .vdd(vdd), .A(_11536_), .Y(_11536__bF_buf3) );
BUFX4 BUFX4_295 ( .gnd(gnd), .vdd(vdd), .A(_11536_), .Y(_11536__bF_buf2) );
BUFX4 BUFX4_296 ( .gnd(gnd), .vdd(vdd), .A(_11536_), .Y(_11536__bF_buf1) );
BUFX4 BUFX4_297 ( .gnd(gnd), .vdd(vdd), .A(_11536_), .Y(_11536__bF_buf0) );
BUFX4 BUFX4_298 ( .gnd(gnd), .vdd(vdd), .A(_10519_), .Y(_10519__bF_buf5) );
BUFX4 BUFX4_299 ( .gnd(gnd), .vdd(vdd), .A(_10519_), .Y(_10519__bF_buf4) );
BUFX4 BUFX4_300 ( .gnd(gnd), .vdd(vdd), .A(_10519_), .Y(_10519__bF_buf3) );
BUFX4 BUFX4_301 ( .gnd(gnd), .vdd(vdd), .A(_10519_), .Y(_10519__bF_buf2) );
BUFX4 BUFX4_302 ( .gnd(gnd), .vdd(vdd), .A(_10519_), .Y(_10519__bF_buf1) );
BUFX4 BUFX4_303 ( .gnd(gnd), .vdd(vdd), .A(_10519_), .Y(_10519__bF_buf0) );
BUFX4 BUFX4_304 ( .gnd(gnd), .vdd(vdd), .A(_5125_), .Y(_5125__bF_buf3) );
BUFX4 BUFX4_305 ( .gnd(gnd), .vdd(vdd), .A(_5125_), .Y(_5125__bF_buf2) );
BUFX4 BUFX4_306 ( .gnd(gnd), .vdd(vdd), .A(_5125_), .Y(_5125__bF_buf1) );
BUFX4 BUFX4_307 ( .gnd(gnd), .vdd(vdd), .A(_5125_), .Y(_5125__bF_buf0) );
BUFX4 BUFX4_308 ( .gnd(gnd), .vdd(vdd), .A(_8705_), .Y(_8705__bF_buf13) );
BUFX4 BUFX4_309 ( .gnd(gnd), .vdd(vdd), .A(_8705_), .Y(_8705__bF_buf12) );
BUFX4 BUFX4_310 ( .gnd(gnd), .vdd(vdd), .A(_8705_), .Y(_8705__bF_buf11) );
BUFX4 BUFX4_311 ( .gnd(gnd), .vdd(vdd), .A(_8705_), .Y(_8705__bF_buf10) );
BUFX4 BUFX4_312 ( .gnd(gnd), .vdd(vdd), .A(_8705_), .Y(_8705__bF_buf9) );
BUFX4 BUFX4_313 ( .gnd(gnd), .vdd(vdd), .A(_8705_), .Y(_8705__bF_buf8) );
BUFX4 BUFX4_314 ( .gnd(gnd), .vdd(vdd), .A(_8705_), .Y(_8705__bF_buf7) );
BUFX4 BUFX4_315 ( .gnd(gnd), .vdd(vdd), .A(_8705_), .Y(_8705__bF_buf6) );
BUFX4 BUFX4_316 ( .gnd(gnd), .vdd(vdd), .A(_8705_), .Y(_8705__bF_buf5) );
BUFX4 BUFX4_317 ( .gnd(gnd), .vdd(vdd), .A(_8705_), .Y(_8705__bF_buf4) );
BUFX4 BUFX4_318 ( .gnd(gnd), .vdd(vdd), .A(_8705_), .Y(_8705__bF_buf3) );
BUFX4 BUFX4_319 ( .gnd(gnd), .vdd(vdd), .A(_8705_), .Y(_8705__bF_buf2) );
BUFX4 BUFX4_320 ( .gnd(gnd), .vdd(vdd), .A(_8705_), .Y(_8705__bF_buf1) );
BUFX4 BUFX4_321 ( .gnd(gnd), .vdd(vdd), .A(_8705_), .Y(_8705__bF_buf0) );
BUFX4 BUFX4_322 ( .gnd(gnd), .vdd(vdd), .A(_911_), .Y(_911__bF_buf4) );
BUFX4 BUFX4_323 ( .gnd(gnd), .vdd(vdd), .A(_911_), .Y(_911__bF_buf3) );
BUFX4 BUFX4_324 ( .gnd(gnd), .vdd(vdd), .A(_911_), .Y(_911__bF_buf2) );
BUFX4 BUFX4_325 ( .gnd(gnd), .vdd(vdd), .A(_911_), .Y(_911__bF_buf1) );
BUFX4 BUFX4_326 ( .gnd(gnd), .vdd(vdd), .A(_911_), .Y(_911__bF_buf0) );
BUFX4 BUFX4_327 ( .gnd(gnd), .vdd(vdd), .A(_2306_), .Y(_2306__bF_buf3) );
BUFX4 BUFX4_328 ( .gnd(gnd), .vdd(vdd), .A(_2306_), .Y(_2306__bF_buf2) );
BUFX4 BUFX4_329 ( .gnd(gnd), .vdd(vdd), .A(_2306_), .Y(_2306__bF_buf1) );
BUFX4 BUFX4_330 ( .gnd(gnd), .vdd(vdd), .A(_2306_), .Y(_2306__bF_buf0) );
BUFX4 BUFX4_331 ( .gnd(gnd), .vdd(vdd), .A(_908_), .Y(_908__bF_buf4) );
BUFX4 BUFX4_332 ( .gnd(gnd), .vdd(vdd), .A(_908_), .Y(_908__bF_buf3) );
BUFX4 BUFX4_333 ( .gnd(gnd), .vdd(vdd), .A(_908_), .Y(_908__bF_buf2) );
BUFX4 BUFX4_334 ( .gnd(gnd), .vdd(vdd), .A(_908_), .Y(_908__bF_buf1) );
BUFX4 BUFX4_335 ( .gnd(gnd), .vdd(vdd), .A(_908_), .Y(_908__bF_buf0) );
BUFX4 BUFX4_336 ( .gnd(gnd), .vdd(vdd), .A(_890_), .Y(_890__bF_buf4) );
BUFX4 BUFX4_337 ( .gnd(gnd), .vdd(vdd), .A(_890_), .Y(_890__bF_buf3) );
BUFX4 BUFX4_338 ( .gnd(gnd), .vdd(vdd), .A(_890_), .Y(_890__bF_buf2) );
BUFX4 BUFX4_339 ( .gnd(gnd), .vdd(vdd), .A(_890_), .Y(_890__bF_buf1) );
BUFX4 BUFX4_340 ( .gnd(gnd), .vdd(vdd), .A(_890_), .Y(_890__bF_buf0) );
BUFX4 BUFX4_341 ( .gnd(gnd), .vdd(vdd), .A(finished_1), .Y(finished_1_bF_buf4) );
BUFX4 BUFX4_342 ( .gnd(gnd), .vdd(vdd), .A(finished_1), .Y(finished_1_bF_buf3) );
BUFX4 BUFX4_343 ( .gnd(gnd), .vdd(vdd), .A(finished_1), .Y(finished_1_bF_buf2) );
BUFX4 BUFX4_344 ( .gnd(gnd), .vdd(vdd), .A(finished_1), .Y(finished_1_bF_buf1) );
BUFX4 BUFX4_345 ( .gnd(gnd), .vdd(vdd), .A(finished_1), .Y(finished_1_bF_buf0) );
BUFX4 BUFX4_346 ( .gnd(gnd), .vdd(vdd), .A(finished_2), .Y(finished_2_bF_buf4) );
BUFX4 BUFX4_347 ( .gnd(gnd), .vdd(vdd), .A(finished_2), .Y(finished_2_bF_buf3) );
BUFX4 BUFX4_348 ( .gnd(gnd), .vdd(vdd), .A(finished_2), .Y(finished_2_bF_buf2) );
BUFX4 BUFX4_349 ( .gnd(gnd), .vdd(vdd), .A(finished_2), .Y(finished_2_bF_buf1) );
BUFX4 BUFX4_350 ( .gnd(gnd), .vdd(vdd), .A(finished_2), .Y(finished_2_bF_buf0) );
BUFX4 BUFX4_351 ( .gnd(gnd), .vdd(vdd), .A(finished_3), .Y(finished_3_bF_buf4) );
BUFX4 BUFX4_352 ( .gnd(gnd), .vdd(vdd), .A(finished_3), .Y(finished_3_bF_buf3) );
BUFX4 BUFX4_353 ( .gnd(gnd), .vdd(vdd), .A(finished_3), .Y(finished_3_bF_buf2) );
BUFX4 BUFX4_354 ( .gnd(gnd), .vdd(vdd), .A(finished_3), .Y(finished_3_bF_buf1) );
BUFX4 BUFX4_355 ( .gnd(gnd), .vdd(vdd), .A(finished_3), .Y(finished_3_bF_buf0) );
BUFX4 BUFX4_356 ( .gnd(gnd), .vdd(vdd), .A(_5122_), .Y(_5122__bF_buf4) );
BUFX4 BUFX4_357 ( .gnd(gnd), .vdd(vdd), .A(_5122_), .Y(_5122__bF_buf3) );
BUFX4 BUFX4_358 ( .gnd(gnd), .vdd(vdd), .A(_5122_), .Y(_5122__bF_buf2) );
BUFX4 BUFX4_359 ( .gnd(gnd), .vdd(vdd), .A(_5122_), .Y(_5122__bF_buf1) );
BUFX4 BUFX4_360 ( .gnd(gnd), .vdd(vdd), .A(_5122_), .Y(_5122__bF_buf0) );
BUFX4 BUFX4_361 ( .gnd(gnd), .vdd(vdd), .A(_11283_), .Y(_11283__bF_buf5) );
BUFX4 BUFX4_362 ( .gnd(gnd), .vdd(vdd), .A(_11283_), .Y(_11283__bF_buf4) );
BUFX4 BUFX4_363 ( .gnd(gnd), .vdd(vdd), .A(_11283_), .Y(_11283__bF_buf3) );
BUFX4 BUFX4_364 ( .gnd(gnd), .vdd(vdd), .A(_11283_), .Y(_11283__bF_buf2) );
BUFX4 BUFX4_365 ( .gnd(gnd), .vdd(vdd), .A(_11283_), .Y(_11283__bF_buf1) );
BUFX4 BUFX4_366 ( .gnd(gnd), .vdd(vdd), .A(_11283_), .Y(_11283__bF_buf0) );
BUFX4 BUFX4_367 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe50), .Y(micro_hash_ucr_2_pipe50_bF_buf3) );
BUFX4 BUFX4_368 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe50), .Y(micro_hash_ucr_2_pipe50_bF_buf2) );
BUFX4 BUFX4_369 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe50), .Y(micro_hash_ucr_2_pipe50_bF_buf1) );
BUFX4 BUFX4_370 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe50), .Y(micro_hash_ucr_2_pipe50_bF_buf0) );
BUFX4 BUFX4_371 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe52), .Y(micro_hash_ucr_2_pipe52_bF_buf3) );
BUFX4 BUFX4_372 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe52), .Y(micro_hash_ucr_2_pipe52_bF_buf2) );
BUFX4 BUFX4_373 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe52), .Y(micro_hash_ucr_2_pipe52_bF_buf1) );
BUFX4 BUFX4_374 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe52), .Y(micro_hash_ucr_2_pipe52_bF_buf0) );
BUFX4 BUFX4_375 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe53), .Y(micro_hash_ucr_2_pipe53_bF_buf3) );
BUFX4 BUFX4_376 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe53), .Y(micro_hash_ucr_2_pipe53_bF_buf2) );
BUFX4 BUFX4_377 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe53), .Y(micro_hash_ucr_2_pipe53_bF_buf1) );
BUFX4 BUFX4_378 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe53), .Y(micro_hash_ucr_2_pipe53_bF_buf0) );
BUFX4 BUFX4_379 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe54), .Y(micro_hash_ucr_2_pipe54_bF_buf4) );
BUFX4 BUFX4_380 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe54), .Y(micro_hash_ucr_2_pipe54_bF_buf3) );
BUFX4 BUFX4_381 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe54), .Y(micro_hash_ucr_2_pipe54_bF_buf2) );
BUFX4 BUFX4_382 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe54), .Y(micro_hash_ucr_2_pipe54_bF_buf1) );
BUFX4 BUFX4_383 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe54), .Y(micro_hash_ucr_2_pipe54_bF_buf0) );
BUFX4 BUFX4_384 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe56), .Y(micro_hash_ucr_2_pipe56_bF_buf3) );
BUFX4 BUFX4_385 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe56), .Y(micro_hash_ucr_2_pipe56_bF_buf2) );
BUFX4 BUFX4_386 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe56), .Y(micro_hash_ucr_2_pipe56_bF_buf1) );
BUFX4 BUFX4_387 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe56), .Y(micro_hash_ucr_2_pipe56_bF_buf0) );
BUFX4 BUFX4_388 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe57), .Y(micro_hash_ucr_2_pipe57_bF_buf3) );
BUFX4 BUFX4_389 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe57), .Y(micro_hash_ucr_2_pipe57_bF_buf2) );
BUFX4 BUFX4_390 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe57), .Y(micro_hash_ucr_2_pipe57_bF_buf1) );
BUFX4 BUFX4_391 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe57), .Y(micro_hash_ucr_2_pipe57_bF_buf0) );
BUFX4 BUFX4_392 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe58), .Y(micro_hash_ucr_2_pipe58_bF_buf4) );
BUFX4 BUFX4_393 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe58), .Y(micro_hash_ucr_2_pipe58_bF_buf3) );
BUFX4 BUFX4_394 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe58), .Y(micro_hash_ucr_2_pipe58_bF_buf2) );
BUFX4 BUFX4_395 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe58), .Y(micro_hash_ucr_2_pipe58_bF_buf1) );
BUFX4 BUFX4_396 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe58), .Y(micro_hash_ucr_2_pipe58_bF_buf0) );
BUFX4 BUFX4_397 ( .gnd(gnd), .vdd(vdd), .A(_4622_), .Y(_4622__bF_buf3) );
BUFX4 BUFX4_398 ( .gnd(gnd), .vdd(vdd), .A(_4622_), .Y(_4622__bF_buf2) );
BUFX4 BUFX4_399 ( .gnd(gnd), .vdd(vdd), .A(_4622_), .Y(_4622__bF_buf1) );
BUFX4 BUFX4_400 ( .gnd(gnd), .vdd(vdd), .A(_4622_), .Y(_4622__bF_buf0) );
BUFX4 BUFX4_401 ( .gnd(gnd), .vdd(vdd), .A(_6785_), .Y(_6785__bF_buf4) );
BUFX4 BUFX4_402 ( .gnd(gnd), .vdd(vdd), .A(_6785_), .Y(_6785__bF_buf3) );
BUFX4 BUFX4_403 ( .gnd(gnd), .vdd(vdd), .A(_6785_), .Y(_6785__bF_buf2) );
BUFX4 BUFX4_404 ( .gnd(gnd), .vdd(vdd), .A(_6785_), .Y(_6785__bF_buf1) );
BUFX4 BUFX4_405 ( .gnd(gnd), .vdd(vdd), .A(_6785_), .Y(_6785__bF_buf0) );
BUFX4 BUFX4_406 ( .gnd(gnd), .vdd(vdd), .A(_887_), .Y(_887__bF_buf3) );
BUFX4 BUFX4_407 ( .gnd(gnd), .vdd(vdd), .A(_887_), .Y(_887__bF_buf2) );
BUFX4 BUFX4_408 ( .gnd(gnd), .vdd(vdd), .A(_887_), .Y(_887__bF_buf1) );
BUFX4 BUFX4_409 ( .gnd(gnd), .vdd(vdd), .A(_887_), .Y(_887__bF_buf0) );
BUFX4 BUFX4_410 ( .gnd(gnd), .vdd(vdd), .A(_9334_), .Y(_9334__bF_buf3) );
BUFX4 BUFX4_411 ( .gnd(gnd), .vdd(vdd), .A(_9334_), .Y(_9334__bF_buf2) );
BUFX4 BUFX4_412 ( .gnd(gnd), .vdd(vdd), .A(_9334_), .Y(_9334__bF_buf1) );
BUFX4 BUFX4_413 ( .gnd(gnd), .vdd(vdd), .A(_9334_), .Y(_9334__bF_buf0) );
BUFX4 BUFX4_414 ( .gnd(gnd), .vdd(vdd), .A(_905_), .Y(_905__bF_buf3) );
BUFX4 BUFX4_415 ( .gnd(gnd), .vdd(vdd), .A(_905_), .Y(_905__bF_buf2) );
BUFX4 BUFX4_416 ( .gnd(gnd), .vdd(vdd), .A(_905_), .Y(_905__bF_buf1) );
BUFX4 BUFX4_417 ( .gnd(gnd), .vdd(vdd), .A(_905_), .Y(_905__bF_buf0) );
BUFX4 BUFX4_418 ( .gnd(gnd), .vdd(vdd), .A(_2570_), .Y(_2570__bF_buf4) );
BUFX4 BUFX4_419 ( .gnd(gnd), .vdd(vdd), .A(_2570_), .Y(_2570__bF_buf3) );
BUFX4 BUFX4_420 ( .gnd(gnd), .vdd(vdd), .A(_2570_), .Y(_2570__bF_buf2) );
BUFX4 BUFX4_421 ( .gnd(gnd), .vdd(vdd), .A(_2570_), .Y(_2570__bF_buf1) );
BUFX4 BUFX4_422 ( .gnd(gnd), .vdd(vdd), .A(_2570_), .Y(_2570__bF_buf0) );
BUFX4 BUFX4_423 ( .gnd(gnd), .vdd(vdd), .A(_5921_), .Y(_5921__bF_buf3) );
BUFX4 BUFX4_424 ( .gnd(gnd), .vdd(vdd), .A(_5921_), .Y(_5921__bF_buf2) );
BUFX4 BUFX4_425 ( .gnd(gnd), .vdd(vdd), .A(_5921_), .Y(_5921__bF_buf1) );
BUFX4 BUFX4_426 ( .gnd(gnd), .vdd(vdd), .A(_5921_), .Y(_5921__bF_buf0) );
BUFX4 BUFX4_427 ( .gnd(gnd), .vdd(vdd), .A(_5098_), .Y(_5098__bF_buf4) );
BUFX4 BUFX4_428 ( .gnd(gnd), .vdd(vdd), .A(_5098_), .Y(_5098__bF_buf3) );
BUFX4 BUFX4_429 ( .gnd(gnd), .vdd(vdd), .A(_5098_), .Y(_5098__bF_buf2) );
BUFX4 BUFX4_430 ( .gnd(gnd), .vdd(vdd), .A(_5098_), .Y(_5098__bF_buf1) );
BUFX4 BUFX4_431 ( .gnd(gnd), .vdd(vdd), .A(_5098_), .Y(_5098__bF_buf0) );
BUFX4 BUFX4_432 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe20), .Y(micro_hash_ucr_2_pipe20_bF_buf3) );
BUFX4 BUFX4_433 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe20), .Y(micro_hash_ucr_2_pipe20_bF_buf2) );
BUFX4 BUFX4_434 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe20), .Y(micro_hash_ucr_2_pipe20_bF_buf1) );
BUFX4 BUFX4_435 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe20), .Y(micro_hash_ucr_2_pipe20_bF_buf0) );
BUFX4 BUFX4_436 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe21), .Y(micro_hash_ucr_2_pipe21_bF_buf3) );
BUFX4 BUFX4_437 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe21), .Y(micro_hash_ucr_2_pipe21_bF_buf2) );
BUFX4 BUFX4_438 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe21), .Y(micro_hash_ucr_2_pipe21_bF_buf1) );
BUFX4 BUFX4_439 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe21), .Y(micro_hash_ucr_2_pipe21_bF_buf0) );
BUFX4 BUFX4_440 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe22), .Y(micro_hash_ucr_2_pipe22_bF_buf4) );
BUFX4 BUFX4_441 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe22), .Y(micro_hash_ucr_2_pipe22_bF_buf3) );
BUFX4 BUFX4_442 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe22), .Y(micro_hash_ucr_2_pipe22_bF_buf2) );
BUFX4 BUFX4_443 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe22), .Y(micro_hash_ucr_2_pipe22_bF_buf1) );
BUFX4 BUFX4_444 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe22), .Y(micro_hash_ucr_2_pipe22_bF_buf0) );
BUFX4 BUFX4_445 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe24), .Y(micro_hash_ucr_2_pipe24_bF_buf3) );
BUFX4 BUFX4_446 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe24), .Y(micro_hash_ucr_2_pipe24_bF_buf2) );
BUFX4 BUFX4_447 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe24), .Y(micro_hash_ucr_2_pipe24_bF_buf1) );
BUFX4 BUFX4_448 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe24), .Y(micro_hash_ucr_2_pipe24_bF_buf0) );
BUFX4 BUFX4_449 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe26), .Y(micro_hash_ucr_2_pipe26_bF_buf3) );
BUFX4 BUFX4_450 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe26), .Y(micro_hash_ucr_2_pipe26_bF_buf2) );
BUFX4 BUFX4_451 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe26), .Y(micro_hash_ucr_2_pipe26_bF_buf1) );
BUFX4 BUFX4_452 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe26), .Y(micro_hash_ucr_2_pipe26_bF_buf0) );
BUFX4 BUFX4_453 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe28), .Y(micro_hash_ucr_2_pipe28_bF_buf3) );
BUFX4 BUFX4_454 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe28), .Y(micro_hash_ucr_2_pipe28_bF_buf2) );
BUFX4 BUFX4_455 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe28), .Y(micro_hash_ucr_2_pipe28_bF_buf1) );
BUFX4 BUFX4_456 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe28), .Y(micro_hash_ucr_2_pipe28_bF_buf0) );
BUFX4 BUFX4_457 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe29), .Y(micro_hash_ucr_2_pipe29_bF_buf3) );
BUFX4 BUFX4_458 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe29), .Y(micro_hash_ucr_2_pipe29_bF_buf2) );
BUFX4 BUFX4_459 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe29), .Y(micro_hash_ucr_2_pipe29_bF_buf1) );
BUFX4 BUFX4_460 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe29), .Y(micro_hash_ucr_2_pipe29_bF_buf0) );
BUFX4 BUFX4_461 ( .gnd(gnd), .vdd(vdd), .A(_884_), .Y(_884__bF_buf4) );
BUFX4 BUFX4_462 ( .gnd(gnd), .vdd(vdd), .A(_884_), .Y(_884__bF_buf3) );
BUFX4 BUFX4_463 ( .gnd(gnd), .vdd(vdd), .A(_884_), .Y(_884__bF_buf2) );
BUFX4 BUFX4_464 ( .gnd(gnd), .vdd(vdd), .A(_884_), .Y(_884__bF_buf1) );
BUFX4 BUFX4_465 ( .gnd(gnd), .vdd(vdd), .A(_884_), .Y(_884__bF_buf0) );
BUFX4 BUFX4_466 ( .gnd(gnd), .vdd(vdd), .A(_5116_), .Y(_5116__bF_buf4) );
BUFX4 BUFX4_467 ( .gnd(gnd), .vdd(vdd), .A(_5116_), .Y(_5116__bF_buf3) );
BUFX4 BUFX4_468 ( .gnd(gnd), .vdd(vdd), .A(_5116_), .Y(_5116__bF_buf2) );
BUFX4 BUFX4_469 ( .gnd(gnd), .vdd(vdd), .A(_5116_), .Y(_5116__bF_buf1) );
BUFX4 BUFX4_470 ( .gnd(gnd), .vdd(vdd), .A(_5116_), .Y(_5116__bF_buf0) );
BUFX4 BUFX4_471 ( .gnd(gnd), .vdd(vdd), .A(_10739_), .Y(_10739__bF_buf3) );
BUFX4 BUFX4_472 ( .gnd(gnd), .vdd(vdd), .A(_10739_), .Y(_10739__bF_buf2) );
BUFX4 BUFX4_473 ( .gnd(gnd), .vdd(vdd), .A(_10739_), .Y(_10739__bF_buf1) );
BUFX4 BUFX4_474 ( .gnd(gnd), .vdd(vdd), .A(_10739_), .Y(_10739__bF_buf0) );
BUFX4 BUFX4_475 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_7_), .Y(micro_hash_ucr_2_b_7_bF_buf3_) );
BUFX4 BUFX4_476 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_7_), .Y(micro_hash_ucr_2_b_7_bF_buf2_) );
BUFX4 BUFX4_477 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_7_), .Y(micro_hash_ucr_2_b_7_bF_buf1_) );
BUFX4 BUFX4_478 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_7_), .Y(micro_hash_ucr_2_b_7_bF_buf0_) );
BUFX4 BUFX4_479 ( .gnd(gnd), .vdd(vdd), .A(_4654_), .Y(_4654__bF_buf3) );
BUFX4 BUFX4_480 ( .gnd(gnd), .vdd(vdd), .A(_4654_), .Y(_4654__bF_buf2) );
BUFX4 BUFX4_481 ( .gnd(gnd), .vdd(vdd), .A(_4654_), .Y(_4654__bF_buf1) );
BUFX4 BUFX4_482 ( .gnd(gnd), .vdd(vdd), .A(_4654_), .Y(_4654__bF_buf0) );
BUFX4 BUFX4_483 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe70), .Y(micro_hash_ucr_3_pipe70_bF_buf3) );
BUFX4 BUFX4_484 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe70), .Y(micro_hash_ucr_3_pipe70_bF_buf2) );
BUFX4 BUFX4_485 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe70), .Y(micro_hash_ucr_3_pipe70_bF_buf1) );
BUFX4 BUFX4_486 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe70), .Y(micro_hash_ucr_3_pipe70_bF_buf0) );
BUFX4 BUFX4_487 ( .gnd(gnd), .vdd(vdd), .A(_9328_), .Y(_9328__bF_buf3) );
BUFX4 BUFX4_488 ( .gnd(gnd), .vdd(vdd), .A(_9328_), .Y(_9328__bF_buf2) );
BUFX4 BUFX4_489 ( .gnd(gnd), .vdd(vdd), .A(_9328_), .Y(_9328__bF_buf1) );
BUFX4 BUFX4_490 ( .gnd(gnd), .vdd(vdd), .A(_9328_), .Y(_9328__bF_buf0) );
BUFX4 BUFX4_491 ( .gnd(gnd), .vdd(vdd), .A(_902_), .Y(_902__bF_buf4) );
BUFX4 BUFX4_492 ( .gnd(gnd), .vdd(vdd), .A(_902_), .Y(_902__bF_buf3) );
BUFX4 BUFX4_493 ( .gnd(gnd), .vdd(vdd), .A(_902_), .Y(_902__bF_buf2) );
BUFX4 BUFX4_494 ( .gnd(gnd), .vdd(vdd), .A(_902_), .Y(_902__bF_buf1) );
BUFX4 BUFX4_495 ( .gnd(gnd), .vdd(vdd), .A(_902_), .Y(_902__bF_buf0) );
BUFX4 BUFX4_496 ( .gnd(gnd), .vdd(vdd), .A(_3352_), .Y(_3352__bF_buf4) );
BUFX4 BUFX4_497 ( .gnd(gnd), .vdd(vdd), .A(_3352_), .Y(_3352__bF_buf3) );
BUFX4 BUFX4_498 ( .gnd(gnd), .vdd(vdd), .A(_3352_), .Y(_3352__bF_buf2) );
BUFX4 BUFX4_499 ( .gnd(gnd), .vdd(vdd), .A(_3352_), .Y(_3352__bF_buf1) );
BUFX4 BUFX4_500 ( .gnd(gnd), .vdd(vdd), .A(_3352_), .Y(_3352__bF_buf0) );
BUFX4 BUFX4_501 ( .gnd(gnd), .vdd(vdd), .A(_6512_), .Y(_6512__bF_buf3) );
BUFX4 BUFX4_502 ( .gnd(gnd), .vdd(vdd), .A(_6512_), .Y(_6512__bF_buf2) );
BUFX4 BUFX4_503 ( .gnd(gnd), .vdd(vdd), .A(_6512_), .Y(_6512__bF_buf1) );
BUFX4 BUFX4_504 ( .gnd(gnd), .vdd(vdd), .A(_6512_), .Y(_6512__bF_buf0) );
BUFX4 BUFX4_505 ( .gnd(gnd), .vdd(vdd), .A(_11791_), .Y(_11791__bF_buf5) );
BUFX4 BUFX4_506 ( .gnd(gnd), .vdd(vdd), .A(_11791_), .Y(_11791__bF_buf4) );
BUFX4 BUFX4_507 ( .gnd(gnd), .vdd(vdd), .A(_11791_), .Y(_11791__bF_buf3) );
BUFX4 BUFX4_508 ( .gnd(gnd), .vdd(vdd), .A(_11791_), .Y(_11791__bF_buf2) );
BUFX4 BUFX4_509 ( .gnd(gnd), .vdd(vdd), .A(_11791_), .Y(_11791__bF_buf1) );
BUFX4 BUFX4_510 ( .gnd(gnd), .vdd(vdd), .A(_11791_), .Y(_11791__bF_buf0) );
BUFX4 BUFX4_511 ( .gnd(gnd), .vdd(vdd), .A(comparador_next), .Y(comparador_next_bF_buf3) );
BUFX4 BUFX4_512 ( .gnd(gnd), .vdd(vdd), .A(comparador_next), .Y(comparador_next_bF_buf2) );
BUFX4 BUFX4_513 ( .gnd(gnd), .vdd(vdd), .A(comparador_next), .Y(comparador_next_bF_buf1) );
BUFX4 BUFX4_514 ( .gnd(gnd), .vdd(vdd), .A(comparador_next), .Y(comparador_next_bF_buf0) );
BUFX4 BUFX4_515 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_1_), .Y(micro_hash_ucr_2_c_1_bF_buf3_) );
BUFX4 BUFX4_516 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_1_), .Y(micro_hash_ucr_2_c_1_bF_buf2_) );
BUFX4 BUFX4_517 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_1_), .Y(micro_hash_ucr_2_c_1_bF_buf1_) );
BUFX4 BUFX4_518 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_1_), .Y(micro_hash_ucr_2_c_1_bF_buf0_) );
BUFX4 BUFX4_519 ( .gnd(gnd), .vdd(vdd), .A(_5915_), .Y(_5915__bF_buf3) );
BUFX4 BUFX4_520 ( .gnd(gnd), .vdd(vdd), .A(_5915_), .Y(_5915__bF_buf2) );
BUFX4 BUFX4_521 ( .gnd(gnd), .vdd(vdd), .A(_5915_), .Y(_5915__bF_buf1) );
BUFX4 BUFX4_522 ( .gnd(gnd), .vdd(vdd), .A(_5915_), .Y(_5915__bF_buf0) );
BUFX4 BUFX4_523 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_4_), .Y(micro_hash_ucr_2_b_4_bF_buf3_) );
BUFX4 BUFX4_524 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_4_), .Y(micro_hash_ucr_2_b_4_bF_buf2_) );
BUFX4 BUFX4_525 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_4_), .Y(micro_hash_ucr_2_b_4_bF_buf1_) );
BUFX4 BUFX4_526 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_4_), .Y(micro_hash_ucr_2_b_4_bF_buf0_) );
BUFX4 BUFX4_527 ( .gnd(gnd), .vdd(vdd), .A(_5818_), .Y(_5818__bF_buf3) );
BUFX4 BUFX4_528 ( .gnd(gnd), .vdd(vdd), .A(_5818_), .Y(_5818__bF_buf2) );
BUFX4 BUFX4_529 ( .gnd(gnd), .vdd(vdd), .A(_5818_), .Y(_5818__bF_buf1) );
BUFX4 BUFX4_530 ( .gnd(gnd), .vdd(vdd), .A(_5818_), .Y(_5818__bF_buf0) );
BUFX4 BUFX4_531 ( .gnd(gnd), .vdd(vdd), .A(_5380_), .Y(_5380__bF_buf3) );
BUFX4 BUFX4_532 ( .gnd(gnd), .vdd(vdd), .A(_5380_), .Y(_5380__bF_buf2) );
BUFX4 BUFX4_533 ( .gnd(gnd), .vdd(vdd), .A(_5380_), .Y(_5380__bF_buf1) );
BUFX4 BUFX4_534 ( .gnd(gnd), .vdd(vdd), .A(_5380_), .Y(_5380__bF_buf0) );
BUFX4 BUFX4_535 ( .gnd(gnd), .vdd(vdd), .A(_878_), .Y(_878__bF_buf4) );
BUFX4 BUFX4_536 ( .gnd(gnd), .vdd(vdd), .A(_878_), .Y(_878__bF_buf3) );
BUFX4 BUFX4_537 ( .gnd(gnd), .vdd(vdd), .A(_878_), .Y(_878__bF_buf2) );
BUFX4 BUFX4_538 ( .gnd(gnd), .vdd(vdd), .A(_878_), .Y(_878__bF_buf1) );
BUFX4 BUFX4_539 ( .gnd(gnd), .vdd(vdd), .A(_878_), .Y(_878__bF_buf0) );
BUFX4 BUFX4_540 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe40), .Y(micro_hash_ucr_3_pipe40_bF_buf4) );
BUFX4 BUFX4_541 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe40), .Y(micro_hash_ucr_3_pipe40_bF_buf3) );
BUFX4 BUFX4_542 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe40), .Y(micro_hash_ucr_3_pipe40_bF_buf2) );
BUFX4 BUFX4_543 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe40), .Y(micro_hash_ucr_3_pipe40_bF_buf1) );
BUFX4 BUFX4_544 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe40), .Y(micro_hash_ucr_3_pipe40_bF_buf0) );
BUFX4 BUFX4_545 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe41), .Y(micro_hash_ucr_3_pipe41_bF_buf3) );
BUFX4 BUFX4_546 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe41), .Y(micro_hash_ucr_3_pipe41_bF_buf2) );
BUFX4 BUFX4_547 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe41), .Y(micro_hash_ucr_3_pipe41_bF_buf1) );
BUFX4 BUFX4_548 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe41), .Y(micro_hash_ucr_3_pipe41_bF_buf0) );
BUFX4 BUFX4_549 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe42), .Y(micro_hash_ucr_3_pipe42_bF_buf3) );
BUFX4 BUFX4_550 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe42), .Y(micro_hash_ucr_3_pipe42_bF_buf2) );
BUFX4 BUFX4_551 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe42), .Y(micro_hash_ucr_3_pipe42_bF_buf1) );
BUFX4 BUFX4_552 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe42), .Y(micro_hash_ucr_3_pipe42_bF_buf0) );
BUFX4 BUFX4_553 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe44), .Y(micro_hash_ucr_3_pipe44_bF_buf3) );
BUFX4 BUFX4_554 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe44), .Y(micro_hash_ucr_3_pipe44_bF_buf2) );
BUFX4 BUFX4_555 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe44), .Y(micro_hash_ucr_3_pipe44_bF_buf1) );
BUFX4 BUFX4_556 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe44), .Y(micro_hash_ucr_3_pipe44_bF_buf0) );
BUFX4 BUFX4_557 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe45), .Y(micro_hash_ucr_3_pipe45_bF_buf3) );
BUFX4 BUFX4_558 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe45), .Y(micro_hash_ucr_3_pipe45_bF_buf2) );
BUFX4 BUFX4_559 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe45), .Y(micro_hash_ucr_3_pipe45_bF_buf1) );
BUFX4 BUFX4_560 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe45), .Y(micro_hash_ucr_3_pipe45_bF_buf0) );
BUFX4 BUFX4_561 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe46), .Y(micro_hash_ucr_3_pipe46_bF_buf4) );
BUFX4 BUFX4_562 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe46), .Y(micro_hash_ucr_3_pipe46_bF_buf3) );
BUFX4 BUFX4_563 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe46), .Y(micro_hash_ucr_3_pipe46_bF_buf2) );
BUFX4 BUFX4_564 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe46), .Y(micro_hash_ucr_3_pipe46_bF_buf1) );
BUFX4 BUFX4_565 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe46), .Y(micro_hash_ucr_3_pipe46_bF_buf0) );
BUFX4 BUFX4_566 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe48), .Y(micro_hash_ucr_3_pipe48_bF_buf4) );
BUFX4 BUFX4_567 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe48), .Y(micro_hash_ucr_3_pipe48_bF_buf3) );
BUFX4 BUFX4_568 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe48), .Y(micro_hash_ucr_3_pipe48_bF_buf2) );
BUFX4 BUFX4_569 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe48), .Y(micro_hash_ucr_3_pipe48_bF_buf1) );
BUFX4 BUFX4_570 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe48), .Y(micro_hash_ucr_3_pipe48_bF_buf0) );
BUFX4 BUFX4_571 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe49), .Y(micro_hash_ucr_3_pipe49_bF_buf3) );
BUFX4 BUFX4_572 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe49), .Y(micro_hash_ucr_3_pipe49_bF_buf2) );
BUFX4 BUFX4_573 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe49), .Y(micro_hash_ucr_3_pipe49_bF_buf1) );
BUFX4 BUFX4_574 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe49), .Y(micro_hash_ucr_3_pipe49_bF_buf0) );
BUFX4 BUFX4_575 ( .gnd(gnd), .vdd(vdd), .A(_9325_), .Y(_9325__bF_buf3) );
BUFX4 BUFX4_576 ( .gnd(gnd), .vdd(vdd), .A(_9325_), .Y(_9325__bF_buf2) );
BUFX4 BUFX4_577 ( .gnd(gnd), .vdd(vdd), .A(_9325_), .Y(_9325__bF_buf1) );
BUFX4 BUFX4_578 ( .gnd(gnd), .vdd(vdd), .A(_9325_), .Y(_9325__bF_buf0) );
BUFX4 BUFX4_579 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_5_), .Y(micro_hash_ucr_3_b_5_bF_buf3_) );
BUFX4 BUFX4_580 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_5_), .Y(micro_hash_ucr_3_b_5_bF_buf2_) );
BUFX4 BUFX4_581 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_5_), .Y(micro_hash_ucr_3_b_5_bF_buf1_) );
BUFX4 BUFX4_582 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_5_), .Y(micro_hash_ucr_3_b_5_bF_buf0_) );
BUFX4 BUFX4_583 ( .gnd(gnd), .vdd(vdd), .A(_5092_), .Y(_5092__bF_buf4) );
BUFX4 BUFX4_584 ( .gnd(gnd), .vdd(vdd), .A(_5092_), .Y(_5092__bF_buf3) );
BUFX4 BUFX4_585 ( .gnd(gnd), .vdd(vdd), .A(_5092_), .Y(_5092__bF_buf2) );
BUFX4 BUFX4_586 ( .gnd(gnd), .vdd(vdd), .A(_5092_), .Y(_5092__bF_buf1) );
BUFX4 BUFX4_587 ( .gnd(gnd), .vdd(vdd), .A(_5092_), .Y(_5092__bF_buf0) );
BUFX4 BUFX4_588 ( .gnd(gnd), .vdd(vdd), .A(_7561_), .Y(_7561__bF_buf4) );
BUFX4 BUFX4_589 ( .gnd(gnd), .vdd(vdd), .A(_7561_), .Y(_7561__bF_buf3) );
BUFX4 BUFX4_590 ( .gnd(gnd), .vdd(vdd), .A(_7561_), .Y(_7561__bF_buf2) );
BUFX4 BUFX4_591 ( .gnd(gnd), .vdd(vdd), .A(_7561_), .Y(_7561__bF_buf1) );
BUFX4 BUFX4_592 ( .gnd(gnd), .vdd(vdd), .A(_7561_), .Y(_7561__bF_buf0) );
BUFX4 BUFX4_593 ( .gnd(gnd), .vdd(vdd), .A(_5089_), .Y(_5089__bF_buf3) );
BUFX4 BUFX4_594 ( .gnd(gnd), .vdd(vdd), .A(_5089_), .Y(_5089__bF_buf2) );
BUFX4 BUFX4_595 ( .gnd(gnd), .vdd(vdd), .A(_5089_), .Y(_5089__bF_buf1) );
BUFX4 BUFX4_596 ( .gnd(gnd), .vdd(vdd), .A(_5089_), .Y(_5089__bF_buf0) );
BUFX4 BUFX4_597 ( .gnd(gnd), .vdd(vdd), .A(_5110_), .Y(_5110__bF_buf3) );
BUFX4 BUFX4_598 ( .gnd(gnd), .vdd(vdd), .A(_5110_), .Y(_5110__bF_buf2) );
BUFX4 BUFX4_599 ( .gnd(gnd), .vdd(vdd), .A(_5110_), .Y(_5110__bF_buf1) );
BUFX4 BUFX4_600 ( .gnd(gnd), .vdd(vdd), .A(_5110_), .Y(_5110__bF_buf0) );
BUFX4 BUFX4_601 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_1_), .Y(micro_hash_ucr_2_b_1_bF_buf3_) );
BUFX4 BUFX4_602 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_1_), .Y(micro_hash_ucr_2_b_1_bF_buf2_) );
BUFX4 BUFX4_603 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_1_), .Y(micro_hash_ucr_2_b_1_bF_buf1_) );
BUFX4 BUFX4_604 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_1_), .Y(micro_hash_ucr_2_b_1_bF_buf0_) );
BUFX4 BUFX4_605 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe10), .Y(micro_hash_ucr_3_pipe10_bF_buf3) );
BUFX4 BUFX4_606 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe10), .Y(micro_hash_ucr_3_pipe10_bF_buf2) );
BUFX4 BUFX4_607 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe10), .Y(micro_hash_ucr_3_pipe10_bF_buf1) );
BUFX4 BUFX4_608 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe10), .Y(micro_hash_ucr_3_pipe10_bF_buf0) );
BUFX4 BUFX4_609 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe14), .Y(micro_hash_ucr_3_pipe14_bF_buf3) );
BUFX4 BUFX4_610 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe14), .Y(micro_hash_ucr_3_pipe14_bF_buf2) );
BUFX4 BUFX4_611 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe14), .Y(micro_hash_ucr_3_pipe14_bF_buf1) );
BUFX4 BUFX4_612 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe14), .Y(micro_hash_ucr_3_pipe14_bF_buf0) );
BUFX4 BUFX4_613 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe15), .Y(micro_hash_ucr_3_pipe15_bF_buf3) );
BUFX4 BUFX4_614 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe15), .Y(micro_hash_ucr_3_pipe15_bF_buf2) );
BUFX4 BUFX4_615 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe15), .Y(micro_hash_ucr_3_pipe15_bF_buf1) );
BUFX4 BUFX4_616 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe15), .Y(micro_hash_ucr_3_pipe15_bF_buf0) );
BUFX4 BUFX4_617 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe16), .Y(micro_hash_ucr_3_pipe16_bF_buf4) );
BUFX4 BUFX4_618 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe16), .Y(micro_hash_ucr_3_pipe16_bF_buf3) );
BUFX4 BUFX4_619 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe16), .Y(micro_hash_ucr_3_pipe16_bF_buf2) );
BUFX4 BUFX4_620 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe16), .Y(micro_hash_ucr_3_pipe16_bF_buf1) );
BUFX4 BUFX4_621 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe16), .Y(micro_hash_ucr_3_pipe16_bF_buf0) );
BUFX4 BUFX4_622 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe17), .Y(micro_hash_ucr_3_pipe17_bF_buf3) );
BUFX4 BUFX4_623 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe17), .Y(micro_hash_ucr_3_pipe17_bF_buf2) );
BUFX4 BUFX4_624 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe17), .Y(micro_hash_ucr_3_pipe17_bF_buf1) );
BUFX4 BUFX4_625 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe17), .Y(micro_hash_ucr_3_pipe17_bF_buf0) );
BUFX4 BUFX4_626 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe18), .Y(micro_hash_ucr_3_pipe18_bF_buf4) );
BUFX4 BUFX4_627 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe18), .Y(micro_hash_ucr_3_pipe18_bF_buf3) );
BUFX4 BUFX4_628 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe18), .Y(micro_hash_ucr_3_pipe18_bF_buf2) );
BUFX4 BUFX4_629 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe18), .Y(micro_hash_ucr_3_pipe18_bF_buf1) );
BUFX4 BUFX4_630 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe18), .Y(micro_hash_ucr_3_pipe18_bF_buf0) );
BUFX4 BUFX4_631 ( .gnd(gnd), .vdd(vdd), .A(_9322_), .Y(_9322__bF_buf3) );
BUFX4 BUFX4_632 ( .gnd(gnd), .vdd(vdd), .A(_9322_), .Y(_9322__bF_buf2) );
BUFX4 BUFX4_633 ( .gnd(gnd), .vdd(vdd), .A(_9322_), .Y(_9322__bF_buf1) );
BUFX4 BUFX4_634 ( .gnd(gnd), .vdd(vdd), .A(_9322_), .Y(_9322__bF_buf0) );
BUFX4 BUFX4_635 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_2_), .Y(micro_hash_ucr_3_b_2_bF_buf3_) );
BUFX4 BUFX4_636 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_2_), .Y(micro_hash_ucr_3_b_2_bF_buf2_) );
BUFX4 BUFX4_637 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_2_), .Y(micro_hash_ucr_3_b_2_bF_buf1_) );
BUFX4 BUFX4_638 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_2_), .Y(micro_hash_ucr_3_b_2_bF_buf0_) );
BUFX4 BUFX4_639 ( .gnd(gnd), .vdd(vdd), .A(_6294_), .Y(_6294__bF_buf4) );
BUFX4 BUFX4_640 ( .gnd(gnd), .vdd(vdd), .A(_6294_), .Y(_6294__bF_buf3) );
BUFX4 BUFX4_641 ( .gnd(gnd), .vdd(vdd), .A(_6294_), .Y(_6294__bF_buf2) );
BUFX4 BUFX4_642 ( .gnd(gnd), .vdd(vdd), .A(_6294_), .Y(_6294__bF_buf1) );
BUFX4 BUFX4_643 ( .gnd(gnd), .vdd(vdd), .A(_6294_), .Y(_6294__bF_buf0) );
BUFX4 BUFX4_644 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_5_), .Y(micro_hash_ucr_3_a_5_bF_buf3_) );
BUFX4 BUFX4_645 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_5_), .Y(micro_hash_ucr_3_a_5_bF_buf2_) );
BUFX4 BUFX4_646 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_5_), .Y(micro_hash_ucr_3_a_5_bF_buf1_) );
BUFX4 BUFX4_647 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_5_), .Y(micro_hash_ucr_3_a_5_bF_buf0_) );
BUFX4 BUFX4_648 ( .gnd(gnd), .vdd(vdd), .A(_10386_), .Y(_10386__bF_buf5) );
BUFX4 BUFX4_649 ( .gnd(gnd), .vdd(vdd), .A(_10386_), .Y(_10386__bF_buf4) );
BUFX4 BUFX4_650 ( .gnd(gnd), .vdd(vdd), .A(_10386_), .Y(_10386__bF_buf3) );
BUFX4 BUFX4_651 ( .gnd(gnd), .vdd(vdd), .A(_10386_), .Y(_10386__bF_buf2) );
BUFX4 BUFX4_652 ( .gnd(gnd), .vdd(vdd), .A(_10386_), .Y(_10386__bF_buf1) );
BUFX4 BUFX4_653 ( .gnd(gnd), .vdd(vdd), .A(_10386_), .Y(_10386__bF_buf0) );
BUFX4 BUFX4_654 ( .gnd(gnd), .vdd(vdd), .A(_5086_), .Y(_5086__bF_buf3) );
BUFX4 BUFX4_655 ( .gnd(gnd), .vdd(vdd), .A(_5086_), .Y(_5086__bF_buf2) );
BUFX4 BUFX4_656 ( .gnd(gnd), .vdd(vdd), .A(_5086_), .Y(_5086__bF_buf1) );
BUFX4 BUFX4_657 ( .gnd(gnd), .vdd(vdd), .A(_5086_), .Y(_5086__bF_buf0) );
BUFX4 BUFX4_658 ( .gnd(gnd), .vdd(vdd), .A(_414_), .Y(_414__bF_buf3) );
BUFX4 BUFX4_659 ( .gnd(gnd), .vdd(vdd), .A(_414_), .Y(_414__bF_buf2) );
BUFX4 BUFX4_660 ( .gnd(gnd), .vdd(vdd), .A(_414_), .Y(_414__bF_buf1) );
BUFX4 BUFX4_661 ( .gnd(gnd), .vdd(vdd), .A(_414_), .Y(_414__bF_buf0) );
BUFX4 BUFX4_662 ( .gnd(gnd), .vdd(vdd), .A(_9701_), .Y(_9701__bF_buf3) );
BUFX4 BUFX4_663 ( .gnd(gnd), .vdd(vdd), .A(_9701_), .Y(_9701__bF_buf2) );
BUFX4 BUFX4_664 ( .gnd(gnd), .vdd(vdd), .A(_9701_), .Y(_9701__bF_buf1) );
BUFX4 BUFX4_665 ( .gnd(gnd), .vdd(vdd), .A(_9701_), .Y(_9701__bF_buf0) );
BUFX4 BUFX4_666 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe70), .Y(micro_hash_ucr_pipe70_bF_buf3) );
BUFX4 BUFX4_667 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe70), .Y(micro_hash_ucr_pipe70_bF_buf2) );
BUFX4 BUFX4_668 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe70), .Y(micro_hash_ucr_pipe70_bF_buf1) );
BUFX4 BUFX4_669 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe70), .Y(micro_hash_ucr_pipe70_bF_buf0) );
BUFX4 BUFX4_670 ( .gnd(gnd), .vdd(vdd), .A(_9298_), .Y(_9298__bF_buf4) );
BUFX4 BUFX4_671 ( .gnd(gnd), .vdd(vdd), .A(_9298_), .Y(_9298__bF_buf3) );
BUFX4 BUFX4_672 ( .gnd(gnd), .vdd(vdd), .A(_9298_), .Y(_9298__bF_buf2) );
BUFX4 BUFX4_673 ( .gnd(gnd), .vdd(vdd), .A(_9298_), .Y(_9298__bF_buf1) );
BUFX4 BUFX4_674 ( .gnd(gnd), .vdd(vdd), .A(_9298_), .Y(_9298__bF_buf0) );
BUFX4 BUFX4_675 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_1_), .Y(micro_hash_ucr_2_a_1_bF_buf3_) );
BUFX4 BUFX4_676 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_1_), .Y(micro_hash_ucr_2_a_1_bF_buf2_) );
BUFX4 BUFX4_677 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_1_), .Y(micro_hash_ucr_2_a_1_bF_buf1_) );
BUFX4 BUFX4_678 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_1_), .Y(micro_hash_ucr_2_a_1_bF_buf0_) );
BUFX4 BUFX4_679 ( .gnd(gnd), .vdd(vdd), .A(_5104_), .Y(_5104__bF_buf4) );
BUFX4 BUFX4_680 ( .gnd(gnd), .vdd(vdd), .A(_5104_), .Y(_5104__bF_buf3) );
BUFX4 BUFX4_681 ( .gnd(gnd), .vdd(vdd), .A(_5104_), .Y(_5104__bF_buf2) );
BUFX4 BUFX4_682 ( .gnd(gnd), .vdd(vdd), .A(_5104_), .Y(_5104__bF_buf1) );
BUFX4 BUFX4_683 ( .gnd(gnd), .vdd(vdd), .A(_5104_), .Y(_5104__bF_buf0) );
BUFX4 BUFX4_684 ( .gnd(gnd), .vdd(vdd), .A(_10994_), .Y(_10994__bF_buf4) );
BUFX4 BUFX4_685 ( .gnd(gnd), .vdd(vdd), .A(_10994_), .Y(_10994__bF_buf3) );
BUFX4 BUFX4_686 ( .gnd(gnd), .vdd(vdd), .A(_10994_), .Y(_10994__bF_buf2) );
BUFX4 BUFX4_687 ( .gnd(gnd), .vdd(vdd), .A(_10994_), .Y(_10994__bF_buf1) );
BUFX4 BUFX4_688 ( .gnd(gnd), .vdd(vdd), .A(_10994_), .Y(_10994__bF_buf0) );
BUFX4 BUFX4_689 ( .gnd(gnd), .vdd(vdd), .A(_9316_), .Y(_9316__bF_buf3) );
BUFX4 BUFX4_690 ( .gnd(gnd), .vdd(vdd), .A(_9316_), .Y(_9316__bF_buf2) );
BUFX4 BUFX4_691 ( .gnd(gnd), .vdd(vdd), .A(_9316_), .Y(_9316__bF_buf1) );
BUFX4 BUFX4_692 ( .gnd(gnd), .vdd(vdd), .A(_9316_), .Y(_9316__bF_buf0) );
BUFX4 BUFX4_693 ( .gnd(gnd), .vdd(vdd), .A(_13217_), .Y(_13217__bF_buf4) );
BUFX4 BUFX4_694 ( .gnd(gnd), .vdd(vdd), .A(_13217_), .Y(_13217__bF_buf3) );
BUFX4 BUFX4_695 ( .gnd(gnd), .vdd(vdd), .A(_13217_), .Y(_13217__bF_buf2) );
BUFX4 BUFX4_696 ( .gnd(gnd), .vdd(vdd), .A(_13217_), .Y(_13217__bF_buf1) );
BUFX4 BUFX4_697 ( .gnd(gnd), .vdd(vdd), .A(_13217_), .Y(_13217__bF_buf0) );
BUFX4 BUFX4_698 ( .gnd(gnd), .vdd(vdd), .A(_5139_), .Y(_5139__bF_buf3) );
BUFX4 BUFX4_699 ( .gnd(gnd), .vdd(vdd), .A(_5139_), .Y(_5139__bF_buf2) );
BUFX4 BUFX4_700 ( .gnd(gnd), .vdd(vdd), .A(_5139_), .Y(_5139__bF_buf1) );
BUFX4 BUFX4_701 ( .gnd(gnd), .vdd(vdd), .A(_5139_), .Y(_5139__bF_buf0) );
BUFX4 BUFX4_702 ( .gnd(gnd), .vdd(vdd), .A(_12908_), .Y(_12908__bF_buf3) );
BUFX4 BUFX4_703 ( .gnd(gnd), .vdd(vdd), .A(_12908_), .Y(_12908__bF_buf2) );
BUFX4 BUFX4_704 ( .gnd(gnd), .vdd(vdd), .A(_12908_), .Y(_12908__bF_buf1) );
BUFX4 BUFX4_705 ( .gnd(gnd), .vdd(vdd), .A(_12908_), .Y(_12908__bF_buf0) );
BUFX4 BUFX4_706 ( .gnd(gnd), .vdd(vdd), .A(_13484_), .Y(_13484__bF_buf3) );
BUFX4 BUFX4_707 ( .gnd(gnd), .vdd(vdd), .A(_13484_), .Y(_13484__bF_buf2) );
BUFX4 BUFX4_708 ( .gnd(gnd), .vdd(vdd), .A(_13484_), .Y(_13484__bF_buf1) );
BUFX4 BUFX4_709 ( .gnd(gnd), .vdd(vdd), .A(_13484_), .Y(_13484__bF_buf0) );
BUFX4 BUFX4_710 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe40), .Y(micro_hash_ucr_pipe40_bF_buf4) );
BUFX4 BUFX4_711 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe40), .Y(micro_hash_ucr_pipe40_bF_buf3) );
BUFX4 BUFX4_712 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe40), .Y(micro_hash_ucr_pipe40_bF_buf2) );
BUFX4 BUFX4_713 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe40), .Y(micro_hash_ucr_pipe40_bF_buf1) );
BUFX4 BUFX4_714 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe40), .Y(micro_hash_ucr_pipe40_bF_buf0) );
BUFX4 BUFX4_715 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe42), .Y(micro_hash_ucr_pipe42_bF_buf3) );
BUFX4 BUFX4_716 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe42), .Y(micro_hash_ucr_pipe42_bF_buf2) );
BUFX4 BUFX4_717 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe42), .Y(micro_hash_ucr_pipe42_bF_buf1) );
BUFX4 BUFX4_718 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe42), .Y(micro_hash_ucr_pipe42_bF_buf0) );
BUFX4 BUFX4_719 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe45), .Y(micro_hash_ucr_pipe45_bF_buf3) );
BUFX4 BUFX4_720 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe45), .Y(micro_hash_ucr_pipe45_bF_buf2) );
BUFX4 BUFX4_721 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe45), .Y(micro_hash_ucr_pipe45_bF_buf1) );
BUFX4 BUFX4_722 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe45), .Y(micro_hash_ucr_pipe45_bF_buf0) );
BUFX4 BUFX4_723 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe46), .Y(micro_hash_ucr_pipe46_bF_buf4) );
BUFX4 BUFX4_724 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe46), .Y(micro_hash_ucr_pipe46_bF_buf3) );
BUFX4 BUFX4_725 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe46), .Y(micro_hash_ucr_pipe46_bF_buf2) );
BUFX4 BUFX4_726 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe46), .Y(micro_hash_ucr_pipe46_bF_buf1) );
BUFX4 BUFX4_727 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe46), .Y(micro_hash_ucr_pipe46_bF_buf0) );
BUFX4 BUFX4_728 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe48), .Y(micro_hash_ucr_pipe48_bF_buf3) );
BUFX4 BUFX4_729 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe48), .Y(micro_hash_ucr_pipe48_bF_buf2) );
BUFX4 BUFX4_730 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe48), .Y(micro_hash_ucr_pipe48_bF_buf1) );
BUFX4 BUFX4_731 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe48), .Y(micro_hash_ucr_pipe48_bF_buf0) );
BUFX4 BUFX4_732 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_2_), .Y(micro_hash_ucr_c_2_bF_buf3_) );
BUFX4 BUFX4_733 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_2_), .Y(micro_hash_ucr_c_2_bF_buf2_) );
BUFX4 BUFX4_734 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_2_), .Y(micro_hash_ucr_c_2_bF_buf1_) );
BUFX4 BUFX4_735 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_2_), .Y(micro_hash_ucr_c_2_bF_buf0_) );
BUFX4 BUFX4_736 ( .gnd(gnd), .vdd(vdd), .A(_925_), .Y(_925__bF_buf4) );
BUFX4 BUFX4_737 ( .gnd(gnd), .vdd(vdd), .A(_925_), .Y(_925__bF_buf3) );
BUFX4 BUFX4_738 ( .gnd(gnd), .vdd(vdd), .A(_925_), .Y(_925__bF_buf2) );
BUFX4 BUFX4_739 ( .gnd(gnd), .vdd(vdd), .A(_925_), .Y(_925__bF_buf1) );
BUFX4 BUFX4_740 ( .gnd(gnd), .vdd(vdd), .A(_925_), .Y(_925__bF_buf0) );
BUFX4 BUFX4_741 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_5_), .Y(micro_hash_ucr_b_5_bF_buf3_) );
BUFX4 BUFX4_742 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_5_), .Y(micro_hash_ucr_b_5_bF_buf2_) );
BUFX4 BUFX4_743 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_5_), .Y(micro_hash_ucr_b_5_bF_buf1_) );
BUFX4 BUFX4_744 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_5_), .Y(micro_hash_ucr_b_5_bF_buf0_) );
BUFX4 BUFX4_745 ( .gnd(gnd), .vdd(vdd), .A(comparador_2_valid), .Y(comparador_2_valid_bF_buf4) );
BUFX4 BUFX4_746 ( .gnd(gnd), .vdd(vdd), .A(comparador_2_valid), .Y(comparador_2_valid_bF_buf3) );
BUFX4 BUFX4_747 ( .gnd(gnd), .vdd(vdd), .A(comparador_2_valid), .Y(comparador_2_valid_bF_buf2) );
BUFX4 BUFX4_748 ( .gnd(gnd), .vdd(vdd), .A(comparador_2_valid), .Y(comparador_2_valid_bF_buf1) );
BUFX4 BUFX4_749 ( .gnd(gnd), .vdd(vdd), .A(comparador_2_valid), .Y(comparador_2_valid_bF_buf0) );
BUFX4 BUFX4_750 ( .gnd(gnd), .vdd(vdd), .A(_6153_), .Y(_6153__bF_buf5) );
BUFX4 BUFX4_751 ( .gnd(gnd), .vdd(vdd), .A(_6153_), .Y(_6153__bF_buf4) );
BUFX4 BUFX4_752 ( .gnd(gnd), .vdd(vdd), .A(_6153_), .Y(_6153__bF_buf3) );
BUFX4 BUFX4_753 ( .gnd(gnd), .vdd(vdd), .A(_6153_), .Y(_6153__bF_buf2) );
BUFX4 BUFX4_754 ( .gnd(gnd), .vdd(vdd), .A(_6153_), .Y(_6153__bF_buf1) );
BUFX4 BUFX4_755 ( .gnd(gnd), .vdd(vdd), .A(_6153_), .Y(_6153__bF_buf0) );
BUFX4 BUFX4_756 ( .gnd(gnd), .vdd(vdd), .A(_5080_), .Y(_5080__bF_buf3) );
BUFX4 BUFX4_757 ( .gnd(gnd), .vdd(vdd), .A(_5080_), .Y(_5080__bF_buf2) );
BUFX4 BUFX4_758 ( .gnd(gnd), .vdd(vdd), .A(_5080_), .Y(_5080__bF_buf1) );
BUFX4 BUFX4_759 ( .gnd(gnd), .vdd(vdd), .A(_5080_), .Y(_5080__bF_buf0) );
BUFX4 BUFX4_760 ( .gnd(gnd), .vdd(vdd), .A(_5365_), .Y(_5365__bF_buf3) );
BUFX4 BUFX4_761 ( .gnd(gnd), .vdd(vdd), .A(_5365_), .Y(_5365__bF_buf2) );
BUFX4 BUFX4_762 ( .gnd(gnd), .vdd(vdd), .A(_5365_), .Y(_5365__bF_buf1) );
BUFX4 BUFX4_763 ( .gnd(gnd), .vdd(vdd), .A(_5365_), .Y(_5365__bF_buf0) );
BUFX4 BUFX4_764 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe14), .Y(micro_hash_ucr_pipe14_bF_buf4) );
BUFX4 BUFX4_765 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe14), .Y(micro_hash_ucr_pipe14_bF_buf3) );
BUFX4 BUFX4_766 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe14), .Y(micro_hash_ucr_pipe14_bF_buf2) );
BUFX4 BUFX4_767 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe14), .Y(micro_hash_ucr_pipe14_bF_buf1) );
BUFX4 BUFX4_768 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe14), .Y(micro_hash_ucr_pipe14_bF_buf0) );
BUFX4 BUFX4_769 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe15), .Y(micro_hash_ucr_pipe15_bF_buf3) );
BUFX4 BUFX4_770 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe15), .Y(micro_hash_ucr_pipe15_bF_buf2) );
BUFX4 BUFX4_771 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe15), .Y(micro_hash_ucr_pipe15_bF_buf1) );
BUFX4 BUFX4_772 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe15), .Y(micro_hash_ucr_pipe15_bF_buf0) );
BUFX4 BUFX4_773 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe16), .Y(micro_hash_ucr_pipe16_bF_buf3) );
BUFX4 BUFX4_774 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe16), .Y(micro_hash_ucr_pipe16_bF_buf2) );
BUFX4 BUFX4_775 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe16), .Y(micro_hash_ucr_pipe16_bF_buf1) );
BUFX4 BUFX4_776 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe16), .Y(micro_hash_ucr_pipe16_bF_buf0) );
BUFX4 BUFX4_777 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe17), .Y(micro_hash_ucr_pipe17_bF_buf3) );
BUFX4 BUFX4_778 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe17), .Y(micro_hash_ucr_pipe17_bF_buf2) );
BUFX4 BUFX4_779 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe17), .Y(micro_hash_ucr_pipe17_bF_buf1) );
BUFX4 BUFX4_780 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe17), .Y(micro_hash_ucr_pipe17_bF_buf0) );
BUFX4 BUFX4_781 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe18), .Y(micro_hash_ucr_pipe18_bF_buf4) );
BUFX4 BUFX4_782 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe18), .Y(micro_hash_ucr_pipe18_bF_buf3) );
BUFX4 BUFX4_783 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe18), .Y(micro_hash_ucr_pipe18_bF_buf2) );
BUFX4 BUFX4_784 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe18), .Y(micro_hash_ucr_pipe18_bF_buf1) );
BUFX4 BUFX4_785 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe18), .Y(micro_hash_ucr_pipe18_bF_buf0) );
BUFX4 BUFX4_786 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe19), .Y(micro_hash_ucr_pipe19_bF_buf3) );
BUFX4 BUFX4_787 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe19), .Y(micro_hash_ucr_pipe19_bF_buf2) );
BUFX4 BUFX4_788 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe19), .Y(micro_hash_ucr_pipe19_bF_buf1) );
BUFX4 BUFX4_789 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe19), .Y(micro_hash_ucr_pipe19_bF_buf0) );
BUFX4 BUFX4_790 ( .gnd(gnd), .vdd(vdd), .A(_4674_), .Y(_4674__bF_buf3) );
BUFX4 BUFX4_791 ( .gnd(gnd), .vdd(vdd), .A(_4674_), .Y(_4674__bF_buf2) );
BUFX4 BUFX4_792 ( .gnd(gnd), .vdd(vdd), .A(_4674_), .Y(_4674__bF_buf1) );
BUFX4 BUFX4_793 ( .gnd(gnd), .vdd(vdd), .A(_4674_), .Y(_4674__bF_buf0) );
BUFX4 BUFX4_794 ( .gnd(gnd), .vdd(vdd), .A(_9292_), .Y(_9292__bF_buf3) );
BUFX4 BUFX4_795 ( .gnd(gnd), .vdd(vdd), .A(_9292_), .Y(_9292__bF_buf2) );
BUFX4 BUFX4_796 ( .gnd(gnd), .vdd(vdd), .A(_9292_), .Y(_9292__bF_buf1) );
BUFX4 BUFX4_797 ( .gnd(gnd), .vdd(vdd), .A(_9292_), .Y(_9292__bF_buf0) );
BUFX4 BUFX4_798 ( .gnd(gnd), .vdd(vdd), .A(_5077_), .Y(_5077__bF_buf3) );
BUFX4 BUFX4_799 ( .gnd(gnd), .vdd(vdd), .A(_5077_), .Y(_5077__bF_buf2) );
BUFX4 BUFX4_800 ( .gnd(gnd), .vdd(vdd), .A(_5077_), .Y(_5077__bF_buf1) );
BUFX4 BUFX4_801 ( .gnd(gnd), .vdd(vdd), .A(_5077_), .Y(_5077__bF_buf0) );
BUFX4 BUFX4_802 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_2_), .Y(micro_hash_ucr_b_2_bF_buf3_) );
BUFX4 BUFX4_803 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_2_), .Y(micro_hash_ucr_b_2_bF_buf2_) );
BUFX4 BUFX4_804 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_2_), .Y(micro_hash_ucr_b_2_bF_buf1_) );
BUFX4 BUFX4_805 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_2_), .Y(micro_hash_ucr_b_2_bF_buf0_) );
BUFX4 BUFX4_806 ( .gnd(gnd), .vdd(vdd), .A(_9289_), .Y(_9289__bF_buf3) );
BUFX4 BUFX4_807 ( .gnd(gnd), .vdd(vdd), .A(_9289_), .Y(_9289__bF_buf2) );
BUFX4 BUFX4_808 ( .gnd(gnd), .vdd(vdd), .A(_9289_), .Y(_9289__bF_buf1) );
BUFX4 BUFX4_809 ( .gnd(gnd), .vdd(vdd), .A(_9289_), .Y(_9289__bF_buf0) );
BUFX4 BUFX4_810 ( .gnd(gnd), .vdd(vdd), .A(_919_), .Y(_919__bF_buf4) );
BUFX4 BUFX4_811 ( .gnd(gnd), .vdd(vdd), .A(_919_), .Y(_919__bF_buf3) );
BUFX4 BUFX4_812 ( .gnd(gnd), .vdd(vdd), .A(_919_), .Y(_919__bF_buf2) );
BUFX4 BUFX4_813 ( .gnd(gnd), .vdd(vdd), .A(_919_), .Y(_919__bF_buf1) );
BUFX4 BUFX4_814 ( .gnd(gnd), .vdd(vdd), .A(_919_), .Y(_919__bF_buf0) );
BUFX4 BUFX4_815 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_5_), .Y(micro_hash_ucr_a_5_bF_buf3_) );
BUFX4 BUFX4_816 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_5_), .Y(micro_hash_ucr_a_5_bF_buf2_) );
BUFX4 BUFX4_817 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_5_), .Y(micro_hash_ucr_a_5_bF_buf1_) );
BUFX4 BUFX4_818 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_5_), .Y(micro_hash_ucr_a_5_bF_buf0_) );
BUFX4 BUFX4_819 ( .gnd(gnd), .vdd(vdd), .A(_8789_), .Y(_8789__bF_buf3) );
BUFX4 BUFX4_820 ( .gnd(gnd), .vdd(vdd), .A(_8789_), .Y(_8789__bF_buf2) );
BUFX4 BUFX4_821 ( .gnd(gnd), .vdd(vdd), .A(_8789_), .Y(_8789__bF_buf1) );
BUFX4 BUFX4_822 ( .gnd(gnd), .vdd(vdd), .A(_8789_), .Y(_8789__bF_buf0) );
BUFX4 BUFX4_823 ( .gnd(gnd), .vdd(vdd), .A(_9310_), .Y(_9310__bF_buf4) );
BUFX4 BUFX4_824 ( .gnd(gnd), .vdd(vdd), .A(_9310_), .Y(_9310__bF_buf3) );
BUFX4 BUFX4_825 ( .gnd(gnd), .vdd(vdd), .A(_9310_), .Y(_9310__bF_buf2) );
BUFX4 BUFX4_826 ( .gnd(gnd), .vdd(vdd), .A(_9310_), .Y(_9310__bF_buf1) );
BUFX4 BUFX4_827 ( .gnd(gnd), .vdd(vdd), .A(_9310_), .Y(_9310__bF_buf0) );
BUFX4 BUFX4_828 ( .gnd(gnd), .vdd(vdd), .A(_7067_), .Y(_7067__bF_buf5) );
BUFX4 BUFX4_829 ( .gnd(gnd), .vdd(vdd), .A(_7067_), .Y(_7067__bF_buf4) );
BUFX4 BUFX4_830 ( .gnd(gnd), .vdd(vdd), .A(_7067_), .Y(_7067__bF_buf3) );
BUFX4 BUFX4_831 ( .gnd(gnd), .vdd(vdd), .A(_7067_), .Y(_7067__bF_buf2) );
BUFX4 BUFX4_832 ( .gnd(gnd), .vdd(vdd), .A(_7067_), .Y(_7067__bF_buf1) );
BUFX4 BUFX4_833 ( .gnd(gnd), .vdd(vdd), .A(_7067_), .Y(_7067__bF_buf0) );
BUFX4 BUFX4_834 ( .gnd(gnd), .vdd(vdd), .A(_5074_), .Y(_5074__bF_buf3) );
BUFX4 BUFX4_835 ( .gnd(gnd), .vdd(vdd), .A(_5074_), .Y(_5074__bF_buf2) );
BUFX4 BUFX4_836 ( .gnd(gnd), .vdd(vdd), .A(_5074_), .Y(_5074__bF_buf1) );
BUFX4 BUFX4_837 ( .gnd(gnd), .vdd(vdd), .A(_5074_), .Y(_5074__bF_buf0) );
BUFX4 BUFX4_838 ( .gnd(gnd), .vdd(vdd), .A(_4668_), .Y(_4668__bF_buf3) );
BUFX4 BUFX4_839 ( .gnd(gnd), .vdd(vdd), .A(_4668_), .Y(_4668__bF_buf2) );
BUFX4 BUFX4_840 ( .gnd(gnd), .vdd(vdd), .A(_4668_), .Y(_4668__bF_buf1) );
BUFX4 BUFX4_841 ( .gnd(gnd), .vdd(vdd), .A(_4668_), .Y(_4668__bF_buf0) );
BUFX4 BUFX4_842 ( .gnd(gnd), .vdd(vdd), .A(_9286_), .Y(_9286__bF_buf3) );
BUFX4 BUFX4_843 ( .gnd(gnd), .vdd(vdd), .A(_9286_), .Y(_9286__bF_buf2) );
BUFX4 BUFX4_844 ( .gnd(gnd), .vdd(vdd), .A(_9286_), .Y(_9286__bF_buf1) );
BUFX4 BUFX4_845 ( .gnd(gnd), .vdd(vdd), .A(_9286_), .Y(_9286__bF_buf0) );
BUFX4 BUFX4_846 ( .gnd(gnd), .vdd(vdd), .A(_1717_), .Y(_1717__bF_buf3) );
BUFX4 BUFX4_847 ( .gnd(gnd), .vdd(vdd), .A(_1717_), .Y(_1717__bF_buf2) );
BUFX4 BUFX4_848 ( .gnd(gnd), .vdd(vdd), .A(_1717_), .Y(_1717__bF_buf1) );
BUFX4 BUFX4_849 ( .gnd(gnd), .vdd(vdd), .A(_1717_), .Y(_1717__bF_buf0) );
BUFX4 BUFX4_850 ( .gnd(gnd), .vdd(vdd), .A(_9304_), .Y(_9304__bF_buf3) );
BUFX4 BUFX4_851 ( .gnd(gnd), .vdd(vdd), .A(_9304_), .Y(_9304__bF_buf2) );
BUFX4 BUFX4_852 ( .gnd(gnd), .vdd(vdd), .A(_9304_), .Y(_9304__bF_buf1) );
BUFX4 BUFX4_853 ( .gnd(gnd), .vdd(vdd), .A(_9304_), .Y(_9304__bF_buf0) );
BUFX4 BUFX4_854 ( .gnd(gnd), .vdd(vdd), .A(_895_), .Y(_895__bF_buf4) );
BUFX4 BUFX4_855 ( .gnd(gnd), .vdd(vdd), .A(_895_), .Y(_895__bF_buf3) );
BUFX4 BUFX4_856 ( .gnd(gnd), .vdd(vdd), .A(_895_), .Y(_895__bF_buf2) );
BUFX4 BUFX4_857 ( .gnd(gnd), .vdd(vdd), .A(_895_), .Y(_895__bF_buf1) );
BUFX4 BUFX4_858 ( .gnd(gnd), .vdd(vdd), .A(_895_), .Y(_895__bF_buf0) );
BUFX4 BUFX4_859 ( .gnd(gnd), .vdd(vdd), .A(_0_), .Y(_0__bF_buf9) );
BUFX4 BUFX4_860 ( .gnd(gnd), .vdd(vdd), .A(_0_), .Y(_0__bF_buf8) );
BUFX4 BUFX4_861 ( .gnd(gnd), .vdd(vdd), .A(_0_), .Y(_0__bF_buf7) );
BUFX4 BUFX4_862 ( .gnd(gnd), .vdd(vdd), .A(_0_), .Y(_0__bF_buf6) );
BUFX4 BUFX4_863 ( .gnd(gnd), .vdd(vdd), .A(_0_), .Y(_0__bF_buf5) );
BUFX4 BUFX4_864 ( .gnd(gnd), .vdd(vdd), .A(_0_), .Y(_0__bF_buf4) );
BUFX4 BUFX4_865 ( .gnd(gnd), .vdd(vdd), .A(_0_), .Y(_0__bF_buf3) );
BUFX4 BUFX4_866 ( .gnd(gnd), .vdd(vdd), .A(_0_), .Y(_0__bF_buf2) );
BUFX4 BUFX4_867 ( .gnd(gnd), .vdd(vdd), .A(_0_), .Y(_0__bF_buf1) );
BUFX4 BUFX4_868 ( .gnd(gnd), .vdd(vdd), .A(_0_), .Y(_0__bF_buf0) );
BUFX4 BUFX4_869 ( .gnd(gnd), .vdd(vdd), .A(_5127_), .Y(_5127__bF_buf3) );
BUFX4 BUFX4_870 ( .gnd(gnd), .vdd(vdd), .A(_5127_), .Y(_5127__bF_buf2) );
BUFX4 BUFX4_871 ( .gnd(gnd), .vdd(vdd), .A(_5127_), .Y(_5127__bF_buf1) );
BUFX4 BUFX4_872 ( .gnd(gnd), .vdd(vdd), .A(_5127_), .Y(_5127__bF_buf0) );
BUFX4 BUFX4_873 ( .gnd(gnd), .vdd(vdd), .A(_7311_), .Y(_7311__bF_buf3) );
BUFX4 BUFX4_874 ( .gnd(gnd), .vdd(vdd), .A(_7311_), .Y(_7311__bF_buf2) );
BUFX4 BUFX4_875 ( .gnd(gnd), .vdd(vdd), .A(_7311_), .Y(_7311__bF_buf1) );
BUFX4 BUFX4_876 ( .gnd(gnd), .vdd(vdd), .A(_7311_), .Y(_7311__bF_buf0) );
BUFX4 BUFX4_877 ( .gnd(gnd), .vdd(vdd), .A(_9283_), .Y(_9283__bF_buf3) );
BUFX4 BUFX4_878 ( .gnd(gnd), .vdd(vdd), .A(_9283_), .Y(_9283__bF_buf2) );
BUFX4 BUFX4_879 ( .gnd(gnd), .vdd(vdd), .A(_9283_), .Y(_9283__bF_buf1) );
BUFX4 BUFX4_880 ( .gnd(gnd), .vdd(vdd), .A(_9283_), .Y(_9283__bF_buf0) );
BUFX4 BUFX4_881 ( .gnd(gnd), .vdd(vdd), .A(_913_), .Y(_913__bF_buf4) );
BUFX4 BUFX4_882 ( .gnd(gnd), .vdd(vdd), .A(_913_), .Y(_913__bF_buf3) );
BUFX4 BUFX4_883 ( .gnd(gnd), .vdd(vdd), .A(_913_), .Y(_913__bF_buf2) );
BUFX4 BUFX4_884 ( .gnd(gnd), .vdd(vdd), .A(_913_), .Y(_913__bF_buf1) );
BUFX4 BUFX4_885 ( .gnd(gnd), .vdd(vdd), .A(_913_), .Y(_913__bF_buf0) );
BUFX4 BUFX4_886 ( .gnd(gnd), .vdd(vdd), .A(_302_), .Y(_302__bF_buf13) );
BUFX4 BUFX4_887 ( .gnd(gnd), .vdd(vdd), .A(_302_), .Y(_302__bF_buf12) );
BUFX4 BUFX4_888 ( .gnd(gnd), .vdd(vdd), .A(_302_), .Y(_302__bF_buf11) );
BUFX4 BUFX4_889 ( .gnd(gnd), .vdd(vdd), .A(_302_), .Y(_302__bF_buf10) );
BUFX4 BUFX4_890 ( .gnd(gnd), .vdd(vdd), .A(_302_), .Y(_302__bF_buf9) );
BUFX4 BUFX4_891 ( .gnd(gnd), .vdd(vdd), .A(_302_), .Y(_302__bF_buf8) );
BUFX4 BUFX4_892 ( .gnd(gnd), .vdd(vdd), .A(_302_), .Y(_302__bF_buf7) );
BUFX4 BUFX4_893 ( .gnd(gnd), .vdd(vdd), .A(_302_), .Y(_302__bF_buf6) );
BUFX4 BUFX4_894 ( .gnd(gnd), .vdd(vdd), .A(_302_), .Y(_302__bF_buf5) );
BUFX4 BUFX4_895 ( .gnd(gnd), .vdd(vdd), .A(_302_), .Y(_302__bF_buf4) );
BUFX4 BUFX4_896 ( .gnd(gnd), .vdd(vdd), .A(_302_), .Y(_302__bF_buf3) );
BUFX4 BUFX4_897 ( .gnd(gnd), .vdd(vdd), .A(_302_), .Y(_302__bF_buf2) );
BUFX4 BUFX4_898 ( .gnd(gnd), .vdd(vdd), .A(_302_), .Y(_302__bF_buf1) );
BUFX4 BUFX4_899 ( .gnd(gnd), .vdd(vdd), .A(_302_), .Y(_302__bF_buf0) );
BUFX4 BUFX4_900 ( .gnd(gnd), .vdd(vdd), .A(_6808_), .Y(_6808__bF_buf4) );
BUFX4 BUFX4_901 ( .gnd(gnd), .vdd(vdd), .A(_6808_), .Y(_6808__bF_buf3) );
BUFX4 BUFX4_902 ( .gnd(gnd), .vdd(vdd), .A(_6808_), .Y(_6808__bF_buf2) );
BUFX4 BUFX4_903 ( .gnd(gnd), .vdd(vdd), .A(_6808_), .Y(_6808__bF_buf1) );
BUFX4 BUFX4_904 ( .gnd(gnd), .vdd(vdd), .A(_6808_), .Y(_6808__bF_buf0) );
BUFX4 BUFX4_905 ( .gnd(gnd), .vdd(vdd), .A(_9301_), .Y(_9301__bF_buf3) );
BUFX4 BUFX4_906 ( .gnd(gnd), .vdd(vdd), .A(_9301_), .Y(_9301__bF_buf2) );
BUFX4 BUFX4_907 ( .gnd(gnd), .vdd(vdd), .A(_9301_), .Y(_9301__bF_buf1) );
BUFX4 BUFX4_908 ( .gnd(gnd), .vdd(vdd), .A(_9301_), .Y(_9301__bF_buf0) );
BUFX4 BUFX4_909 ( .gnd(gnd), .vdd(vdd), .A(_5124_), .Y(_5124__bF_buf3) );
BUFX4 BUFX4_910 ( .gnd(gnd), .vdd(vdd), .A(_5124_), .Y(_5124__bF_buf2) );
BUFX4 BUFX4_911 ( .gnd(gnd), .vdd(vdd), .A(_5124_), .Y(_5124__bF_buf1) );
BUFX4 BUFX4_912 ( .gnd(gnd), .vdd(vdd), .A(_5124_), .Y(_5124__bF_buf0) );
BUFX4 BUFX4_913 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe70), .Y(micro_hash_ucr_2_pipe70_bF_buf3) );
BUFX4 BUFX4_914 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe70), .Y(micro_hash_ucr_2_pipe70_bF_buf2) );
BUFX4 BUFX4_915 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe70), .Y(micro_hash_ucr_2_pipe70_bF_buf1) );
BUFX4 BUFX4_916 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe70), .Y(micro_hash_ucr_2_pipe70_bF_buf0) );
BUFX4 BUFX4_917 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe6), .Y(micro_hash_ucr_3_pipe6_bF_buf3) );
BUFX4 BUFX4_918 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe6), .Y(micro_hash_ucr_3_pipe6_bF_buf2) );
BUFX4 BUFX4_919 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe6), .Y(micro_hash_ucr_3_pipe6_bF_buf1) );
BUFX4 BUFX4_920 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe6), .Y(micro_hash_ucr_3_pipe6_bF_buf0) );
BUFX4 BUFX4_921 ( .gnd(gnd), .vdd(vdd), .A(_889_), .Y(_889__bF_buf4) );
BUFX4 BUFX4_922 ( .gnd(gnd), .vdd(vdd), .A(_889_), .Y(_889__bF_buf3) );
BUFX4 BUFX4_923 ( .gnd(gnd), .vdd(vdd), .A(_889_), .Y(_889__bF_buf2) );
BUFX4 BUFX4_924 ( .gnd(gnd), .vdd(vdd), .A(_889_), .Y(_889__bF_buf1) );
BUFX4 BUFX4_925 ( .gnd(gnd), .vdd(vdd), .A(_889_), .Y(_889__bF_buf0) );
BUFX4 BUFX4_926 ( .gnd(gnd), .vdd(vdd), .A(_9336_), .Y(_9336__bF_buf3) );
BUFX4 BUFX4_927 ( .gnd(gnd), .vdd(vdd), .A(_9336_), .Y(_9336__bF_buf2) );
BUFX4 BUFX4_928 ( .gnd(gnd), .vdd(vdd), .A(_9336_), .Y(_9336__bF_buf1) );
BUFX4 BUFX4_929 ( .gnd(gnd), .vdd(vdd), .A(_9336_), .Y(_9336__bF_buf0) );
BUFX4 BUFX4_930 ( .gnd(gnd), .vdd(vdd), .A(_2305_), .Y(_2305__bF_buf3) );
BUFX4 BUFX4_931 ( .gnd(gnd), .vdd(vdd), .A(_2305_), .Y(_2305__bF_buf2) );
BUFX4 BUFX4_932 ( .gnd(gnd), .vdd(vdd), .A(_2305_), .Y(_2305__bF_buf1) );
BUFX4 BUFX4_933 ( .gnd(gnd), .vdd(vdd), .A(_2305_), .Y(_2305__bF_buf0) );
BUFX4 BUFX4_934 ( .gnd(gnd), .vdd(vdd), .A(_907_), .Y(_907__bF_buf4) );
BUFX4 BUFX4_935 ( .gnd(gnd), .vdd(vdd), .A(_907_), .Y(_907__bF_buf3) );
BUFX4 BUFX4_936 ( .gnd(gnd), .vdd(vdd), .A(_907_), .Y(_907__bF_buf2) );
BUFX4 BUFX4_937 ( .gnd(gnd), .vdd(vdd), .A(_907_), .Y(_907__bF_buf1) );
BUFX4 BUFX4_938 ( .gnd(gnd), .vdd(vdd), .A(_907_), .Y(_907__bF_buf0) );
BUFX4 BUFX4_939 ( .gnd(gnd), .vdd(vdd), .A(_6517_), .Y(_6517__bF_buf5) );
BUFX4 BUFX4_940 ( .gnd(gnd), .vdd(vdd), .A(_6517_), .Y(_6517__bF_buf4) );
BUFX4 BUFX4_941 ( .gnd(gnd), .vdd(vdd), .A(_6517_), .Y(_6517__bF_buf3) );
BUFX4 BUFX4_942 ( .gnd(gnd), .vdd(vdd), .A(_6517_), .Y(_6517__bF_buf2) );
BUFX4 BUFX4_943 ( .gnd(gnd), .vdd(vdd), .A(_6517_), .Y(_6517__bF_buf1) );
BUFX4 BUFX4_944 ( .gnd(gnd), .vdd(vdd), .A(_6517_), .Y(_6517__bF_buf0) );
BUFX4 BUFX4_945 ( .gnd(gnd), .vdd(vdd), .A(_2857_), .Y(_2857__bF_buf5) );
BUFX4 BUFX4_946 ( .gnd(gnd), .vdd(vdd), .A(_2857_), .Y(_2857__bF_buf4) );
BUFX4 BUFX4_947 ( .gnd(gnd), .vdd(vdd), .A(_2857_), .Y(_2857__bF_buf3) );
BUFX4 BUFX4_948 ( .gnd(gnd), .vdd(vdd), .A(_2857_), .Y(_2857__bF_buf2) );
BUFX4 BUFX4_949 ( .gnd(gnd), .vdd(vdd), .A(_2857_), .Y(_2857__bF_buf1) );
BUFX4 BUFX4_950 ( .gnd(gnd), .vdd(vdd), .A(_2857_), .Y(_2857__bF_buf0) );
BUFX4 BUFX4_951 ( .gnd(gnd), .vdd(vdd), .A(_5121_), .Y(_5121__bF_buf4) );
BUFX4 BUFX4_952 ( .gnd(gnd), .vdd(vdd), .A(_5121_), .Y(_5121__bF_buf3) );
BUFX4 BUFX4_953 ( .gnd(gnd), .vdd(vdd), .A(_5121_), .Y(_5121__bF_buf2) );
BUFX4 BUFX4_954 ( .gnd(gnd), .vdd(vdd), .A(_5121_), .Y(_5121__bF_buf1) );
BUFX4 BUFX4_955 ( .gnd(gnd), .vdd(vdd), .A(_5121_), .Y(_5121__bF_buf0) );
BUFX4 BUFX4_956 ( .gnd(gnd), .vdd(vdd), .A(_428_), .Y(_428__bF_buf3) );
BUFX4 BUFX4_957 ( .gnd(gnd), .vdd(vdd), .A(_428_), .Y(_428__bF_buf2) );
BUFX4 BUFX4_958 ( .gnd(gnd), .vdd(vdd), .A(_428_), .Y(_428__bF_buf1) );
BUFX4 BUFX4_959 ( .gnd(gnd), .vdd(vdd), .A(_428_), .Y(_428__bF_buf0) );
BUFX4 BUFX4_960 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe40), .Y(micro_hash_ucr_2_pipe40_bF_buf4) );
BUFX4 BUFX4_961 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe40), .Y(micro_hash_ucr_2_pipe40_bF_buf3) );
BUFX4 BUFX4_962 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe40), .Y(micro_hash_ucr_2_pipe40_bF_buf2) );
BUFX4 BUFX4_963 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe40), .Y(micro_hash_ucr_2_pipe40_bF_buf1) );
BUFX4 BUFX4_964 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe40), .Y(micro_hash_ucr_2_pipe40_bF_buf0) );
BUFX4 BUFX4_965 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe41), .Y(micro_hash_ucr_2_pipe41_bF_buf3) );
BUFX4 BUFX4_966 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe41), .Y(micro_hash_ucr_2_pipe41_bF_buf2) );
BUFX4 BUFX4_967 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe41), .Y(micro_hash_ucr_2_pipe41_bF_buf1) );
BUFX4 BUFX4_968 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe41), .Y(micro_hash_ucr_2_pipe41_bF_buf0) );
BUFX4 BUFX4_969 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe42), .Y(micro_hash_ucr_2_pipe42_bF_buf3) );
BUFX4 BUFX4_970 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe42), .Y(micro_hash_ucr_2_pipe42_bF_buf2) );
BUFX4 BUFX4_971 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe42), .Y(micro_hash_ucr_2_pipe42_bF_buf1) );
BUFX4 BUFX4_972 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe42), .Y(micro_hash_ucr_2_pipe42_bF_buf0) );
BUFX4 BUFX4_973 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe44), .Y(micro_hash_ucr_2_pipe44_bF_buf3) );
BUFX4 BUFX4_974 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe44), .Y(micro_hash_ucr_2_pipe44_bF_buf2) );
BUFX4 BUFX4_975 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe44), .Y(micro_hash_ucr_2_pipe44_bF_buf1) );
BUFX4 BUFX4_976 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe44), .Y(micro_hash_ucr_2_pipe44_bF_buf0) );
BUFX4 BUFX4_977 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe45), .Y(micro_hash_ucr_2_pipe45_bF_buf3) );
BUFX4 BUFX4_978 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe45), .Y(micro_hash_ucr_2_pipe45_bF_buf2) );
BUFX4 BUFX4_979 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe45), .Y(micro_hash_ucr_2_pipe45_bF_buf1) );
BUFX4 BUFX4_980 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe45), .Y(micro_hash_ucr_2_pipe45_bF_buf0) );
BUFX4 BUFX4_981 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe46), .Y(micro_hash_ucr_2_pipe46_bF_buf4) );
BUFX4 BUFX4_982 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe46), .Y(micro_hash_ucr_2_pipe46_bF_buf3) );
BUFX4 BUFX4_983 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe46), .Y(micro_hash_ucr_2_pipe46_bF_buf2) );
BUFX4 BUFX4_984 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe46), .Y(micro_hash_ucr_2_pipe46_bF_buf1) );
BUFX4 BUFX4_985 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe46), .Y(micro_hash_ucr_2_pipe46_bF_buf0) );
BUFX4 BUFX4_986 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe48), .Y(micro_hash_ucr_2_pipe48_bF_buf4) );
BUFX4 BUFX4_987 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe48), .Y(micro_hash_ucr_2_pipe48_bF_buf3) );
BUFX4 BUFX4_988 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe48), .Y(micro_hash_ucr_2_pipe48_bF_buf2) );
BUFX4 BUFX4_989 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe48), .Y(micro_hash_ucr_2_pipe48_bF_buf1) );
BUFX4 BUFX4_990 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe48), .Y(micro_hash_ucr_2_pipe48_bF_buf0) );
BUFX4 BUFX4_991 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe49), .Y(micro_hash_ucr_2_pipe49_bF_buf3) );
BUFX4 BUFX4_992 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe49), .Y(micro_hash_ucr_2_pipe49_bF_buf2) );
BUFX4 BUFX4_993 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe49), .Y(micro_hash_ucr_2_pipe49_bF_buf1) );
BUFX4 BUFX4_994 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe49), .Y(micro_hash_ucr_2_pipe49_bF_buf0) );
BUFX4 BUFX4_995 ( .gnd(gnd), .vdd(vdd), .A(_6135_), .Y(_6135__bF_buf3) );
BUFX4 BUFX4_996 ( .gnd(gnd), .vdd(vdd), .A(_6135_), .Y(_6135__bF_buf2) );
BUFX4 BUFX4_997 ( .gnd(gnd), .vdd(vdd), .A(_6135_), .Y(_6135__bF_buf1) );
BUFX4 BUFX4_998 ( .gnd(gnd), .vdd(vdd), .A(_6135_), .Y(_6135__bF_buf0) );
BUFX4 BUFX4_999 ( .gnd(gnd), .vdd(vdd), .A(_6784_), .Y(_6784__bF_buf4) );
BUFX4 BUFX4_1000 ( .gnd(gnd), .vdd(vdd), .A(_6784_), .Y(_6784__bF_buf3) );
BUFX4 BUFX4_1001 ( .gnd(gnd), .vdd(vdd), .A(_6784_), .Y(_6784__bF_buf2) );
BUFX4 BUFX4_1002 ( .gnd(gnd), .vdd(vdd), .A(_6784_), .Y(_6784__bF_buf1) );
BUFX4 BUFX4_1003 ( .gnd(gnd), .vdd(vdd), .A(_6784_), .Y(_6784__bF_buf0) );
BUFX4 BUFX4_1004 ( .gnd(gnd), .vdd(vdd), .A(target[7]), .Y(target_7_bF_buf3_) );
BUFX4 BUFX4_1005 ( .gnd(gnd), .vdd(vdd), .A(target[7]), .Y(target_7_bF_buf2_) );
BUFX4 BUFX4_1006 ( .gnd(gnd), .vdd(vdd), .A(target[7]), .Y(target_7_bF_buf1_) );
BUFX4 BUFX4_1007 ( .gnd(gnd), .vdd(vdd), .A(target[7]), .Y(target_7_bF_buf0_) );
BUFX4 BUFX4_1008 ( .gnd(gnd), .vdd(vdd), .A(_2569_), .Y(_2569__bF_buf4) );
BUFX4 BUFX4_1009 ( .gnd(gnd), .vdd(vdd), .A(_2569_), .Y(_2569__bF_buf3) );
BUFX4 BUFX4_1010 ( .gnd(gnd), .vdd(vdd), .A(_2569_), .Y(_2569__bF_buf2) );
BUFX4 BUFX4_1011 ( .gnd(gnd), .vdd(vdd), .A(_2569_), .Y(_2569__bF_buf1) );
BUFX4 BUFX4_1012 ( .gnd(gnd), .vdd(vdd), .A(_2569_), .Y(_2569__bF_buf0) );
BUFX4 BUFX4_1013 ( .gnd(gnd), .vdd(vdd), .A(_9333_), .Y(_9333__bF_buf3) );
BUFX4 BUFX4_1014 ( .gnd(gnd), .vdd(vdd), .A(_9333_), .Y(_9333__bF_buf2) );
BUFX4 BUFX4_1015 ( .gnd(gnd), .vdd(vdd), .A(_9333_), .Y(_9333__bF_buf1) );
BUFX4 BUFX4_1016 ( .gnd(gnd), .vdd(vdd), .A(_9333_), .Y(_9333__bF_buf0) );
BUFX4 BUFX4_1017 ( .gnd(gnd), .vdd(vdd), .A(_5118_), .Y(_5118__bF_buf3) );
BUFX4 BUFX4_1018 ( .gnd(gnd), .vdd(vdd), .A(_5118_), .Y(_5118__bF_buf2) );
BUFX4 BUFX4_1019 ( .gnd(gnd), .vdd(vdd), .A(_5118_), .Y(_5118__bF_buf1) );
BUFX4 BUFX4_1020 ( .gnd(gnd), .vdd(vdd), .A(_5118_), .Y(_5118__bF_buf0) );
BUFX4 BUFX4_1021 ( .gnd(gnd), .vdd(vdd), .A(_904_), .Y(_904__bF_buf3) );
BUFX4 BUFX4_1022 ( .gnd(gnd), .vdd(vdd), .A(_904_), .Y(_904__bF_buf2) );
BUFX4 BUFX4_1023 ( .gnd(gnd), .vdd(vdd), .A(_904_), .Y(_904__bF_buf1) );
BUFX4 BUFX4_1024 ( .gnd(gnd), .vdd(vdd), .A(_904_), .Y(_904__bF_buf0) );
BUFX4 BUFX4_1025 ( .gnd(gnd), .vdd(vdd), .A(_11852_), .Y(_11852__bF_buf3) );
BUFX4 BUFX4_1026 ( .gnd(gnd), .vdd(vdd), .A(_11852_), .Y(_11852__bF_buf2) );
BUFX4 BUFX4_1027 ( .gnd(gnd), .vdd(vdd), .A(_11852_), .Y(_11852__bF_buf1) );
BUFX4 BUFX4_1028 ( .gnd(gnd), .vdd(vdd), .A(_11852_), .Y(_11852__bF_buf0) );
BUFX4 BUFX4_1029 ( .gnd(gnd), .vdd(vdd), .A(_5097_), .Y(_5097__bF_buf3) );
BUFX4 BUFX4_1030 ( .gnd(gnd), .vdd(vdd), .A(_5097_), .Y(_5097__bF_buf2) );
BUFX4 BUFX4_1031 ( .gnd(gnd), .vdd(vdd), .A(_5097_), .Y(_5097__bF_buf1) );
BUFX4 BUFX4_1032 ( .gnd(gnd), .vdd(vdd), .A(_5097_), .Y(_5097__bF_buf0) );
BUFX4 BUFX4_1033 ( .gnd(gnd), .vdd(vdd), .A(_8868_), .Y(_8868__bF_buf3) );
BUFX4 BUFX4_1034 ( .gnd(gnd), .vdd(vdd), .A(_8868_), .Y(_8868__bF_buf2) );
BUFX4 BUFX4_1035 ( .gnd(gnd), .vdd(vdd), .A(_8868_), .Y(_8868__bF_buf1) );
BUFX4 BUFX4_1036 ( .gnd(gnd), .vdd(vdd), .A(_8868_), .Y(_8868__bF_buf0) );
BUFX4 BUFX4_1037 ( .gnd(gnd), .vdd(vdd), .A(_6514_), .Y(_6514__bF_buf3) );
BUFX4 BUFX4_1038 ( .gnd(gnd), .vdd(vdd), .A(_6514_), .Y(_6514__bF_buf2) );
BUFX4 BUFX4_1039 ( .gnd(gnd), .vdd(vdd), .A(_6514_), .Y(_6514__bF_buf1) );
BUFX4 BUFX4_1040 ( .gnd(gnd), .vdd(vdd), .A(_6514_), .Y(_6514__bF_buf0) );
BUFX4 BUFX4_1041 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe12), .Y(micro_hash_ucr_2_pipe12_bF_buf3) );
BUFX4 BUFX4_1042 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe12), .Y(micro_hash_ucr_2_pipe12_bF_buf2) );
BUFX4 BUFX4_1043 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe12), .Y(micro_hash_ucr_2_pipe12_bF_buf1) );
BUFX4 BUFX4_1044 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe12), .Y(micro_hash_ucr_2_pipe12_bF_buf0) );
BUFX4 BUFX4_1045 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe14), .Y(micro_hash_ucr_2_pipe14_bF_buf4) );
BUFX4 BUFX4_1046 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe14), .Y(micro_hash_ucr_2_pipe14_bF_buf3) );
BUFX4 BUFX4_1047 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe14), .Y(micro_hash_ucr_2_pipe14_bF_buf2) );
BUFX4 BUFX4_1048 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe14), .Y(micro_hash_ucr_2_pipe14_bF_buf1) );
BUFX4 BUFX4_1049 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe14), .Y(micro_hash_ucr_2_pipe14_bF_buf0) );
BUFX4 BUFX4_1050 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe16), .Y(micro_hash_ucr_2_pipe16_bF_buf4) );
BUFX4 BUFX4_1051 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe16), .Y(micro_hash_ucr_2_pipe16_bF_buf3) );
BUFX4 BUFX4_1052 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe16), .Y(micro_hash_ucr_2_pipe16_bF_buf2) );
BUFX4 BUFX4_1053 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe16), .Y(micro_hash_ucr_2_pipe16_bF_buf1) );
BUFX4 BUFX4_1054 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe16), .Y(micro_hash_ucr_2_pipe16_bF_buf0) );
BUFX4 BUFX4_1055 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe17), .Y(micro_hash_ucr_2_pipe17_bF_buf3) );
BUFX4 BUFX4_1056 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe17), .Y(micro_hash_ucr_2_pipe17_bF_buf2) );
BUFX4 BUFX4_1057 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe17), .Y(micro_hash_ucr_2_pipe17_bF_buf1) );
BUFX4 BUFX4_1058 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe17), .Y(micro_hash_ucr_2_pipe17_bF_buf0) );
BUFX4 BUFX4_1059 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe18), .Y(micro_hash_ucr_2_pipe18_bF_buf4) );
BUFX4 BUFX4_1060 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe18), .Y(micro_hash_ucr_2_pipe18_bF_buf3) );
BUFX4 BUFX4_1061 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe18), .Y(micro_hash_ucr_2_pipe18_bF_buf2) );
BUFX4 BUFX4_1062 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe18), .Y(micro_hash_ucr_2_pipe18_bF_buf1) );
BUFX4 BUFX4_1063 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe18), .Y(micro_hash_ucr_2_pipe18_bF_buf0) );
BUFX4 BUFX4_1064 ( .gnd(gnd), .vdd(vdd), .A(_883_), .Y(_883__bF_buf3) );
BUFX4 BUFX4_1065 ( .gnd(gnd), .vdd(vdd), .A(_883_), .Y(_883__bF_buf2) );
BUFX4 BUFX4_1066 ( .gnd(gnd), .vdd(vdd), .A(_883_), .Y(_883__bF_buf1) );
BUFX4 BUFX4_1067 ( .gnd(gnd), .vdd(vdd), .A(_883_), .Y(_883__bF_buf0) );
BUFX4 BUFX4_1068 ( .gnd(gnd), .vdd(vdd), .A(_2090_), .Y(_2090__bF_buf4) );
BUFX4 BUFX4_1069 ( .gnd(gnd), .vdd(vdd), .A(_2090_), .Y(_2090__bF_buf3) );
BUFX4 BUFX4_1070 ( .gnd(gnd), .vdd(vdd), .A(_2090_), .Y(_2090__bF_buf2) );
BUFX4 BUFX4_1071 ( .gnd(gnd), .vdd(vdd), .A(_2090_), .Y(_2090__bF_buf1) );
BUFX4 BUFX4_1072 ( .gnd(gnd), .vdd(vdd), .A(_2090_), .Y(_2090__bF_buf0) );
BUFX4 BUFX4_1073 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_3_), .Y(micro_hash_ucr_2_c_3_bF_buf3_) );
BUFX4 BUFX4_1074 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_3_), .Y(micro_hash_ucr_2_c_3_bF_buf2_) );
BUFX4 BUFX4_1075 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_3_), .Y(micro_hash_ucr_2_c_3_bF_buf1_) );
BUFX4 BUFX4_1076 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_3_), .Y(micro_hash_ucr_2_c_3_bF_buf0_) );
BUFX4 BUFX4_1077 ( .gnd(gnd), .vdd(vdd), .A(_9330_), .Y(_9330__bF_buf4) );
BUFX4 BUFX4_1078 ( .gnd(gnd), .vdd(vdd), .A(_9330_), .Y(_9330__bF_buf3) );
BUFX4 BUFX4_1079 ( .gnd(gnd), .vdd(vdd), .A(_9330_), .Y(_9330__bF_buf2) );
BUFX4 BUFX4_1080 ( .gnd(gnd), .vdd(vdd), .A(_9330_), .Y(_9330__bF_buf1) );
BUFX4 BUFX4_1081 ( .gnd(gnd), .vdd(vdd), .A(_9330_), .Y(_9330__bF_buf0) );
BUFX4 BUFX4_1082 ( .gnd(gnd), .vdd(vdd), .A(_5115_), .Y(_5115__bF_buf4) );
BUFX4 BUFX4_1083 ( .gnd(gnd), .vdd(vdd), .A(_5115_), .Y(_5115__bF_buf3) );
BUFX4 BUFX4_1084 ( .gnd(gnd), .vdd(vdd), .A(_5115_), .Y(_5115__bF_buf2) );
BUFX4 BUFX4_1085 ( .gnd(gnd), .vdd(vdd), .A(_5115_), .Y(_5115__bF_buf1) );
BUFX4 BUFX4_1086 ( .gnd(gnd), .vdd(vdd), .A(_5115_), .Y(_5115__bF_buf0) );
BUFX4 BUFX4_1087 ( .gnd(gnd), .vdd(vdd), .A(_10738_), .Y(_10738__bF_buf3) );
BUFX4 BUFX4_1088 ( .gnd(gnd), .vdd(vdd), .A(_10738_), .Y(_10738__bF_buf2) );
BUFX4 BUFX4_1089 ( .gnd(gnd), .vdd(vdd), .A(_10738_), .Y(_10738__bF_buf1) );
BUFX4 BUFX4_1090 ( .gnd(gnd), .vdd(vdd), .A(_10738_), .Y(_10738__bF_buf0) );
BUFX4 BUFX4_1091 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe60), .Y(micro_hash_ucr_3_pipe60_bF_buf4) );
BUFX4 BUFX4_1092 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe60), .Y(micro_hash_ucr_3_pipe60_bF_buf3) );
BUFX4 BUFX4_1093 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe60), .Y(micro_hash_ucr_3_pipe60_bF_buf2) );
BUFX4 BUFX4_1094 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe60), .Y(micro_hash_ucr_3_pipe60_bF_buf1) );
BUFX4 BUFX4_1095 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe60), .Y(micro_hash_ucr_3_pipe60_bF_buf0) );
BUFX4 BUFX4_1096 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe61), .Y(micro_hash_ucr_3_pipe61_bF_buf3) );
BUFX4 BUFX4_1097 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe61), .Y(micro_hash_ucr_3_pipe61_bF_buf2) );
BUFX4 BUFX4_1098 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe61), .Y(micro_hash_ucr_3_pipe61_bF_buf1) );
BUFX4 BUFX4_1099 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe61), .Y(micro_hash_ucr_3_pipe61_bF_buf0) );
BUFX4 BUFX4_1100 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe62), .Y(micro_hash_ucr_3_pipe62_bF_buf3) );
BUFX4 BUFX4_1101 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe62), .Y(micro_hash_ucr_3_pipe62_bF_buf2) );
BUFX4 BUFX4_1102 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe62), .Y(micro_hash_ucr_3_pipe62_bF_buf1) );
BUFX4 BUFX4_1103 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe62), .Y(micro_hash_ucr_3_pipe62_bF_buf0) );
BUFX4 BUFX4_1104 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe64), .Y(micro_hash_ucr_3_pipe64_bF_buf4) );
BUFX4 BUFX4_1105 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe64), .Y(micro_hash_ucr_3_pipe64_bF_buf3) );
BUFX4 BUFX4_1106 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe64), .Y(micro_hash_ucr_3_pipe64_bF_buf2) );
BUFX4 BUFX4_1107 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe64), .Y(micro_hash_ucr_3_pipe64_bF_buf1) );
BUFX4 BUFX4_1108 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe64), .Y(micro_hash_ucr_3_pipe64_bF_buf0) );
BUFX4 BUFX4_1109 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe65), .Y(micro_hash_ucr_3_pipe65_bF_buf3) );
BUFX4 BUFX4_1110 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe65), .Y(micro_hash_ucr_3_pipe65_bF_buf2) );
BUFX4 BUFX4_1111 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe65), .Y(micro_hash_ucr_3_pipe65_bF_buf1) );
BUFX4 BUFX4_1112 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe65), .Y(micro_hash_ucr_3_pipe65_bF_buf0) );
BUFX4 BUFX4_1113 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe66), .Y(micro_hash_ucr_3_pipe66_bF_buf4) );
BUFX4 BUFX4_1114 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe66), .Y(micro_hash_ucr_3_pipe66_bF_buf3) );
BUFX4 BUFX4_1115 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe66), .Y(micro_hash_ucr_3_pipe66_bF_buf2) );
BUFX4 BUFX4_1116 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe66), .Y(micro_hash_ucr_3_pipe66_bF_buf1) );
BUFX4 BUFX4_1117 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe66), .Y(micro_hash_ucr_3_pipe66_bF_buf0) );
BUFX4 BUFX4_1118 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe68), .Y(micro_hash_ucr_3_pipe68_bF_buf3) );
BUFX4 BUFX4_1119 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe68), .Y(micro_hash_ucr_3_pipe68_bF_buf2) );
BUFX4 BUFX4_1120 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe68), .Y(micro_hash_ucr_3_pipe68_bF_buf1) );
BUFX4 BUFX4_1121 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe68), .Y(micro_hash_ucr_3_pipe68_bF_buf0) );
BUFX4 BUFX4_1122 ( .gnd(gnd), .vdd(vdd), .A(_901_), .Y(_901__bF_buf4) );
BUFX4 BUFX4_1123 ( .gnd(gnd), .vdd(vdd), .A(_901_), .Y(_901__bF_buf3) );
BUFX4 BUFX4_1124 ( .gnd(gnd), .vdd(vdd), .A(_901_), .Y(_901__bF_buf2) );
BUFX4 BUFX4_1125 ( .gnd(gnd), .vdd(vdd), .A(_901_), .Y(_901__bF_buf1) );
BUFX4 BUFX4_1126 ( .gnd(gnd), .vdd(vdd), .A(_901_), .Y(_901__bF_buf0) );
BUFX4 BUFX4_1127 ( .gnd(gnd), .vdd(vdd), .A(_1167_), .Y(_1167__bF_buf3) );
BUFX4 BUFX4_1128 ( .gnd(gnd), .vdd(vdd), .A(_1167_), .Y(_1167__bF_buf2) );
BUFX4 BUFX4_1129 ( .gnd(gnd), .vdd(vdd), .A(_1167_), .Y(_1167__bF_buf1) );
BUFX4 BUFX4_1130 ( .gnd(gnd), .vdd(vdd), .A(_1167_), .Y(_1167__bF_buf0) );
BUFX4 BUFX4_1131 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_7_), .Y(micro_hash_ucr_3_b_7_bF_buf3_) );
BUFX4 BUFX4_1132 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_7_), .Y(micro_hash_ucr_3_b_7_bF_buf2_) );
BUFX4 BUFX4_1133 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_7_), .Y(micro_hash_ucr_3_b_7_bF_buf1_) );
BUFX4 BUFX4_1134 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_7_), .Y(micro_hash_ucr_3_b_7_bF_buf0_) );
BUFX4 BUFX4_1135 ( .gnd(gnd), .vdd(vdd), .A(_3351_), .Y(_3351__bF_buf4) );
BUFX4 BUFX4_1136 ( .gnd(gnd), .vdd(vdd), .A(_3351_), .Y(_3351__bF_buf3) );
BUFX4 BUFX4_1137 ( .gnd(gnd), .vdd(vdd), .A(_3351_), .Y(_3351__bF_buf2) );
BUFX4 BUFX4_1138 ( .gnd(gnd), .vdd(vdd), .A(_3351_), .Y(_3351__bF_buf1) );
BUFX4 BUFX4_1139 ( .gnd(gnd), .vdd(vdd), .A(_3351_), .Y(_3351__bF_buf0) );
BUFX4 BUFX4_1140 ( .gnd(gnd), .vdd(vdd), .A(_4594_), .Y(_4594__bF_buf12) );
BUFX4 BUFX4_1141 ( .gnd(gnd), .vdd(vdd), .A(_4594_), .Y(_4594__bF_buf11) );
BUFX4 BUFX4_1142 ( .gnd(gnd), .vdd(vdd), .A(_4594_), .Y(_4594__bF_buf10) );
BUFX4 BUFX4_1143 ( .gnd(gnd), .vdd(vdd), .A(_4594_), .Y(_4594__bF_buf9) );
BUFX4 BUFX4_1144 ( .gnd(gnd), .vdd(vdd), .A(_4594_), .Y(_4594__bF_buf8) );
BUFX4 BUFX4_1145 ( .gnd(gnd), .vdd(vdd), .A(_4594_), .Y(_4594__bF_buf7) );
BUFX4 BUFX4_1146 ( .gnd(gnd), .vdd(vdd), .A(_4594_), .Y(_4594__bF_buf6) );
BUFX4 BUFX4_1147 ( .gnd(gnd), .vdd(vdd), .A(_4594_), .Y(_4594__bF_buf5) );
BUFX4 BUFX4_1148 ( .gnd(gnd), .vdd(vdd), .A(_4594_), .Y(_4594__bF_buf4) );
BUFX4 BUFX4_1149 ( .gnd(gnd), .vdd(vdd), .A(_4594_), .Y(_4594__bF_buf3) );
BUFX4 BUFX4_1150 ( .gnd(gnd), .vdd(vdd), .A(_4594_), .Y(_4594__bF_buf2) );
BUFX4 BUFX4_1151 ( .gnd(gnd), .vdd(vdd), .A(_4594_), .Y(_4594__bF_buf1) );
BUFX4 BUFX4_1152 ( .gnd(gnd), .vdd(vdd), .A(_4594_), .Y(_4594__bF_buf0) );
BUFX4 BUFX4_1153 ( .gnd(gnd), .vdd(vdd), .A(_880_), .Y(_880__bF_buf3) );
BUFX4 BUFX4_1154 ( .gnd(gnd), .vdd(vdd), .A(_880_), .Y(_880__bF_buf2) );
BUFX4 BUFX4_1155 ( .gnd(gnd), .vdd(vdd), .A(_880_), .Y(_880__bF_buf1) );
BUFX4 BUFX4_1156 ( .gnd(gnd), .vdd(vdd), .A(_880_), .Y(_880__bF_buf0) );
BUFX4 BUFX4_1157 ( .gnd(gnd), .vdd(vdd), .A(_460_), .Y(_460__bF_buf3) );
BUFX4 BUFX4_1158 ( .gnd(gnd), .vdd(vdd), .A(_460_), .Y(_460__bF_buf2) );
BUFX4 BUFX4_1159 ( .gnd(gnd), .vdd(vdd), .A(_460_), .Y(_460__bF_buf1) );
BUFX4 BUFX4_1160 ( .gnd(gnd), .vdd(vdd), .A(_460_), .Y(_460__bF_buf0) );
BUFX4 BUFX4_1161 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_0_), .Y(micro_hash_ucr_2_c_0_bF_buf3_) );
BUFX4 BUFX4_1162 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_0_), .Y(micro_hash_ucr_2_c_0_bF_buf2_) );
BUFX4 BUFX4_1163 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_0_), .Y(micro_hash_ucr_2_c_0_bF_buf1_) );
BUFX4 BUFX4_1164 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_0_), .Y(micro_hash_ucr_2_c_0_bF_buf0_) );
BUFX4 BUFX4_1165 ( .gnd(gnd), .vdd(vdd), .A(_5112_), .Y(_5112__bF_buf3) );
BUFX4 BUFX4_1166 ( .gnd(gnd), .vdd(vdd), .A(_5112_), .Y(_5112__bF_buf2) );
BUFX4 BUFX4_1167 ( .gnd(gnd), .vdd(vdd), .A(_5112_), .Y(_5112__bF_buf1) );
BUFX4 BUFX4_1168 ( .gnd(gnd), .vdd(vdd), .A(_5112_), .Y(_5112__bF_buf0) );
BUFX4 BUFX4_1169 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_3_), .Y(micro_hash_ucr_2_b_3_bF_buf3_) );
BUFX4 BUFX4_1170 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_3_), .Y(micro_hash_ucr_2_b_3_bF_buf2_) );
BUFX4 BUFX4_1171 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_3_), .Y(micro_hash_ucr_2_b_3_bF_buf1_) );
BUFX4 BUFX4_1172 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_3_), .Y(micro_hash_ucr_2_b_3_bF_buf0_) );
BUFX4 BUFX4_1173 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_1_), .Y(micro_hash_ucr_3_c_1_bF_buf3_) );
BUFX4 BUFX4_1174 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_1_), .Y(micro_hash_ucr_3_c_1_bF_buf2_) );
BUFX4 BUFX4_1175 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_1_), .Y(micro_hash_ucr_3_c_1_bF_buf1_) );
BUFX4 BUFX4_1176 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_1_), .Y(micro_hash_ucr_3_c_1_bF_buf0_) );
BUFX4 BUFX4_1177 ( .gnd(gnd), .vdd(vdd), .A(_9706_), .Y(_9706__bF_buf3) );
BUFX4 BUFX4_1178 ( .gnd(gnd), .vdd(vdd), .A(_9706_), .Y(_9706__bF_buf2) );
BUFX4 BUFX4_1179 ( .gnd(gnd), .vdd(vdd), .A(_9706_), .Y(_9706__bF_buf1) );
BUFX4 BUFX4_1180 ( .gnd(gnd), .vdd(vdd), .A(_9706_), .Y(_9706__bF_buf0) );
BUFX4 BUFX4_1181 ( .gnd(gnd), .vdd(vdd), .A(_877_), .Y(_877__bF_buf3) );
BUFX4 BUFX4_1182 ( .gnd(gnd), .vdd(vdd), .A(_877_), .Y(_877__bF_buf2) );
BUFX4 BUFX4_1183 ( .gnd(gnd), .vdd(vdd), .A(_877_), .Y(_877__bF_buf1) );
BUFX4 BUFX4_1184 ( .gnd(gnd), .vdd(vdd), .A(_877_), .Y(_877__bF_buf0) );
BUFX4 BUFX4_1185 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe30), .Y(micro_hash_ucr_3_pipe30_bF_buf4) );
BUFX4 BUFX4_1186 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe30), .Y(micro_hash_ucr_3_pipe30_bF_buf3) );
BUFX4 BUFX4_1187 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe30), .Y(micro_hash_ucr_3_pipe30_bF_buf2) );
BUFX4 BUFX4_1188 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe30), .Y(micro_hash_ucr_3_pipe30_bF_buf1) );
BUFX4 BUFX4_1189 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe30), .Y(micro_hash_ucr_3_pipe30_bF_buf0) );
BUFX4 BUFX4_1190 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe32), .Y(micro_hash_ucr_3_pipe32_bF_buf3) );
BUFX4 BUFX4_1191 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe32), .Y(micro_hash_ucr_3_pipe32_bF_buf2) );
BUFX4 BUFX4_1192 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe32), .Y(micro_hash_ucr_3_pipe32_bF_buf1) );
BUFX4 BUFX4_1193 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe32), .Y(micro_hash_ucr_3_pipe32_bF_buf0) );
BUFX4 BUFX4_1194 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe33), .Y(micro_hash_ucr_3_pipe33_bF_buf3) );
BUFX4 BUFX4_1195 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe33), .Y(micro_hash_ucr_3_pipe33_bF_buf2) );
BUFX4 BUFX4_1196 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe33), .Y(micro_hash_ucr_3_pipe33_bF_buf1) );
BUFX4 BUFX4_1197 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe33), .Y(micro_hash_ucr_3_pipe33_bF_buf0) );
BUFX4 BUFX4_1198 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe34), .Y(micro_hash_ucr_3_pipe34_bF_buf4) );
BUFX4 BUFX4_1199 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe34), .Y(micro_hash_ucr_3_pipe34_bF_buf3) );
BUFX4 BUFX4_1200 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe34), .Y(micro_hash_ucr_3_pipe34_bF_buf2) );
BUFX4 BUFX4_1201 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe34), .Y(micro_hash_ucr_3_pipe34_bF_buf1) );
BUFX4 BUFX4_1202 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe34), .Y(micro_hash_ucr_3_pipe34_bF_buf0) );
BUFX4 BUFX4_1203 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe35), .Y(micro_hash_ucr_3_pipe35_bF_buf3) );
BUFX4 BUFX4_1204 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe35), .Y(micro_hash_ucr_3_pipe35_bF_buf2) );
BUFX4 BUFX4_1205 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe35), .Y(micro_hash_ucr_3_pipe35_bF_buf1) );
BUFX4 BUFX4_1206 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe35), .Y(micro_hash_ucr_3_pipe35_bF_buf0) );
BUFX4 BUFX4_1207 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe36), .Y(micro_hash_ucr_3_pipe36_bF_buf4) );
BUFX4 BUFX4_1208 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe36), .Y(micro_hash_ucr_3_pipe36_bF_buf3) );
BUFX4 BUFX4_1209 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe36), .Y(micro_hash_ucr_3_pipe36_bF_buf2) );
BUFX4 BUFX4_1210 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe36), .Y(micro_hash_ucr_3_pipe36_bF_buf1) );
BUFX4 BUFX4_1211 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe36), .Y(micro_hash_ucr_3_pipe36_bF_buf0) );
BUFX4 BUFX4_1212 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe37), .Y(micro_hash_ucr_3_pipe37_bF_buf3) );
BUFX4 BUFX4_1213 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe37), .Y(micro_hash_ucr_3_pipe37_bF_buf2) );
BUFX4 BUFX4_1214 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe37), .Y(micro_hash_ucr_3_pipe37_bF_buf1) );
BUFX4 BUFX4_1215 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe37), .Y(micro_hash_ucr_3_pipe37_bF_buf0) );
BUFX4 BUFX4_1216 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe38), .Y(micro_hash_ucr_3_pipe38_bF_buf3) );
BUFX4 BUFX4_1217 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe38), .Y(micro_hash_ucr_3_pipe38_bF_buf2) );
BUFX4 BUFX4_1218 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe38), .Y(micro_hash_ucr_3_pipe38_bF_buf1) );
BUFX4 BUFX4_1219 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe38), .Y(micro_hash_ucr_3_pipe38_bF_buf0) );
BUFX4 BUFX4_1220 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe39), .Y(micro_hash_ucr_3_pipe39_bF_buf3) );
BUFX4 BUFX4_1221 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe39), .Y(micro_hash_ucr_3_pipe39_bF_buf2) );
BUFX4 BUFX4_1222 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe39), .Y(micro_hash_ucr_3_pipe39_bF_buf1) );
BUFX4 BUFX4_1223 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe39), .Y(micro_hash_ucr_3_pipe39_bF_buf0) );
BUFX4 BUFX4_1224 ( .gnd(gnd), .vdd(vdd), .A(_9324_), .Y(_9324__bF_buf4) );
BUFX4 BUFX4_1225 ( .gnd(gnd), .vdd(vdd), .A(_9324_), .Y(_9324__bF_buf3) );
BUFX4 BUFX4_1226 ( .gnd(gnd), .vdd(vdd), .A(_9324_), .Y(_9324__bF_buf2) );
BUFX4 BUFX4_1227 ( .gnd(gnd), .vdd(vdd), .A(_9324_), .Y(_9324__bF_buf1) );
BUFX4 BUFX4_1228 ( .gnd(gnd), .vdd(vdd), .A(_9324_), .Y(_9324__bF_buf0) );
BUFX4 BUFX4_1229 ( .gnd(gnd), .vdd(vdd), .A(comparador_valid), .Y(comparador_valid_bF_buf4) );
BUFX4 BUFX4_1230 ( .gnd(gnd), .vdd(vdd), .A(comparador_valid), .Y(comparador_valid_bF_buf3) );
BUFX4 BUFX4_1231 ( .gnd(gnd), .vdd(vdd), .A(comparador_valid), .Y(comparador_valid_bF_buf2) );
BUFX4 BUFX4_1232 ( .gnd(gnd), .vdd(vdd), .A(comparador_valid), .Y(comparador_valid_bF_buf1) );
BUFX4 BUFX4_1233 ( .gnd(gnd), .vdd(vdd), .A(comparador_valid), .Y(comparador_valid_bF_buf0) );
BUFX4 BUFX4_1234 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_6_), .Y(micro_hash_ucr_2_a_6_bF_buf3_) );
BUFX4 BUFX4_1235 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_6_), .Y(micro_hash_ucr_2_a_6_bF_buf2_) );
BUFX4 BUFX4_1236 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_6_), .Y(micro_hash_ucr_2_a_6_bF_buf1_) );
BUFX4 BUFX4_1237 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_6_), .Y(micro_hash_ucr_2_a_6_bF_buf0_) );
BUFX4 BUFX4_1238 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_4_), .Y(micro_hash_ucr_3_b_4_bF_buf4_) );
BUFX4 BUFX4_1239 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_4_), .Y(micro_hash_ucr_3_b_4_bF_buf3_) );
BUFX4 BUFX4_1240 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_4_), .Y(micro_hash_ucr_3_b_4_bF_buf2_) );
BUFX4 BUFX4_1241 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_4_), .Y(micro_hash_ucr_3_b_4_bF_buf1_) );
BUFX4 BUFX4_1242 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_4_), .Y(micro_hash_ucr_3_b_4_bF_buf0_) );
BUFX4 BUFX4_1243 ( .gnd(gnd), .vdd(vdd), .A(_5109_), .Y(_5109__bF_buf4) );
BUFX4 BUFX4_1244 ( .gnd(gnd), .vdd(vdd), .A(_5109_), .Y(_5109__bF_buf3) );
BUFX4 BUFX4_1245 ( .gnd(gnd), .vdd(vdd), .A(_5109_), .Y(_5109__bF_buf2) );
BUFX4 BUFX4_1246 ( .gnd(gnd), .vdd(vdd), .A(_5109_), .Y(_5109__bF_buf1) );
BUFX4 BUFX4_1247 ( .gnd(gnd), .vdd(vdd), .A(_5109_), .Y(_5109__bF_buf0) );
BUFX4 BUFX4_1248 ( .gnd(gnd), .vdd(vdd), .A(_5091_), .Y(_5091__bF_buf4) );
BUFX4 BUFX4_1249 ( .gnd(gnd), .vdd(vdd), .A(_5091_), .Y(_5091__bF_buf3) );
BUFX4 BUFX4_1250 ( .gnd(gnd), .vdd(vdd), .A(_5091_), .Y(_5091__bF_buf2) );
BUFX4 BUFX4_1251 ( .gnd(gnd), .vdd(vdd), .A(_5091_), .Y(_5091__bF_buf1) );
BUFX4 BUFX4_1252 ( .gnd(gnd), .vdd(vdd), .A(_5091_), .Y(_5091__bF_buf0) );
BUFX4 BUFX4_1253 ( .gnd(gnd), .vdd(vdd), .A(_8862_), .Y(_8862__bF_buf3) );
BUFX4 BUFX4_1254 ( .gnd(gnd), .vdd(vdd), .A(_8862_), .Y(_8862__bF_buf2) );
BUFX4 BUFX4_1255 ( .gnd(gnd), .vdd(vdd), .A(_8862_), .Y(_8862__bF_buf1) );
BUFX4 BUFX4_1256 ( .gnd(gnd), .vdd(vdd), .A(_8862_), .Y(_8862__bF_buf0) );
BUFX4 BUFX4_1257 ( .gnd(gnd), .vdd(vdd), .A(_12916__hier0_bF_buf5), .Y(_12916__bF_buf42) );
BUFX4 BUFX4_1258 ( .gnd(gnd), .vdd(vdd), .A(_12916__hier0_bF_buf4), .Y(_12916__bF_buf41) );
BUFX4 BUFX4_1259 ( .gnd(gnd), .vdd(vdd), .A(_12916__hier0_bF_buf3), .Y(_12916__bF_buf40) );
BUFX4 BUFX4_1260 ( .gnd(gnd), .vdd(vdd), .A(_12916__hier0_bF_buf2), .Y(_12916__bF_buf39) );
BUFX4 BUFX4_1261 ( .gnd(gnd), .vdd(vdd), .A(_12916__hier0_bF_buf1), .Y(_12916__bF_buf38) );
BUFX4 BUFX4_1262 ( .gnd(gnd), .vdd(vdd), .A(_12916__hier0_bF_buf0), .Y(_12916__bF_buf37) );
BUFX4 BUFX4_1263 ( .gnd(gnd), .vdd(vdd), .A(_12916__hier0_bF_buf5), .Y(_12916__bF_buf36) );
BUFX4 BUFX4_1264 ( .gnd(gnd), .vdd(vdd), .A(_12916__hier0_bF_buf4), .Y(_12916__bF_buf35) );
BUFX4 BUFX4_1265 ( .gnd(gnd), .vdd(vdd), .A(_12916__hier0_bF_buf3), .Y(_12916__bF_buf34) );
BUFX4 BUFX4_1266 ( .gnd(gnd), .vdd(vdd), .A(_12916__hier0_bF_buf2), .Y(_12916__bF_buf33) );
BUFX4 BUFX4_1267 ( .gnd(gnd), .vdd(vdd), .A(_12916__hier0_bF_buf1), .Y(_12916__bF_buf32) );
BUFX4 BUFX4_1268 ( .gnd(gnd), .vdd(vdd), .A(_12916__hier0_bF_buf0), .Y(_12916__bF_buf31) );
BUFX4 BUFX4_1269 ( .gnd(gnd), .vdd(vdd), .A(_12916__hier0_bF_buf5), .Y(_12916__bF_buf30) );
BUFX4 BUFX4_1270 ( .gnd(gnd), .vdd(vdd), .A(_12916__hier0_bF_buf4), .Y(_12916__bF_buf29) );
BUFX4 BUFX4_1271 ( .gnd(gnd), .vdd(vdd), .A(_12916__hier0_bF_buf3), .Y(_12916__bF_buf28) );
BUFX4 BUFX4_1272 ( .gnd(gnd), .vdd(vdd), .A(_12916__hier0_bF_buf2), .Y(_12916__bF_buf27) );
BUFX4 BUFX4_1273 ( .gnd(gnd), .vdd(vdd), .A(_12916__hier0_bF_buf1), .Y(_12916__bF_buf26) );
BUFX4 BUFX4_1274 ( .gnd(gnd), .vdd(vdd), .A(_12916__hier0_bF_buf0), .Y(_12916__bF_buf25) );
BUFX4 BUFX4_1275 ( .gnd(gnd), .vdd(vdd), .A(_12916__hier0_bF_buf5), .Y(_12916__bF_buf24) );
BUFX4 BUFX4_1276 ( .gnd(gnd), .vdd(vdd), .A(_12916__hier0_bF_buf4), .Y(_12916__bF_buf23) );
BUFX4 BUFX4_1277 ( .gnd(gnd), .vdd(vdd), .A(_12916__hier0_bF_buf3), .Y(_12916__bF_buf22) );
BUFX4 BUFX4_1278 ( .gnd(gnd), .vdd(vdd), .A(_12916__hier0_bF_buf2), .Y(_12916__bF_buf21) );
BUFX4 BUFX4_1279 ( .gnd(gnd), .vdd(vdd), .A(_12916__hier0_bF_buf1), .Y(_12916__bF_buf20) );
BUFX4 BUFX4_1280 ( .gnd(gnd), .vdd(vdd), .A(_12916__hier0_bF_buf0), .Y(_12916__bF_buf19) );
BUFX4 BUFX4_1281 ( .gnd(gnd), .vdd(vdd), .A(_12916__hier0_bF_buf5), .Y(_12916__bF_buf18) );
BUFX4 BUFX4_1282 ( .gnd(gnd), .vdd(vdd), .A(_12916__hier0_bF_buf4), .Y(_12916__bF_buf17) );
BUFX4 BUFX4_1283 ( .gnd(gnd), .vdd(vdd), .A(_12916__hier0_bF_buf3), .Y(_12916__bF_buf16) );
BUFX4 BUFX4_1284 ( .gnd(gnd), .vdd(vdd), .A(_12916__hier0_bF_buf2), .Y(_12916__bF_buf15) );
BUFX4 BUFX4_1285 ( .gnd(gnd), .vdd(vdd), .A(_12916__hier0_bF_buf1), .Y(_12916__bF_buf14) );
BUFX4 BUFX4_1286 ( .gnd(gnd), .vdd(vdd), .A(_12916__hier0_bF_buf0), .Y(_12916__bF_buf13) );
BUFX4 BUFX4_1287 ( .gnd(gnd), .vdd(vdd), .A(_12916__hier0_bF_buf5), .Y(_12916__bF_buf12) );
BUFX4 BUFX4_1288 ( .gnd(gnd), .vdd(vdd), .A(_12916__hier0_bF_buf4), .Y(_12916__bF_buf11) );
BUFX4 BUFX4_1289 ( .gnd(gnd), .vdd(vdd), .A(_12916__hier0_bF_buf3), .Y(_12916__bF_buf10) );
BUFX4 BUFX4_1290 ( .gnd(gnd), .vdd(vdd), .A(_12916__hier0_bF_buf2), .Y(_12916__bF_buf9) );
BUFX4 BUFX4_1291 ( .gnd(gnd), .vdd(vdd), .A(_12916__hier0_bF_buf1), .Y(_12916__bF_buf8) );
BUFX4 BUFX4_1292 ( .gnd(gnd), .vdd(vdd), .A(_12916__hier0_bF_buf0), .Y(_12916__bF_buf7) );
BUFX4 BUFX4_1293 ( .gnd(gnd), .vdd(vdd), .A(_12916__hier0_bF_buf5), .Y(_12916__bF_buf6) );
BUFX4 BUFX4_1294 ( .gnd(gnd), .vdd(vdd), .A(_12916__hier0_bF_buf4), .Y(_12916__bF_buf5) );
BUFX4 BUFX4_1295 ( .gnd(gnd), .vdd(vdd), .A(_12916__hier0_bF_buf3), .Y(_12916__bF_buf4) );
BUFX4 BUFX4_1296 ( .gnd(gnd), .vdd(vdd), .A(_12916__hier0_bF_buf2), .Y(_12916__bF_buf3) );
BUFX4 BUFX4_1297 ( .gnd(gnd), .vdd(vdd), .A(_12916__hier0_bF_buf1), .Y(_12916__bF_buf2) );
BUFX4 BUFX4_1298 ( .gnd(gnd), .vdd(vdd), .A(_12916__hier0_bF_buf0), .Y(_12916__bF_buf1) );
BUFX4 BUFX4_1299 ( .gnd(gnd), .vdd(vdd), .A(_12916__hier0_bF_buf5), .Y(_12916__bF_buf0) );
BUFX4 BUFX4_1300 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_7_), .Y(micro_hash_ucr_3_a_7_bF_buf3_) );
BUFX4 BUFX4_1301 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_7_), .Y(micro_hash_ucr_3_a_7_bF_buf2_) );
BUFX4 BUFX4_1302 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_7_), .Y(micro_hash_ucr_3_a_7_bF_buf1_) );
BUFX4 BUFX4_1303 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_7_), .Y(micro_hash_ucr_3_a_7_bF_buf0_) );
BUFX4 BUFX4_1304 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_0_), .Y(micro_hash_ucr_2_b_0_bF_buf3_) );
BUFX4 BUFX4_1305 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_0_), .Y(micro_hash_ucr_2_b_0_bF_buf2_) );
BUFX4 BUFX4_1306 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_0_), .Y(micro_hash_ucr_2_b_0_bF_buf1_) );
BUFX4 BUFX4_1307 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_0_), .Y(micro_hash_ucr_2_b_0_bF_buf0_) );
BUFX4 BUFX4_1308 ( .gnd(gnd), .vdd(vdd), .A(_9321_), .Y(_9321__bF_buf3) );
BUFX4 BUFX4_1309 ( .gnd(gnd), .vdd(vdd), .A(_9321_), .Y(_9321__bF_buf2) );
BUFX4 BUFX4_1310 ( .gnd(gnd), .vdd(vdd), .A(_9321_), .Y(_9321__bF_buf1) );
BUFX4 BUFX4_1311 ( .gnd(gnd), .vdd(vdd), .A(_9321_), .Y(_9321__bF_buf0) );
BUFX4 BUFX4_1312 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_1_), .Y(micro_hash_ucr_3_b_1_bF_buf3_) );
BUFX4 BUFX4_1313 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_1_), .Y(micro_hash_ucr_3_b_1_bF_buf2_) );
BUFX4 BUFX4_1314 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_1_), .Y(micro_hash_ucr_3_b_1_bF_buf1_) );
BUFX4 BUFX4_1315 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_1_), .Y(micro_hash_ucr_3_b_1_bF_buf0_) );
BUFX4 BUFX4_1316 ( .gnd(gnd), .vdd(vdd), .A(_6293_), .Y(_6293__bF_buf4) );
BUFX4 BUFX4_1317 ( .gnd(gnd), .vdd(vdd), .A(_6293_), .Y(_6293__bF_buf3) );
BUFX4 BUFX4_1318 ( .gnd(gnd), .vdd(vdd), .A(_6293_), .Y(_6293__bF_buf2) );
BUFX4 BUFX4_1319 ( .gnd(gnd), .vdd(vdd), .A(_6293_), .Y(_6293__bF_buf1) );
BUFX4 BUFX4_1320 ( .gnd(gnd), .vdd(vdd), .A(_6293_), .Y(_6293__bF_buf0) );
BUFX4 BUFX4_1321 ( .gnd(gnd), .vdd(vdd), .A(_10996_), .Y(_10996__bF_buf4) );
BUFX4 BUFX4_1322 ( .gnd(gnd), .vdd(vdd), .A(_10996_), .Y(_10996__bF_buf3) );
BUFX4 BUFX4_1323 ( .gnd(gnd), .vdd(vdd), .A(_10996_), .Y(_10996__bF_buf2) );
BUFX4 BUFX4_1324 ( .gnd(gnd), .vdd(vdd), .A(_10996_), .Y(_10996__bF_buf1) );
BUFX4 BUFX4_1325 ( .gnd(gnd), .vdd(vdd), .A(_10996_), .Y(_10996__bF_buf0) );
BUFX4 BUFX4_1326 ( .gnd(gnd), .vdd(vdd), .A(_9318_), .Y(_9318__bF_buf4) );
BUFX4 BUFX4_1327 ( .gnd(gnd), .vdd(vdd), .A(_9318_), .Y(_9318__bF_buf3) );
BUFX4 BUFX4_1328 ( .gnd(gnd), .vdd(vdd), .A(_9318_), .Y(_9318__bF_buf2) );
BUFX4 BUFX4_1329 ( .gnd(gnd), .vdd(vdd), .A(_9318_), .Y(_9318__bF_buf1) );
BUFX4 BUFX4_1330 ( .gnd(gnd), .vdd(vdd), .A(_9318_), .Y(_9318__bF_buf0) );
BUFX4 BUFX4_1331 ( .gnd(gnd), .vdd(vdd), .A(_930_), .Y(_930__bF_buf4) );
BUFX4 BUFX4_1332 ( .gnd(gnd), .vdd(vdd), .A(_930_), .Y(_930__bF_buf3) );
BUFX4 BUFX4_1333 ( .gnd(gnd), .vdd(vdd), .A(_930_), .Y(_930__bF_buf2) );
BUFX4 BUFX4_1334 ( .gnd(gnd), .vdd(vdd), .A(_930_), .Y(_930__bF_buf1) );
BUFX4 BUFX4_1335 ( .gnd(gnd), .vdd(vdd), .A(_930_), .Y(_930__bF_buf0) );
BUFX4 BUFX4_1336 ( .gnd(gnd), .vdd(vdd), .A(_5085_), .Y(_5085__bF_buf3) );
BUFX4 BUFX4_1337 ( .gnd(gnd), .vdd(vdd), .A(_5085_), .Y(_5085__bF_buf2) );
BUFX4 BUFX4_1338 ( .gnd(gnd), .vdd(vdd), .A(_5085_), .Y(_5085__bF_buf1) );
BUFX4 BUFX4_1339 ( .gnd(gnd), .vdd(vdd), .A(_5085_), .Y(_5085__bF_buf0) );
BUFX4 BUFX4_1340 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe60), .Y(micro_hash_ucr_pipe60_bF_buf4) );
BUFX4 BUFX4_1341 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe60), .Y(micro_hash_ucr_pipe60_bF_buf3) );
BUFX4 BUFX4_1342 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe60), .Y(micro_hash_ucr_pipe60_bF_buf2) );
BUFX4 BUFX4_1343 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe60), .Y(micro_hash_ucr_pipe60_bF_buf1) );
BUFX4 BUFX4_1344 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe60), .Y(micro_hash_ucr_pipe60_bF_buf0) );
BUFX4 BUFX4_1345 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe61), .Y(micro_hash_ucr_pipe61_bF_buf3) );
BUFX4 BUFX4_1346 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe61), .Y(micro_hash_ucr_pipe61_bF_buf2) );
BUFX4 BUFX4_1347 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe61), .Y(micro_hash_ucr_pipe61_bF_buf1) );
BUFX4 BUFX4_1348 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe61), .Y(micro_hash_ucr_pipe61_bF_buf0) );
BUFX4 BUFX4_1349 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe62), .Y(micro_hash_ucr_pipe62_bF_buf4) );
BUFX4 BUFX4_1350 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe62), .Y(micro_hash_ucr_pipe62_bF_buf3) );
BUFX4 BUFX4_1351 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe62), .Y(micro_hash_ucr_pipe62_bF_buf2) );
BUFX4 BUFX4_1352 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe62), .Y(micro_hash_ucr_pipe62_bF_buf1) );
BUFX4 BUFX4_1353 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe62), .Y(micro_hash_ucr_pipe62_bF_buf0) );
BUFX4 BUFX4_1354 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe64), .Y(micro_hash_ucr_pipe64_bF_buf4) );
BUFX4 BUFX4_1355 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe64), .Y(micro_hash_ucr_pipe64_bF_buf3) );
BUFX4 BUFX4_1356 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe64), .Y(micro_hash_ucr_pipe64_bF_buf2) );
BUFX4 BUFX4_1357 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe64), .Y(micro_hash_ucr_pipe64_bF_buf1) );
BUFX4 BUFX4_1358 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe64), .Y(micro_hash_ucr_pipe64_bF_buf0) );
BUFX4 BUFX4_1359 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe65), .Y(micro_hash_ucr_pipe65_bF_buf3) );
BUFX4 BUFX4_1360 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe65), .Y(micro_hash_ucr_pipe65_bF_buf2) );
BUFX4 BUFX4_1361 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe65), .Y(micro_hash_ucr_pipe65_bF_buf1) );
BUFX4 BUFX4_1362 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe65), .Y(micro_hash_ucr_pipe65_bF_buf0) );
BUFX4 BUFX4_1363 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe66), .Y(micro_hash_ucr_pipe66_bF_buf4) );
BUFX4 BUFX4_1364 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe66), .Y(micro_hash_ucr_pipe66_bF_buf3) );
BUFX4 BUFX4_1365 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe66), .Y(micro_hash_ucr_pipe66_bF_buf2) );
BUFX4 BUFX4_1366 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe66), .Y(micro_hash_ucr_pipe66_bF_buf1) );
BUFX4 BUFX4_1367 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe66), .Y(micro_hash_ucr_pipe66_bF_buf0) );
BUFX4 BUFX4_1368 ( .gnd(gnd), .vdd(vdd), .A(_927_), .Y(_927__bF_buf3) );
BUFX4 BUFX4_1369 ( .gnd(gnd), .vdd(vdd), .A(_927_), .Y(_927__bF_buf2) );
BUFX4 BUFX4_1370 ( .gnd(gnd), .vdd(vdd), .A(_927_), .Y(_927__bF_buf1) );
BUFX4 BUFX4_1371 ( .gnd(gnd), .vdd(vdd), .A(_927_), .Y(_927__bF_buf0) );
BUFX4 BUFX4_1372 ( .gnd(gnd), .vdd(vdd), .A(_5103_), .Y(_5103__bF_buf3) );
BUFX4 BUFX4_1373 ( .gnd(gnd), .vdd(vdd), .A(_5103_), .Y(_5103__bF_buf2) );
BUFX4 BUFX4_1374 ( .gnd(gnd), .vdd(vdd), .A(_5103_), .Y(_5103__bF_buf1) );
BUFX4 BUFX4_1375 ( .gnd(gnd), .vdd(vdd), .A(_5103_), .Y(_5103__bF_buf0) );
BUFX4 BUFX4_1376 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_1_), .Y(micro_hash_ucr_3_a_1_bF_buf3_) );
BUFX4 BUFX4_1377 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_1_), .Y(micro_hash_ucr_3_a_1_bF_buf2_) );
BUFX4 BUFX4_1378 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_1_), .Y(micro_hash_ucr_3_a_1_bF_buf1_) );
BUFX4 BUFX4_1379 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_1_), .Y(micro_hash_ucr_3_a_1_bF_buf0_) );
BUFX4 BUFX4_1380 ( .gnd(gnd), .vdd(vdd), .A(_1957_), .Y(_1957__bF_buf3) );
BUFX4 BUFX4_1381 ( .gnd(gnd), .vdd(vdd), .A(_1957_), .Y(_1957__bF_buf2) );
BUFX4 BUFX4_1382 ( .gnd(gnd), .vdd(vdd), .A(_1957_), .Y(_1957__bF_buf1) );
BUFX4 BUFX4_1383 ( .gnd(gnd), .vdd(vdd), .A(_1957_), .Y(_1957__bF_buf0) );
BUFX4 BUFX4_1384 ( .gnd(gnd), .vdd(vdd), .A(_1290_), .Y(_1290__bF_buf3) );
BUFX4 BUFX4_1385 ( .gnd(gnd), .vdd(vdd), .A(_1290_), .Y(_1290__bF_buf2) );
BUFX4 BUFX4_1386 ( .gnd(gnd), .vdd(vdd), .A(_1290_), .Y(_1290__bF_buf1) );
BUFX4 BUFX4_1387 ( .gnd(gnd), .vdd(vdd), .A(_1290_), .Y(_1290__bF_buf0) );
BUFX4 BUFX4_1388 ( .gnd(gnd), .vdd(vdd), .A(_1058_), .Y(_1058__bF_buf3) );
BUFX4 BUFX4_1389 ( .gnd(gnd), .vdd(vdd), .A(_1058_), .Y(_1058__bF_buf2) );
BUFX4 BUFX4_1390 ( .gnd(gnd), .vdd(vdd), .A(_1058_), .Y(_1058__bF_buf1) );
BUFX4 BUFX4_1391 ( .gnd(gnd), .vdd(vdd), .A(_1058_), .Y(_1058__bF_buf0) );
BUFX4 BUFX4_1392 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe30), .Y(micro_hash_ucr_pipe30_bF_buf3) );
BUFX4 BUFX4_1393 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe30), .Y(micro_hash_ucr_pipe30_bF_buf2) );
BUFX4 BUFX4_1394 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe30), .Y(micro_hash_ucr_pipe30_bF_buf1) );
BUFX4 BUFX4_1395 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe30), .Y(micro_hash_ucr_pipe30_bF_buf0) );
BUFX4 BUFX4_1396 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe32), .Y(micro_hash_ucr_pipe32_bF_buf3) );
BUFX4 BUFX4_1397 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe32), .Y(micro_hash_ucr_pipe32_bF_buf2) );
BUFX4 BUFX4_1398 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe32), .Y(micro_hash_ucr_pipe32_bF_buf1) );
BUFX4 BUFX4_1399 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe32), .Y(micro_hash_ucr_pipe32_bF_buf0) );
BUFX4 BUFX4_1400 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe33), .Y(micro_hash_ucr_pipe33_bF_buf3) );
BUFX4 BUFX4_1401 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe33), .Y(micro_hash_ucr_pipe33_bF_buf2) );
BUFX4 BUFX4_1402 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe33), .Y(micro_hash_ucr_pipe33_bF_buf1) );
BUFX4 BUFX4_1403 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe33), .Y(micro_hash_ucr_pipe33_bF_buf0) );
BUFX4 BUFX4_1404 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe34), .Y(micro_hash_ucr_pipe34_bF_buf3) );
BUFX4 BUFX4_1405 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe34), .Y(micro_hash_ucr_pipe34_bF_buf2) );
BUFX4 BUFX4_1406 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe34), .Y(micro_hash_ucr_pipe34_bF_buf1) );
BUFX4 BUFX4_1407 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe34), .Y(micro_hash_ucr_pipe34_bF_buf0) );
BUFX4 BUFX4_1408 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe36), .Y(micro_hash_ucr_pipe36_bF_buf3) );
BUFX4 BUFX4_1409 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe36), .Y(micro_hash_ucr_pipe36_bF_buf2) );
BUFX4 BUFX4_1410 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe36), .Y(micro_hash_ucr_pipe36_bF_buf1) );
BUFX4 BUFX4_1411 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe36), .Y(micro_hash_ucr_pipe36_bF_buf0) );
BUFX4 BUFX4_1412 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe38), .Y(micro_hash_ucr_pipe38_bF_buf3) );
BUFX4 BUFX4_1413 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe38), .Y(micro_hash_ucr_pipe38_bF_buf2) );
BUFX4 BUFX4_1414 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe38), .Y(micro_hash_ucr_pipe38_bF_buf1) );
BUFX4 BUFX4_1415 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe38), .Y(micro_hash_ucr_pipe38_bF_buf0) );
BUFX4 BUFX4_1416 ( .gnd(gnd), .vdd(vdd), .A(_9294_), .Y(_9294__bF_buf4) );
BUFX4 BUFX4_1417 ( .gnd(gnd), .vdd(vdd), .A(_9294_), .Y(_9294__bF_buf3) );
BUFX4 BUFX4_1418 ( .gnd(gnd), .vdd(vdd), .A(_9294_), .Y(_9294__bF_buf2) );
BUFX4 BUFX4_1419 ( .gnd(gnd), .vdd(vdd), .A(_9294_), .Y(_9294__bF_buf1) );
BUFX4 BUFX4_1420 ( .gnd(gnd), .vdd(vdd), .A(_9294_), .Y(_9294__bF_buf0) );
BUFX4 BUFX4_1421 ( .gnd(gnd), .vdd(vdd), .A(_2322_), .Y(_2322__bF_buf5) );
BUFX4 BUFX4_1422 ( .gnd(gnd), .vdd(vdd), .A(_2322_), .Y(_2322__bF_buf4) );
BUFX4 BUFX4_1423 ( .gnd(gnd), .vdd(vdd), .A(_2322_), .Y(_2322__bF_buf3) );
BUFX4 BUFX4_1424 ( .gnd(gnd), .vdd(vdd), .A(_2322_), .Y(_2322__bF_buf2) );
BUFX4 BUFX4_1425 ( .gnd(gnd), .vdd(vdd), .A(_2322_), .Y(_2322__bF_buf1) );
BUFX4 BUFX4_1426 ( .gnd(gnd), .vdd(vdd), .A(_2322_), .Y(_2322__bF_buf0) );
BUFX4 BUFX4_1427 ( .gnd(gnd), .vdd(vdd), .A(_3107_), .Y(_3107__bF_buf3) );
BUFX4 BUFX4_1428 ( .gnd(gnd), .vdd(vdd), .A(_3107_), .Y(_3107__bF_buf2) );
BUFX4 BUFX4_1429 ( .gnd(gnd), .vdd(vdd), .A(_3107_), .Y(_3107__bF_buf1) );
BUFX4 BUFX4_1430 ( .gnd(gnd), .vdd(vdd), .A(_3107_), .Y(_3107__bF_buf0) );
BUFX4 BUFX4_1431 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_1_), .Y(micro_hash_ucr_c_1_bF_buf3_) );
BUFX4 BUFX4_1432 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_1_), .Y(micro_hash_ucr_c_1_bF_buf2_) );
BUFX4 BUFX4_1433 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_1_), .Y(micro_hash_ucr_c_1_bF_buf1_) );
BUFX4 BUFX4_1434 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_1_), .Y(micro_hash_ucr_c_1_bF_buf0_) );
BUFX4 BUFX4_1435 ( .gnd(gnd), .vdd(vdd), .A(_924_), .Y(_924__bF_buf4) );
BUFX4 BUFX4_1436 ( .gnd(gnd), .vdd(vdd), .A(_924_), .Y(_924__bF_buf3) );
BUFX4 BUFX4_1437 ( .gnd(gnd), .vdd(vdd), .A(_924_), .Y(_924__bF_buf2) );
BUFX4 BUFX4_1438 ( .gnd(gnd), .vdd(vdd), .A(_924_), .Y(_924__bF_buf1) );
BUFX4 BUFX4_1439 ( .gnd(gnd), .vdd(vdd), .A(_924_), .Y(_924__bF_buf0) );
BUFX4 BUFX4_1440 ( .gnd(gnd), .vdd(vdd), .A(_1402_), .Y(_1402__bF_buf3) );
BUFX4 BUFX4_1441 ( .gnd(gnd), .vdd(vdd), .A(_1402_), .Y(_1402__bF_buf2) );
BUFX4 BUFX4_1442 ( .gnd(gnd), .vdd(vdd), .A(_1402_), .Y(_1402__bF_buf1) );
BUFX4 BUFX4_1443 ( .gnd(gnd), .vdd(vdd), .A(_1402_), .Y(_1402__bF_buf0) );
BUFX4 BUFX4_1444 ( .gnd(gnd), .vdd(vdd), .A(_5079_), .Y(_5079__bF_buf4) );
BUFX4 BUFX4_1445 ( .gnd(gnd), .vdd(vdd), .A(_5079_), .Y(_5079__bF_buf3) );
BUFX4 BUFX4_1446 ( .gnd(gnd), .vdd(vdd), .A(_5079_), .Y(_5079__bF_buf2) );
BUFX4 BUFX4_1447 ( .gnd(gnd), .vdd(vdd), .A(_5079_), .Y(_5079__bF_buf1) );
BUFX4 BUFX4_1448 ( .gnd(gnd), .vdd(vdd), .A(_5079_), .Y(_5079__bF_buf0) );
BUFX4 BUFX4_1449 ( .gnd(gnd), .vdd(vdd), .A(_12848_), .Y(_12848__bF_buf3) );
BUFX4 BUFX4_1450 ( .gnd(gnd), .vdd(vdd), .A(_12848_), .Y(_12848__bF_buf2) );
BUFX4 BUFX4_1451 ( .gnd(gnd), .vdd(vdd), .A(_12848_), .Y(_12848__bF_buf1) );
BUFX4 BUFX4_1452 ( .gnd(gnd), .vdd(vdd), .A(_12848_), .Y(_12848__bF_buf0) );
BUFX4 BUFX4_1453 ( .gnd(gnd), .vdd(vdd), .A(_5100_), .Y(_5100__bF_buf3) );
BUFX4 BUFX4_1454 ( .gnd(gnd), .vdd(vdd), .A(_5100_), .Y(_5100__bF_buf2) );
BUFX4 BUFX4_1455 ( .gnd(gnd), .vdd(vdd), .A(_5100_), .Y(_5100__bF_buf1) );
BUFX4 BUFX4_1456 ( .gnd(gnd), .vdd(vdd), .A(_5100_), .Y(_5100__bF_buf0) );
BUFX4 BUFX4_1457 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_4_), .Y(micro_hash_ucr_b_4_bF_buf3_) );
BUFX4 BUFX4_1458 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_4_), .Y(micro_hash_ucr_b_4_bF_buf2_) );
BUFX4 BUFX4_1459 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_4_), .Y(micro_hash_ucr_b_4_bF_buf1_) );
BUFX4 BUFX4_1460 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_4_), .Y(micro_hash_ucr_b_4_bF_buf0_) );
BUFX4 BUFX4_1461 ( .gnd(gnd), .vdd(vdd), .A(_1725_), .Y(_1725__bF_buf3) );
BUFX4 BUFX4_1462 ( .gnd(gnd), .vdd(vdd), .A(_1725_), .Y(_1725__bF_buf2) );
BUFX4 BUFX4_1463 ( .gnd(gnd), .vdd(vdd), .A(_1725_), .Y(_1725__bF_buf1) );
BUFX4 BUFX4_1464 ( .gnd(gnd), .vdd(vdd), .A(_1725_), .Y(_1725__bF_buf0) );
BUFX4 BUFX4_1465 ( .gnd(gnd), .vdd(vdd), .A(_9312_), .Y(_9312__bF_buf3) );
BUFX4 BUFX4_1466 ( .gnd(gnd), .vdd(vdd), .A(_9312_), .Y(_9312__bF_buf2) );
BUFX4 BUFX4_1467 ( .gnd(gnd), .vdd(vdd), .A(_9312_), .Y(_9312__bF_buf1) );
BUFX4 BUFX4_1468 ( .gnd(gnd), .vdd(vdd), .A(_9312_), .Y(_9312__bF_buf0) );
BUFX4 BUFX4_1469 ( .gnd(gnd), .vdd(vdd), .A(_9309_), .Y(_9309__bF_buf3) );
BUFX4 BUFX4_1470 ( .gnd(gnd), .vdd(vdd), .A(_9309_), .Y(_9309__bF_buf2) );
BUFX4 BUFX4_1471 ( .gnd(gnd), .vdd(vdd), .A(_9309_), .Y(_9309__bF_buf1) );
BUFX4 BUFX4_1472 ( .gnd(gnd), .vdd(vdd), .A(_9309_), .Y(_9309__bF_buf0) );
BUFX4 BUFX4_1473 ( .gnd(gnd), .vdd(vdd), .A(_921_), .Y(_921__bF_buf3) );
BUFX4 BUFX4_1474 ( .gnd(gnd), .vdd(vdd), .A(_921_), .Y(_921__bF_buf2) );
BUFX4 BUFX4_1475 ( .gnd(gnd), .vdd(vdd), .A(_921_), .Y(_921__bF_buf1) );
BUFX4 BUFX4_1476 ( .gnd(gnd), .vdd(vdd), .A(_921_), .Y(_921__bF_buf0) );
BUFX4 BUFX4_1477 ( .gnd(gnd), .vdd(vdd), .A(_5076_), .Y(_5076__bF_buf3) );
BUFX4 BUFX4_1478 ( .gnd(gnd), .vdd(vdd), .A(_5076_), .Y(_5076__bF_buf2) );
BUFX4 BUFX4_1479 ( .gnd(gnd), .vdd(vdd), .A(_5076_), .Y(_5076__bF_buf1) );
BUFX4 BUFX4_1480 ( .gnd(gnd), .vdd(vdd), .A(_5076_), .Y(_5076__bF_buf0) );
BUFX4 BUFX4_1481 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_1_), .Y(micro_hash_ucr_b_1_bF_buf3_) );
BUFX4 BUFX4_1482 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_1_), .Y(micro_hash_ucr_b_1_bF_buf2_) );
BUFX4 BUFX4_1483 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_1_), .Y(micro_hash_ucr_b_1_bF_buf1_) );
BUFX4 BUFX4_1484 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_1_), .Y(micro_hash_ucr_b_1_bF_buf0_) );
BUFX4 BUFX4_1485 ( .gnd(gnd), .vdd(vdd), .A(_7316_), .Y(_7316__bF_buf3) );
BUFX4 BUFX4_1486 ( .gnd(gnd), .vdd(vdd), .A(_7316_), .Y(_7316__bF_buf2) );
BUFX4 BUFX4_1487 ( .gnd(gnd), .vdd(vdd), .A(_7316_), .Y(_7316__bF_buf1) );
BUFX4 BUFX4_1488 ( .gnd(gnd), .vdd(vdd), .A(_7316_), .Y(_7316__bF_buf0) );
BUFX4 BUFX4_1489 ( .gnd(gnd), .vdd(vdd), .A(_11543_), .Y(_11543__bF_buf3) );
BUFX4 BUFX4_1490 ( .gnd(gnd), .vdd(vdd), .A(_11543_), .Y(_11543__bF_buf2) );
BUFX4 BUFX4_1491 ( .gnd(gnd), .vdd(vdd), .A(_11543_), .Y(_11543__bF_buf1) );
BUFX4 BUFX4_1492 ( .gnd(gnd), .vdd(vdd), .A(_11543_), .Y(_11543__bF_buf0) );
BUFX4 BUFX4_1493 ( .gnd(gnd), .vdd(vdd), .A(_9288_), .Y(_9288__bF_buf3) );
BUFX4 BUFX4_1494 ( .gnd(gnd), .vdd(vdd), .A(_9288_), .Y(_9288__bF_buf2) );
BUFX4 BUFX4_1495 ( .gnd(gnd), .vdd(vdd), .A(_9288_), .Y(_9288__bF_buf1) );
BUFX4 BUFX4_1496 ( .gnd(gnd), .vdd(vdd), .A(_9288_), .Y(_9288__bF_buf0) );
BUFX4 BUFX4_1497 ( .gnd(gnd), .vdd(vdd), .A(_4479_), .Y(_4479__bF_buf3) );
BUFX4 BUFX4_1498 ( .gnd(gnd), .vdd(vdd), .A(_4479_), .Y(_4479__bF_buf2) );
BUFX4 BUFX4_1499 ( .gnd(gnd), .vdd(vdd), .A(_4479_), .Y(_4479__bF_buf1) );
BUFX4 BUFX4_1500 ( .gnd(gnd), .vdd(vdd), .A(_4479_), .Y(_4479__bF_buf0) );
BUFX4 BUFX4_1501 ( .gnd(gnd), .vdd(vdd), .A(_918_), .Y(_918__bF_buf4) );
BUFX4 BUFX4_1502 ( .gnd(gnd), .vdd(vdd), .A(_918_), .Y(_918__bF_buf3) );
BUFX4 BUFX4_1503 ( .gnd(gnd), .vdd(vdd), .A(_918_), .Y(_918__bF_buf2) );
BUFX4 BUFX4_1504 ( .gnd(gnd), .vdd(vdd), .A(_918_), .Y(_918__bF_buf1) );
BUFX4 BUFX4_1505 ( .gnd(gnd), .vdd(vdd), .A(_918_), .Y(_918__bF_buf0) );
BUFX4 BUFX4_1506 ( .gnd(gnd), .vdd(vdd), .A(_5705_), .Y(_5705__bF_buf3) );
BUFX4 BUFX4_1507 ( .gnd(gnd), .vdd(vdd), .A(_5705_), .Y(_5705__bF_buf2) );
BUFX4 BUFX4_1508 ( .gnd(gnd), .vdd(vdd), .A(_5705_), .Y(_5705__bF_buf1) );
BUFX4 BUFX4_1509 ( .gnd(gnd), .vdd(vdd), .A(_5705_), .Y(_5705__bF_buf0) );
BUFX4 BUFX4_1510 ( .gnd(gnd), .vdd(vdd), .A(_8903_), .Y(_8903__bF_buf3) );
BUFX4 BUFX4_1511 ( .gnd(gnd), .vdd(vdd), .A(_8903_), .Y(_8903__bF_buf2) );
BUFX4 BUFX4_1512 ( .gnd(gnd), .vdd(vdd), .A(_8903_), .Y(_8903__bF_buf1) );
BUFX4 BUFX4_1513 ( .gnd(gnd), .vdd(vdd), .A(_8903_), .Y(_8903__bF_buf0) );
BUFX4 BUFX4_1514 ( .gnd(gnd), .vdd(vdd), .A(_9306_), .Y(_9306__bF_buf3) );
BUFX4 BUFX4_1515 ( .gnd(gnd), .vdd(vdd), .A(_9306_), .Y(_9306__bF_buf2) );
BUFX4 BUFX4_1516 ( .gnd(gnd), .vdd(vdd), .A(_9306_), .Y(_9306__bF_buf1) );
BUFX4 BUFX4_1517 ( .gnd(gnd), .vdd(vdd), .A(_9306_), .Y(_9306__bF_buf0) );
BUFX4 BUFX4_1518 ( .gnd(gnd), .vdd(vdd), .A(_897_), .Y(_897__bF_buf3) );
BUFX4 BUFX4_1519 ( .gnd(gnd), .vdd(vdd), .A(_897_), .Y(_897__bF_buf2) );
BUFX4 BUFX4_1520 ( .gnd(gnd), .vdd(vdd), .A(_897_), .Y(_897__bF_buf1) );
BUFX4 BUFX4_1521 ( .gnd(gnd), .vdd(vdd), .A(_897_), .Y(_897__bF_buf0) );
BUFX4 BUFX4_1522 ( .gnd(gnd), .vdd(vdd), .A(_5073_), .Y(_5073__bF_buf3) );
BUFX4 BUFX4_1523 ( .gnd(gnd), .vdd(vdd), .A(_5073_), .Y(_5073__bF_buf2) );
BUFX4 BUFX4_1524 ( .gnd(gnd), .vdd(vdd), .A(_5073_), .Y(_5073__bF_buf1) );
BUFX4 BUFX4_1525 ( .gnd(gnd), .vdd(vdd), .A(_5073_), .Y(_5073__bF_buf0) );
BUFX4 BUFX4_1526 ( .gnd(gnd), .vdd(vdd), .A(_9285_), .Y(_9285__bF_buf3) );
BUFX4 BUFX4_1527 ( .gnd(gnd), .vdd(vdd), .A(_9285_), .Y(_9285__bF_buf2) );
BUFX4 BUFX4_1528 ( .gnd(gnd), .vdd(vdd), .A(_9285_), .Y(_9285__bF_buf1) );
BUFX4 BUFX4_1529 ( .gnd(gnd), .vdd(vdd), .A(_9285_), .Y(_9285__bF_buf0) );
BUFX4 BUFX4_1530 ( .gnd(gnd), .vdd(vdd), .A(_915_), .Y(_915__bF_buf3) );
BUFX4 BUFX4_1531 ( .gnd(gnd), .vdd(vdd), .A(_915_), .Y(_915__bF_buf2) );
BUFX4 BUFX4_1532 ( .gnd(gnd), .vdd(vdd), .A(_915_), .Y(_915__bF_buf1) );
BUFX4 BUFX4_1533 ( .gnd(gnd), .vdd(vdd), .A(_915_), .Y(_915__bF_buf0) );
BUFX4 BUFX4_1534 ( .gnd(gnd), .vdd(vdd), .A(_8688_), .Y(_8688__bF_buf3) );
BUFX4 BUFX4_1535 ( .gnd(gnd), .vdd(vdd), .A(_8688_), .Y(_8688__bF_buf2) );
BUFX4 BUFX4_1536 ( .gnd(gnd), .vdd(vdd), .A(_8688_), .Y(_8688__bF_buf1) );
BUFX4 BUFX4_1537 ( .gnd(gnd), .vdd(vdd), .A(_8688_), .Y(_8688__bF_buf0) );
BUFX4 BUFX4_1538 ( .gnd(gnd), .vdd(vdd), .A(_11537_), .Y(_11537__bF_buf4) );
BUFX4 BUFX4_1539 ( .gnd(gnd), .vdd(vdd), .A(_11537_), .Y(_11537__bF_buf3) );
BUFX4 BUFX4_1540 ( .gnd(gnd), .vdd(vdd), .A(_11537_), .Y(_11537__bF_buf2) );
BUFX4 BUFX4_1541 ( .gnd(gnd), .vdd(vdd), .A(_11537_), .Y(_11537__bF_buf1) );
BUFX4 BUFX4_1542 ( .gnd(gnd), .vdd(vdd), .A(_11537_), .Y(_11537__bF_buf0) );
BUFX4 BUFX4_1543 ( .gnd(gnd), .vdd(vdd), .A(_894_), .Y(_894__bF_buf3) );
BUFX4 BUFX4_1544 ( .gnd(gnd), .vdd(vdd), .A(_894_), .Y(_894__bF_buf2) );
BUFX4 BUFX4_1545 ( .gnd(gnd), .vdd(vdd), .A(_894_), .Y(_894__bF_buf1) );
BUFX4 BUFX4_1546 ( .gnd(gnd), .vdd(vdd), .A(_894_), .Y(_894__bF_buf0) );
BUFX4 BUFX4_1547 ( .gnd(gnd), .vdd(vdd), .A(_474_), .Y(_474__bF_buf3) );
BUFX4 BUFX4_1548 ( .gnd(gnd), .vdd(vdd), .A(_474_), .Y(_474__bF_buf2) );
BUFX4 BUFX4_1549 ( .gnd(gnd), .vdd(vdd), .A(_474_), .Y(_474__bF_buf1) );
BUFX4 BUFX4_1550 ( .gnd(gnd), .vdd(vdd), .A(_474_), .Y(_474__bF_buf0) );
BUFX4 BUFX4_1551 ( .gnd(gnd), .vdd(vdd), .A(_9282_), .Y(_9282__bF_buf4) );
BUFX4 BUFX4_1552 ( .gnd(gnd), .vdd(vdd), .A(_9282_), .Y(_9282__bF_buf3) );
BUFX4 BUFX4_1553 ( .gnd(gnd), .vdd(vdd), .A(_9282_), .Y(_9282__bF_buf2) );
BUFX4 BUFX4_1554 ( .gnd(gnd), .vdd(vdd), .A(_9282_), .Y(_9282__bF_buf1) );
BUFX4 BUFX4_1555 ( .gnd(gnd), .vdd(vdd), .A(_9282_), .Y(_9282__bF_buf0) );
BUFX4 BUFX4_1556 ( .gnd(gnd), .vdd(vdd), .A(_912_), .Y(_912__bF_buf4) );
BUFX4 BUFX4_1557 ( .gnd(gnd), .vdd(vdd), .A(_912_), .Y(_912__bF_buf3) );
BUFX4 BUFX4_1558 ( .gnd(gnd), .vdd(vdd), .A(_912_), .Y(_912__bF_buf2) );
BUFX4 BUFX4_1559 ( .gnd(gnd), .vdd(vdd), .A(_912_), .Y(_912__bF_buf1) );
BUFX4 BUFX4_1560 ( .gnd(gnd), .vdd(vdd), .A(_912_), .Y(_912__bF_buf0) );
BUFX4 BUFX4_1561 ( .gnd(gnd), .vdd(vdd), .A(_1178_), .Y(_1178__bF_buf3) );
BUFX4 BUFX4_1562 ( .gnd(gnd), .vdd(vdd), .A(_1178_), .Y(_1178__bF_buf2) );
BUFX4 BUFX4_1563 ( .gnd(gnd), .vdd(vdd), .A(_1178_), .Y(_1178__bF_buf1) );
BUFX4 BUFX4_1564 ( .gnd(gnd), .vdd(vdd), .A(_1178_), .Y(_1178__bF_buf0) );
BUFX4 BUFX4_1565 ( .gnd(gnd), .vdd(vdd), .A(_5487_), .Y(_5487__bF_buf3) );
BUFX4 BUFX4_1566 ( .gnd(gnd), .vdd(vdd), .A(_5487_), .Y(_5487__bF_buf2) );
BUFX4 BUFX4_1567 ( .gnd(gnd), .vdd(vdd), .A(_5487_), .Y(_5487__bF_buf1) );
BUFX4 BUFX4_1568 ( .gnd(gnd), .vdd(vdd), .A(_5487_), .Y(_5487__bF_buf0) );
BUFX4 BUFX4_1569 ( .gnd(gnd), .vdd(vdd), .A(_11534_), .Y(_11534__bF_buf3) );
BUFX4 BUFX4_1570 ( .gnd(gnd), .vdd(vdd), .A(_11534_), .Y(_11534__bF_buf2) );
BUFX4 BUFX4_1571 ( .gnd(gnd), .vdd(vdd), .A(_11534_), .Y(_11534__bF_buf1) );
BUFX4 BUFX4_1572 ( .gnd(gnd), .vdd(vdd), .A(_11534_), .Y(_11534__bF_buf0) );
BUFX4 BUFX4_1573 ( .gnd(gnd), .vdd(vdd), .A(_909_), .Y(_909__bF_buf3) );
BUFX4 BUFX4_1574 ( .gnd(gnd), .vdd(vdd), .A(_909_), .Y(_909__bF_buf2) );
BUFX4 BUFX4_1575 ( .gnd(gnd), .vdd(vdd), .A(_909_), .Y(_909__bF_buf1) );
BUFX4 BUFX4_1576 ( .gnd(gnd), .vdd(vdd), .A(_909_), .Y(_909__bF_buf0) );
BUFX4 BUFX4_1577 ( .gnd(gnd), .vdd(vdd), .A(_9300_), .Y(_9300__bF_buf3) );
BUFX4 BUFX4_1578 ( .gnd(gnd), .vdd(vdd), .A(_9300_), .Y(_9300__bF_buf2) );
BUFX4 BUFX4_1579 ( .gnd(gnd), .vdd(vdd), .A(_9300_), .Y(_9300__bF_buf1) );
BUFX4 BUFX4_1580 ( .gnd(gnd), .vdd(vdd), .A(_9300_), .Y(_9300__bF_buf0) );
BUFX4 BUFX4_1581 ( .gnd(gnd), .vdd(vdd), .A(_2574_), .Y(_2574__bF_buf4) );
BUFX4 BUFX4_1582 ( .gnd(gnd), .vdd(vdd), .A(_2574_), .Y(_2574__bF_buf3) );
BUFX4 BUFX4_1583 ( .gnd(gnd), .vdd(vdd), .A(_2574_), .Y(_2574__bF_buf2) );
BUFX4 BUFX4_1584 ( .gnd(gnd), .vdd(vdd), .A(_2574_), .Y(_2574__bF_buf1) );
BUFX4 BUFX4_1585 ( .gnd(gnd), .vdd(vdd), .A(_2574_), .Y(_2574__bF_buf0) );
BUFX4 BUFX4_1586 ( .gnd(gnd), .vdd(vdd), .A(_8800_), .Y(_8800__bF_buf12) );
BUFX4 BUFX4_1587 ( .gnd(gnd), .vdd(vdd), .A(_8800_), .Y(_8800__bF_buf11) );
BUFX4 BUFX4_1588 ( .gnd(gnd), .vdd(vdd), .A(_8800_), .Y(_8800__bF_buf10) );
BUFX4 BUFX4_1589 ( .gnd(gnd), .vdd(vdd), .A(_8800_), .Y(_8800__bF_buf9) );
BUFX4 BUFX4_1590 ( .gnd(gnd), .vdd(vdd), .A(_8800_), .Y(_8800__bF_buf8) );
BUFX4 BUFX4_1591 ( .gnd(gnd), .vdd(vdd), .A(_8800_), .Y(_8800__bF_buf7) );
BUFX4 BUFX4_1592 ( .gnd(gnd), .vdd(vdd), .A(_8800_), .Y(_8800__bF_buf6) );
BUFX4 BUFX4_1593 ( .gnd(gnd), .vdd(vdd), .A(_8800_), .Y(_8800__bF_buf5) );
BUFX4 BUFX4_1594 ( .gnd(gnd), .vdd(vdd), .A(_8800_), .Y(_8800__bF_buf4) );
BUFX4 BUFX4_1595 ( .gnd(gnd), .vdd(vdd), .A(_8800_), .Y(_8800__bF_buf3) );
BUFX4 BUFX4_1596 ( .gnd(gnd), .vdd(vdd), .A(_8800_), .Y(_8800__bF_buf2) );
BUFX4 BUFX4_1597 ( .gnd(gnd), .vdd(vdd), .A(_8800_), .Y(_8800__bF_buf1) );
BUFX4 BUFX4_1598 ( .gnd(gnd), .vdd(vdd), .A(_8800_), .Y(_8800__bF_buf0) );
BUFX4 BUFX4_1599 ( .gnd(gnd), .vdd(vdd), .A(_5123_), .Y(_5123__bF_buf4) );
BUFX4 BUFX4_1600 ( .gnd(gnd), .vdd(vdd), .A(_5123_), .Y(_5123__bF_buf3) );
BUFX4 BUFX4_1601 ( .gnd(gnd), .vdd(vdd), .A(_5123_), .Y(_5123__bF_buf2) );
BUFX4 BUFX4_1602 ( .gnd(gnd), .vdd(vdd), .A(_5123_), .Y(_5123__bF_buf1) );
BUFX4 BUFX4_1603 ( .gnd(gnd), .vdd(vdd), .A(_5123_), .Y(_5123__bF_buf0) );
BUFX4 BUFX4_1604 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe60), .Y(micro_hash_ucr_2_pipe60_bF_buf4) );
BUFX4 BUFX4_1605 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe60), .Y(micro_hash_ucr_2_pipe60_bF_buf3) );
BUFX4 BUFX4_1606 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe60), .Y(micro_hash_ucr_2_pipe60_bF_buf2) );
BUFX4 BUFX4_1607 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe60), .Y(micro_hash_ucr_2_pipe60_bF_buf1) );
BUFX4 BUFX4_1608 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe60), .Y(micro_hash_ucr_2_pipe60_bF_buf0) );
BUFX4 BUFX4_1609 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe61), .Y(micro_hash_ucr_2_pipe61_bF_buf3) );
BUFX4 BUFX4_1610 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe61), .Y(micro_hash_ucr_2_pipe61_bF_buf2) );
BUFX4 BUFX4_1611 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe61), .Y(micro_hash_ucr_2_pipe61_bF_buf1) );
BUFX4 BUFX4_1612 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe61), .Y(micro_hash_ucr_2_pipe61_bF_buf0) );
BUFX4 BUFX4_1613 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe62), .Y(micro_hash_ucr_2_pipe62_bF_buf4) );
BUFX4 BUFX4_1614 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe62), .Y(micro_hash_ucr_2_pipe62_bF_buf3) );
BUFX4 BUFX4_1615 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe62), .Y(micro_hash_ucr_2_pipe62_bF_buf2) );
BUFX4 BUFX4_1616 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe62), .Y(micro_hash_ucr_2_pipe62_bF_buf1) );
BUFX4 BUFX4_1617 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe62), .Y(micro_hash_ucr_2_pipe62_bF_buf0) );
BUFX4 BUFX4_1618 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe64), .Y(micro_hash_ucr_2_pipe64_bF_buf4) );
BUFX4 BUFX4_1619 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe64), .Y(micro_hash_ucr_2_pipe64_bF_buf3) );
BUFX4 BUFX4_1620 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe64), .Y(micro_hash_ucr_2_pipe64_bF_buf2) );
BUFX4 BUFX4_1621 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe64), .Y(micro_hash_ucr_2_pipe64_bF_buf1) );
BUFX4 BUFX4_1622 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe64), .Y(micro_hash_ucr_2_pipe64_bF_buf0) );
BUFX4 BUFX4_1623 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe65), .Y(micro_hash_ucr_2_pipe65_bF_buf3) );
BUFX4 BUFX4_1624 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe65), .Y(micro_hash_ucr_2_pipe65_bF_buf2) );
BUFX4 BUFX4_1625 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe65), .Y(micro_hash_ucr_2_pipe65_bF_buf1) );
BUFX4 BUFX4_1626 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe65), .Y(micro_hash_ucr_2_pipe65_bF_buf0) );
BUFX4 BUFX4_1627 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe66), .Y(micro_hash_ucr_2_pipe66_bF_buf4) );
BUFX4 BUFX4_1628 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe66), .Y(micro_hash_ucr_2_pipe66_bF_buf3) );
BUFX4 BUFX4_1629 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe66), .Y(micro_hash_ucr_2_pipe66_bF_buf2) );
BUFX4 BUFX4_1630 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe66), .Y(micro_hash_ucr_2_pipe66_bF_buf1) );
BUFX4 BUFX4_1631 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe66), .Y(micro_hash_ucr_2_pipe66_bF_buf0) );
BUFX4 BUFX4_1632 ( .gnd(gnd), .vdd(vdd), .A(comparador_3_valid), .Y(comparador_3_valid_bF_buf4) );
BUFX4 BUFX4_1633 ( .gnd(gnd), .vdd(vdd), .A(comparador_3_valid), .Y(comparador_3_valid_bF_buf3) );
BUFX4 BUFX4_1634 ( .gnd(gnd), .vdd(vdd), .A(comparador_3_valid), .Y(comparador_3_valid_bF_buf2) );
BUFX4 BUFX4_1635 ( .gnd(gnd), .vdd(vdd), .A(comparador_3_valid), .Y(comparador_3_valid_bF_buf1) );
BUFX4 BUFX4_1636 ( .gnd(gnd), .vdd(vdd), .A(comparador_3_valid), .Y(comparador_3_valid_bF_buf0) );
BUFX4 BUFX4_1637 ( .gnd(gnd), .vdd(vdd), .A(_888_), .Y(_888__bF_buf3) );
BUFX4 BUFX4_1638 ( .gnd(gnd), .vdd(vdd), .A(_888_), .Y(_888__bF_buf2) );
BUFX4 BUFX4_1639 ( .gnd(gnd), .vdd(vdd), .A(_888_), .Y(_888__bF_buf1) );
BUFX4 BUFX4_1640 ( .gnd(gnd), .vdd(vdd), .A(_888_), .Y(_888__bF_buf0) );
BUFX4 BUFX4_1641 ( .gnd(gnd), .vdd(vdd), .A(_9335_), .Y(_9335__bF_buf3) );
BUFX4 BUFX4_1642 ( .gnd(gnd), .vdd(vdd), .A(_9335_), .Y(_9335__bF_buf2) );
BUFX4 BUFX4_1643 ( .gnd(gnd), .vdd(vdd), .A(_9335_), .Y(_9335__bF_buf1) );
BUFX4 BUFX4_1644 ( .gnd(gnd), .vdd(vdd), .A(_9335_), .Y(_9335__bF_buf0) );
BUFX4 BUFX4_1645 ( .gnd(gnd), .vdd(vdd), .A(_13618_), .Y(_13618__bF_buf4) );
BUFX4 BUFX4_1646 ( .gnd(gnd), .vdd(vdd), .A(_13618_), .Y(_13618__bF_buf3) );
BUFX4 BUFX4_1647 ( .gnd(gnd), .vdd(vdd), .A(_13618_), .Y(_13618__bF_buf2) );
BUFX4 BUFX4_1648 ( .gnd(gnd), .vdd(vdd), .A(_13618_), .Y(_13618__bF_buf1) );
BUFX4 BUFX4_1649 ( .gnd(gnd), .vdd(vdd), .A(_13618_), .Y(_13618__bF_buf0) );
BUFX4 BUFX4_1650 ( .gnd(gnd), .vdd(vdd), .A(_2304_), .Y(_2304__bF_buf3) );
BUFX4 BUFX4_1651 ( .gnd(gnd), .vdd(vdd), .A(_2304_), .Y(_2304__bF_buf2) );
BUFX4 BUFX4_1652 ( .gnd(gnd), .vdd(vdd), .A(_2304_), .Y(_2304__bF_buf1) );
BUFX4 BUFX4_1653 ( .gnd(gnd), .vdd(vdd), .A(_2304_), .Y(_2304__bF_buf0) );
BUFX4 BUFX4_1654 ( .gnd(gnd), .vdd(vdd), .A(_906_), .Y(_906__bF_buf4) );
BUFX4 BUFX4_1655 ( .gnd(gnd), .vdd(vdd), .A(_906_), .Y(_906__bF_buf3) );
BUFX4 BUFX4_1656 ( .gnd(gnd), .vdd(vdd), .A(_906_), .Y(_906__bF_buf2) );
BUFX4 BUFX4_1657 ( .gnd(gnd), .vdd(vdd), .A(_906_), .Y(_906__bF_buf1) );
BUFX4 BUFX4_1658 ( .gnd(gnd), .vdd(vdd), .A(_906_), .Y(_906__bF_buf0) );
BUFX4 BUFX4_1659 ( .gnd(gnd), .vdd(vdd), .A(_944_), .Y(_944__bF_buf3) );
BUFX4 BUFX4_1660 ( .gnd(gnd), .vdd(vdd), .A(_944_), .Y(_944__bF_buf2) );
BUFX4 BUFX4_1661 ( .gnd(gnd), .vdd(vdd), .A(_944_), .Y(_944__bF_buf1) );
BUFX4 BUFX4_1662 ( .gnd(gnd), .vdd(vdd), .A(_944_), .Y(_944__bF_buf0) );
BUFX4 BUFX4_1663 ( .gnd(gnd), .vdd(vdd), .A(_5099_), .Y(_5099__bF_buf4) );
BUFX4 BUFX4_1664 ( .gnd(gnd), .vdd(vdd), .A(_5099_), .Y(_5099__bF_buf3) );
BUFX4 BUFX4_1665 ( .gnd(gnd), .vdd(vdd), .A(_5099_), .Y(_5099__bF_buf2) );
BUFX4 BUFX4_1666 ( .gnd(gnd), .vdd(vdd), .A(_5099_), .Y(_5099__bF_buf1) );
BUFX4 BUFX4_1667 ( .gnd(gnd), .vdd(vdd), .A(_5099_), .Y(_5099__bF_buf0) );
BUFX4 BUFX4_1668 ( .gnd(gnd), .vdd(vdd), .A(_5120_), .Y(_5120__bF_buf3) );
BUFX4 BUFX4_1669 ( .gnd(gnd), .vdd(vdd), .A(_5120_), .Y(_5120__bF_buf2) );
BUFX4 BUFX4_1670 ( .gnd(gnd), .vdd(vdd), .A(_5120_), .Y(_5120__bF_buf1) );
BUFX4 BUFX4_1671 ( .gnd(gnd), .vdd(vdd), .A(_5120_), .Y(_5120__bF_buf0) );
BUFX4 BUFX4_1672 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe30), .Y(micro_hash_ucr_2_pipe30_bF_buf4) );
BUFX4 BUFX4_1673 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe30), .Y(micro_hash_ucr_2_pipe30_bF_buf3) );
BUFX4 BUFX4_1674 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe30), .Y(micro_hash_ucr_2_pipe30_bF_buf2) );
BUFX4 BUFX4_1675 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe30), .Y(micro_hash_ucr_2_pipe30_bF_buf1) );
BUFX4 BUFX4_1676 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe30), .Y(micro_hash_ucr_2_pipe30_bF_buf0) );
BUFX4 BUFX4_1677 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe32), .Y(micro_hash_ucr_2_pipe32_bF_buf3) );
BUFX4 BUFX4_1678 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe32), .Y(micro_hash_ucr_2_pipe32_bF_buf2) );
BUFX4 BUFX4_1679 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe32), .Y(micro_hash_ucr_2_pipe32_bF_buf1) );
BUFX4 BUFX4_1680 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe32), .Y(micro_hash_ucr_2_pipe32_bF_buf0) );
BUFX4 BUFX4_1681 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe33), .Y(micro_hash_ucr_2_pipe33_bF_buf3) );
BUFX4 BUFX4_1682 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe33), .Y(micro_hash_ucr_2_pipe33_bF_buf2) );
BUFX4 BUFX4_1683 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe33), .Y(micro_hash_ucr_2_pipe33_bF_buf1) );
BUFX4 BUFX4_1684 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe33), .Y(micro_hash_ucr_2_pipe33_bF_buf0) );
BUFX4 BUFX4_1685 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe34), .Y(micro_hash_ucr_2_pipe34_bF_buf3) );
BUFX4 BUFX4_1686 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe34), .Y(micro_hash_ucr_2_pipe34_bF_buf2) );
BUFX4 BUFX4_1687 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe34), .Y(micro_hash_ucr_2_pipe34_bF_buf1) );
BUFX4 BUFX4_1688 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe34), .Y(micro_hash_ucr_2_pipe34_bF_buf0) );
BUFX4 BUFX4_1689 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe36), .Y(micro_hash_ucr_2_pipe36_bF_buf3) );
BUFX4 BUFX4_1690 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe36), .Y(micro_hash_ucr_2_pipe36_bF_buf2) );
BUFX4 BUFX4_1691 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe36), .Y(micro_hash_ucr_2_pipe36_bF_buf1) );
BUFX4 BUFX4_1692 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe36), .Y(micro_hash_ucr_2_pipe36_bF_buf0) );
BUFX4 BUFX4_1693 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe38), .Y(micro_hash_ucr_2_pipe38_bF_buf3) );
BUFX4 BUFX4_1694 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe38), .Y(micro_hash_ucr_2_pipe38_bF_buf2) );
BUFX4 BUFX4_1695 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe38), .Y(micro_hash_ucr_2_pipe38_bF_buf1) );
BUFX4 BUFX4_1696 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe38), .Y(micro_hash_ucr_2_pipe38_bF_buf0) );
BUFX4 BUFX4_1697 ( .gnd(gnd), .vdd(vdd), .A(_13615_), .Y(_13615__bF_buf4) );
BUFX4 BUFX4_1698 ( .gnd(gnd), .vdd(vdd), .A(_13615_), .Y(_13615__bF_buf3) );
BUFX4 BUFX4_1699 ( .gnd(gnd), .vdd(vdd), .A(_13615_), .Y(_13615__bF_buf2) );
BUFX4 BUFX4_1700 ( .gnd(gnd), .vdd(vdd), .A(_13615_), .Y(_13615__bF_buf1) );
BUFX4 BUFX4_1701 ( .gnd(gnd), .vdd(vdd), .A(_13615_), .Y(_13615__bF_buf0) );
BUFX4 BUFX4_1702 ( .gnd(gnd), .vdd(vdd), .A(_5117_), .Y(_5117__bF_buf4) );
BUFX4 BUFX4_1703 ( .gnd(gnd), .vdd(vdd), .A(_5117_), .Y(_5117__bF_buf3) );
BUFX4 BUFX4_1704 ( .gnd(gnd), .vdd(vdd), .A(_5117_), .Y(_5117__bF_buf2) );
BUFX4 BUFX4_1705 ( .gnd(gnd), .vdd(vdd), .A(_5117_), .Y(_5117__bF_buf1) );
BUFX4 BUFX4_1706 ( .gnd(gnd), .vdd(vdd), .A(_5117_), .Y(_5117__bF_buf0) );
BUFX4 BUFX4_1707 ( .gnd(gnd), .vdd(vdd), .A(_7301_), .Y(_7301__bF_buf3) );
BUFX4 BUFX4_1708 ( .gnd(gnd), .vdd(vdd), .A(_7301_), .Y(_7301__bF_buf2) );
BUFX4 BUFX4_1709 ( .gnd(gnd), .vdd(vdd), .A(_7301_), .Y(_7301__bF_buf1) );
BUFX4 BUFX4_1710 ( .gnd(gnd), .vdd(vdd), .A(_7301_), .Y(_7301__bF_buf0) );
BUFX4 BUFX4_1711 ( .gnd(gnd), .vdd(vdd), .A(_2089_), .Y(_2089__bF_buf5) );
BUFX4 BUFX4_1712 ( .gnd(gnd), .vdd(vdd), .A(_2089_), .Y(_2089__bF_buf4) );
BUFX4 BUFX4_1713 ( .gnd(gnd), .vdd(vdd), .A(_2089_), .Y(_2089__bF_buf3) );
BUFX4 BUFX4_1714 ( .gnd(gnd), .vdd(vdd), .A(_2089_), .Y(_2089__bF_buf2) );
BUFX4 BUFX4_1715 ( .gnd(gnd), .vdd(vdd), .A(_2089_), .Y(_2089__bF_buf1) );
BUFX4 BUFX4_1716 ( .gnd(gnd), .vdd(vdd), .A(_2089_), .Y(_2089__bF_buf0) );
BUFX4 BUFX4_1717 ( .gnd(gnd), .vdd(vdd), .A(_9329_), .Y(_9329__bF_buf4) );
BUFX4 BUFX4_1718 ( .gnd(gnd), .vdd(vdd), .A(_9329_), .Y(_9329__bF_buf3) );
BUFX4 BUFX4_1719 ( .gnd(gnd), .vdd(vdd), .A(_9329_), .Y(_9329__bF_buf2) );
BUFX4 BUFX4_1720 ( .gnd(gnd), .vdd(vdd), .A(_9329_), .Y(_9329__bF_buf1) );
BUFX4 BUFX4_1721 ( .gnd(gnd), .vdd(vdd), .A(_9329_), .Y(_9329__bF_buf0) );
BUFX4 BUFX4_1722 ( .gnd(gnd), .vdd(vdd), .A(_903_), .Y(_903__bF_buf3) );
BUFX4 BUFX4_1723 ( .gnd(gnd), .vdd(vdd), .A(_903_), .Y(_903__bF_buf2) );
BUFX4 BUFX4_1724 ( .gnd(gnd), .vdd(vdd), .A(_903_), .Y(_903__bF_buf1) );
BUFX4 BUFX4_1725 ( .gnd(gnd), .vdd(vdd), .A(_903_), .Y(_903__bF_buf0) );
BUFX4 BUFX4_1726 ( .gnd(gnd), .vdd(vdd), .A(_5096_), .Y(_5096__bF_buf3) );
BUFX4 BUFX4_1727 ( .gnd(gnd), .vdd(vdd), .A(_5096_), .Y(_5096__bF_buf2) );
BUFX4 BUFX4_1728 ( .gnd(gnd), .vdd(vdd), .A(_5096_), .Y(_5096__bF_buf1) );
BUFX4 BUFX4_1729 ( .gnd(gnd), .vdd(vdd), .A(_5096_), .Y(_5096__bF_buf0) );
BUFX4 BUFX4_1730 ( .gnd(gnd), .vdd(vdd), .A(_882_), .Y(_882__bF_buf3) );
BUFX4 BUFX4_1731 ( .gnd(gnd), .vdd(vdd), .A(_882_), .Y(_882__bF_buf2) );
BUFX4 BUFX4_1732 ( .gnd(gnd), .vdd(vdd), .A(_882_), .Y(_882__bF_buf1) );
BUFX4 BUFX4_1733 ( .gnd(gnd), .vdd(vdd), .A(_882_), .Y(_882__bF_buf0) );
BUFX4 BUFX4_1734 ( .gnd(gnd), .vdd(vdd), .A(_11008_), .Y(_11008__bF_buf4) );
BUFX4 BUFX4_1735 ( .gnd(gnd), .vdd(vdd), .A(_11008_), .Y(_11008__bF_buf3) );
BUFX4 BUFX4_1736 ( .gnd(gnd), .vdd(vdd), .A(_11008_), .Y(_11008__bF_buf2) );
BUFX4 BUFX4_1737 ( .gnd(gnd), .vdd(vdd), .A(_11008_), .Y(_11008__bF_buf1) );
BUFX4 BUFX4_1738 ( .gnd(gnd), .vdd(vdd), .A(_11008_), .Y(_11008__bF_buf0) );
BUFX4 BUFX4_1739 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_2_), .Y(micro_hash_ucr_2_c_2_bF_buf3_) );
BUFX4 BUFX4_1740 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_2_), .Y(micro_hash_ucr_2_c_2_bF_buf2_) );
BUFX4 BUFX4_1741 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_2_), .Y(micro_hash_ucr_2_c_2_bF_buf1_) );
BUFX4 BUFX4_1742 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_2_), .Y(micro_hash_ucr_2_c_2_bF_buf0_) );
BUFX4 BUFX4_1743 ( .gnd(gnd), .vdd(vdd), .A(_10737_), .Y(_10737__bF_buf3) );
BUFX4 BUFX4_1744 ( .gnd(gnd), .vdd(vdd), .A(_10737_), .Y(_10737__bF_buf2) );
BUFX4 BUFX4_1745 ( .gnd(gnd), .vdd(vdd), .A(_10737_), .Y(_10737__bF_buf1) );
BUFX4 BUFX4_1746 ( .gnd(gnd), .vdd(vdd), .A(_10737_), .Y(_10737__bF_buf0) );
BUFX4 BUFX4_1747 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_5_), .Y(micro_hash_ucr_2_b_5_bF_buf3_) );
BUFX4 BUFX4_1748 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_5_), .Y(micro_hash_ucr_2_b_5_bF_buf2_) );
BUFX4 BUFX4_1749 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_5_), .Y(micro_hash_ucr_2_b_5_bF_buf1_) );
BUFX4 BUFX4_1750 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_5_), .Y(micro_hash_ucr_2_b_5_bF_buf0_) );
BUFX4 BUFX4_1751 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_3_), .Y(micro_hash_ucr_3_c_3_bF_buf3_) );
BUFX4 BUFX4_1752 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_3_), .Y(micro_hash_ucr_3_c_3_bF_buf2_) );
BUFX4 BUFX4_1753 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_3_), .Y(micro_hash_ucr_3_c_3_bF_buf1_) );
BUFX4 BUFX4_1754 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_3_), .Y(micro_hash_ucr_3_c_3_bF_buf0_) );
BUFX4 BUFX4_1755 ( .gnd(gnd), .vdd(vdd), .A(_4423_), .Y(_4423__bF_buf3) );
BUFX4 BUFX4_1756 ( .gnd(gnd), .vdd(vdd), .A(_4423_), .Y(_4423__bF_buf2) );
BUFX4 BUFX4_1757 ( .gnd(gnd), .vdd(vdd), .A(_4423_), .Y(_4423__bF_buf1) );
BUFX4 BUFX4_1758 ( .gnd(gnd), .vdd(vdd), .A(_4423_), .Y(_4423__bF_buf0) );
BUFX4 BUFX4_1759 ( .gnd(gnd), .vdd(vdd), .A(_879_), .Y(_879__bF_buf3) );
BUFX4 BUFX4_1760 ( .gnd(gnd), .vdd(vdd), .A(_879_), .Y(_879__bF_buf2) );
BUFX4 BUFX4_1761 ( .gnd(gnd), .vdd(vdd), .A(_879_), .Y(_879__bF_buf1) );
BUFX4 BUFX4_1762 ( .gnd(gnd), .vdd(vdd), .A(_879_), .Y(_879__bF_buf0) );
BUFX4 BUFX4_1763 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe50), .Y(micro_hash_ucr_3_pipe50_bF_buf4) );
BUFX4 BUFX4_1764 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe50), .Y(micro_hash_ucr_3_pipe50_bF_buf3) );
BUFX4 BUFX4_1765 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe50), .Y(micro_hash_ucr_3_pipe50_bF_buf2) );
BUFX4 BUFX4_1766 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe50), .Y(micro_hash_ucr_3_pipe50_bF_buf1) );
BUFX4 BUFX4_1767 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe50), .Y(micro_hash_ucr_3_pipe50_bF_buf0) );
BUFX4 BUFX4_1768 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe52), .Y(micro_hash_ucr_3_pipe52_bF_buf4) );
BUFX4 BUFX4_1769 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe52), .Y(micro_hash_ucr_3_pipe52_bF_buf3) );
BUFX4 BUFX4_1770 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe52), .Y(micro_hash_ucr_3_pipe52_bF_buf2) );
BUFX4 BUFX4_1771 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe52), .Y(micro_hash_ucr_3_pipe52_bF_buf1) );
BUFX4 BUFX4_1772 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe52), .Y(micro_hash_ucr_3_pipe52_bF_buf0) );
BUFX4 BUFX4_1773 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe54), .Y(micro_hash_ucr_3_pipe54_bF_buf3) );
BUFX4 BUFX4_1774 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe54), .Y(micro_hash_ucr_3_pipe54_bF_buf2) );
BUFX4 BUFX4_1775 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe54), .Y(micro_hash_ucr_3_pipe54_bF_buf1) );
BUFX4 BUFX4_1776 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe54), .Y(micro_hash_ucr_3_pipe54_bF_buf0) );
BUFX4 BUFX4_1777 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe56), .Y(micro_hash_ucr_3_pipe56_bF_buf4) );
BUFX4 BUFX4_1778 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe56), .Y(micro_hash_ucr_3_pipe56_bF_buf3) );
BUFX4 BUFX4_1779 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe56), .Y(micro_hash_ucr_3_pipe56_bF_buf2) );
BUFX4 BUFX4_1780 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe56), .Y(micro_hash_ucr_3_pipe56_bF_buf1) );
BUFX4 BUFX4_1781 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe56), .Y(micro_hash_ucr_3_pipe56_bF_buf0) );
BUFX4 BUFX4_1782 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe57), .Y(micro_hash_ucr_3_pipe57_bF_buf3) );
BUFX4 BUFX4_1783 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe57), .Y(micro_hash_ucr_3_pipe57_bF_buf2) );
BUFX4 BUFX4_1784 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe57), .Y(micro_hash_ucr_3_pipe57_bF_buf1) );
BUFX4 BUFX4_1785 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe57), .Y(micro_hash_ucr_3_pipe57_bF_buf0) );
BUFX4 BUFX4_1786 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe58), .Y(micro_hash_ucr_3_pipe58_bF_buf3) );
BUFX4 BUFX4_1787 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe58), .Y(micro_hash_ucr_3_pipe58_bF_buf2) );
BUFX4 BUFX4_1788 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe58), .Y(micro_hash_ucr_3_pipe58_bF_buf1) );
BUFX4 BUFX4_1789 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe58), .Y(micro_hash_ucr_3_pipe58_bF_buf0) );
BUFX4 BUFX4_1790 ( .gnd(gnd), .vdd(vdd), .A(_9326_), .Y(_9326__bF_buf3) );
BUFX4 BUFX4_1791 ( .gnd(gnd), .vdd(vdd), .A(_9326_), .Y(_9326__bF_buf2) );
BUFX4 BUFX4_1792 ( .gnd(gnd), .vdd(vdd), .A(_9326_), .Y(_9326__bF_buf1) );
BUFX4 BUFX4_1793 ( .gnd(gnd), .vdd(vdd), .A(_9326_), .Y(_9326__bF_buf0) );
BUFX4 BUFX4_1794 ( .gnd(gnd), .vdd(vdd), .A(_900_), .Y(_900__bF_buf3) );
BUFX4 BUFX4_1795 ( .gnd(gnd), .vdd(vdd), .A(_900_), .Y(_900__bF_buf2) );
BUFX4 BUFX4_1796 ( .gnd(gnd), .vdd(vdd), .A(_900_), .Y(_900__bF_buf1) );
BUFX4 BUFX4_1797 ( .gnd(gnd), .vdd(vdd), .A(_900_), .Y(_900__bF_buf0) );
BUFX4 BUFX4_1798 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_6_), .Y(micro_hash_ucr_3_b_6_bF_buf3_) );
BUFX4 BUFX4_1799 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_6_), .Y(micro_hash_ucr_3_b_6_bF_buf2_) );
BUFX4 BUFX4_1800 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_6_), .Y(micro_hash_ucr_3_b_6_bF_buf1_) );
BUFX4 BUFX4_1801 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_6_), .Y(micro_hash_ucr_3_b_6_bF_buf0_) );
BUFX4 BUFX4_1802 ( .gnd(gnd), .vdd(vdd), .A(_9593_), .Y(_9593__bF_buf3) );
BUFX4 BUFX4_1803 ( .gnd(gnd), .vdd(vdd), .A(_9593_), .Y(_9593__bF_buf2) );
BUFX4 BUFX4_1804 ( .gnd(gnd), .vdd(vdd), .A(_9593_), .Y(_9593__bF_buf1) );
BUFX4 BUFX4_1805 ( .gnd(gnd), .vdd(vdd), .A(_9593_), .Y(_9593__bF_buf0) );
BUFX4 BUFX4_1806 ( .gnd(gnd), .vdd(vdd), .A(_5093_), .Y(_5093__bF_buf4) );
BUFX4 BUFX4_1807 ( .gnd(gnd), .vdd(vdd), .A(_5093_), .Y(_5093__bF_buf3) );
BUFX4 BUFX4_1808 ( .gnd(gnd), .vdd(vdd), .A(_5093_), .Y(_5093__bF_buf2) );
BUFX4 BUFX4_1809 ( .gnd(gnd), .vdd(vdd), .A(_5093_), .Y(_5093__bF_buf1) );
BUFX4 BUFX4_1810 ( .gnd(gnd), .vdd(vdd), .A(_5093_), .Y(_5093__bF_buf0) );
BUFX4 BUFX4_1811 ( .gnd(gnd), .vdd(vdd), .A(reset), .Y(reset_bF_buf10) );
BUFX4 BUFX4_1812 ( .gnd(gnd), .vdd(vdd), .A(reset), .Y(reset_bF_buf9) );
BUFX4 BUFX4_1813 ( .gnd(gnd), .vdd(vdd), .A(reset), .Y(reset_bF_buf8) );
BUFX4 BUFX4_1814 ( .gnd(gnd), .vdd(vdd), .A(reset), .Y(reset_bF_buf7) );
BUFX4 BUFX4_1815 ( .gnd(gnd), .vdd(vdd), .A(reset), .Y(reset_bF_buf6) );
BUFX4 BUFX4_1816 ( .gnd(gnd), .vdd(vdd), .A(reset), .Y(reset_bF_buf5) );
BUFX4 BUFX4_1817 ( .gnd(gnd), .vdd(vdd), .A(reset), .Y(reset_bF_buf4) );
BUFX4 BUFX4_1818 ( .gnd(gnd), .vdd(vdd), .A(reset), .Y(reset_bF_buf3) );
BUFX4 BUFX4_1819 ( .gnd(gnd), .vdd(vdd), .A(reset), .Y(reset_bF_buf2) );
BUFX4 BUFX4_1820 ( .gnd(gnd), .vdd(vdd), .A(reset), .Y(reset_bF_buf1) );
BUFX4 BUFX4_1821 ( .gnd(gnd), .vdd(vdd), .A(reset), .Y(reset_bF_buf0) );
BUFX4 BUFX4_1822 ( .gnd(gnd), .vdd(vdd), .A(_7562_), .Y(_7562__bF_buf4) );
BUFX4 BUFX4_1823 ( .gnd(gnd), .vdd(vdd), .A(_7562_), .Y(_7562__bF_buf3) );
BUFX4 BUFX4_1824 ( .gnd(gnd), .vdd(vdd), .A(_7562_), .Y(_7562__bF_buf2) );
BUFX4 BUFX4_1825 ( .gnd(gnd), .vdd(vdd), .A(_7562_), .Y(_7562__bF_buf1) );
BUFX4 BUFX4_1826 ( .gnd(gnd), .vdd(vdd), .A(_7562_), .Y(_7562__bF_buf0) );
BUFX4 BUFX4_1827 ( .gnd(gnd), .vdd(vdd), .A(_11560_), .Y(_11560__bF_buf3) );
BUFX4 BUFX4_1828 ( .gnd(gnd), .vdd(vdd), .A(_11560_), .Y(_11560__bF_buf2) );
BUFX4 BUFX4_1829 ( .gnd(gnd), .vdd(vdd), .A(_11560_), .Y(_11560__bF_buf1) );
BUFX4 BUFX4_1830 ( .gnd(gnd), .vdd(vdd), .A(_11560_), .Y(_11560__bF_buf0) );
BUFX4 BUFX4_1831 ( .gnd(gnd), .vdd(vdd), .A(_4496_), .Y(_4496__bF_buf13) );
BUFX4 BUFX4_1832 ( .gnd(gnd), .vdd(vdd), .A(_4496_), .Y(_4496__bF_buf12) );
BUFX4 BUFX4_1833 ( .gnd(gnd), .vdd(vdd), .A(_4496_), .Y(_4496__bF_buf11) );
BUFX4 BUFX4_1834 ( .gnd(gnd), .vdd(vdd), .A(_4496_), .Y(_4496__bF_buf10) );
BUFX4 BUFX4_1835 ( .gnd(gnd), .vdd(vdd), .A(_4496_), .Y(_4496__bF_buf9) );
BUFX4 BUFX4_1836 ( .gnd(gnd), .vdd(vdd), .A(_4496_), .Y(_4496__bF_buf8) );
BUFX4 BUFX4_1837 ( .gnd(gnd), .vdd(vdd), .A(_4496_), .Y(_4496__bF_buf7) );
BUFX4 BUFX4_1838 ( .gnd(gnd), .vdd(vdd), .A(_4496_), .Y(_4496__bF_buf6) );
BUFX4 BUFX4_1839 ( .gnd(gnd), .vdd(vdd), .A(_4496_), .Y(_4496__bF_buf5) );
BUFX4 BUFX4_1840 ( .gnd(gnd), .vdd(vdd), .A(_4496_), .Y(_4496__bF_buf4) );
BUFX4 BUFX4_1841 ( .gnd(gnd), .vdd(vdd), .A(_4496_), .Y(_4496__bF_buf3) );
BUFX4 BUFX4_1842 ( .gnd(gnd), .vdd(vdd), .A(_4496_), .Y(_4496__bF_buf2) );
BUFX4 BUFX4_1843 ( .gnd(gnd), .vdd(vdd), .A(_4496_), .Y(_4496__bF_buf1) );
BUFX4 BUFX4_1844 ( .gnd(gnd), .vdd(vdd), .A(_4496_), .Y(_4496__bF_buf0) );
BUFX4 BUFX4_1845 ( .gnd(gnd), .vdd(vdd), .A(_3576_), .Y(_3576__bF_buf4) );
BUFX4 BUFX4_1846 ( .gnd(gnd), .vdd(vdd), .A(_3576_), .Y(_3576__bF_buf3) );
BUFX4 BUFX4_1847 ( .gnd(gnd), .vdd(vdd), .A(_3576_), .Y(_3576__bF_buf2) );
BUFX4 BUFX4_1848 ( .gnd(gnd), .vdd(vdd), .A(_3576_), .Y(_3576__bF_buf1) );
BUFX4 BUFX4_1849 ( .gnd(gnd), .vdd(vdd), .A(_3576_), .Y(_3576__bF_buf0) );
BUFX4 BUFX4_1850 ( .gnd(gnd), .vdd(vdd), .A(_5111_), .Y(_5111__bF_buf4) );
BUFX4 BUFX4_1851 ( .gnd(gnd), .vdd(vdd), .A(_5111_), .Y(_5111__bF_buf3) );
BUFX4 BUFX4_1852 ( .gnd(gnd), .vdd(vdd), .A(_5111_), .Y(_5111__bF_buf2) );
BUFX4 BUFX4_1853 ( .gnd(gnd), .vdd(vdd), .A(_5111_), .Y(_5111__bF_buf1) );
BUFX4 BUFX4_1854 ( .gnd(gnd), .vdd(vdd), .A(_5111_), .Y(_5111__bF_buf0) );
BUFX4 BUFX4_1855 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_2_), .Y(micro_hash_ucr_2_b_2_bF_buf3_) );
BUFX4 BUFX4_1856 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_2_), .Y(micro_hash_ucr_2_b_2_bF_buf2_) );
BUFX4 BUFX4_1857 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_2_), .Y(micro_hash_ucr_2_b_2_bF_buf1_) );
BUFX4 BUFX4_1858 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_2_), .Y(micro_hash_ucr_2_b_2_bF_buf0_) );
BUFX4 BUFX4_1859 ( .gnd(gnd), .vdd(vdd), .A(_9705_), .Y(_9705__bF_buf3) );
BUFX4 BUFX4_1860 ( .gnd(gnd), .vdd(vdd), .A(_9705_), .Y(_9705__bF_buf2) );
BUFX4 BUFX4_1861 ( .gnd(gnd), .vdd(vdd), .A(_9705_), .Y(_9705__bF_buf1) );
BUFX4 BUFX4_1862 ( .gnd(gnd), .vdd(vdd), .A(_9705_), .Y(_9705__bF_buf0) );
BUFX4 BUFX4_1863 ( .gnd(gnd), .vdd(vdd), .A(_876_), .Y(_876__bF_buf3) );
BUFX4 BUFX4_1864 ( .gnd(gnd), .vdd(vdd), .A(_876_), .Y(_876__bF_buf2) );
BUFX4 BUFX4_1865 ( .gnd(gnd), .vdd(vdd), .A(_876_), .Y(_876__bF_buf1) );
BUFX4 BUFX4_1866 ( .gnd(gnd), .vdd(vdd), .A(_876_), .Y(_876__bF_buf0) );
BUFX4 BUFX4_1867 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe20), .Y(micro_hash_ucr_3_pipe20_bF_buf4) );
BUFX4 BUFX4_1868 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe20), .Y(micro_hash_ucr_3_pipe20_bF_buf3) );
BUFX4 BUFX4_1869 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe20), .Y(micro_hash_ucr_3_pipe20_bF_buf2) );
BUFX4 BUFX4_1870 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe20), .Y(micro_hash_ucr_3_pipe20_bF_buf1) );
BUFX4 BUFX4_1871 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe20), .Y(micro_hash_ucr_3_pipe20_bF_buf0) );
BUFX4 BUFX4_1872 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe21), .Y(micro_hash_ucr_3_pipe21_bF_buf3) );
BUFX4 BUFX4_1873 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe21), .Y(micro_hash_ucr_3_pipe21_bF_buf2) );
BUFX4 BUFX4_1874 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe21), .Y(micro_hash_ucr_3_pipe21_bF_buf1) );
BUFX4 BUFX4_1875 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe21), .Y(micro_hash_ucr_3_pipe21_bF_buf0) );
BUFX4 BUFX4_1876 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe22), .Y(micro_hash_ucr_3_pipe22_bF_buf4) );
BUFX4 BUFX4_1877 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe22), .Y(micro_hash_ucr_3_pipe22_bF_buf3) );
BUFX4 BUFX4_1878 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe22), .Y(micro_hash_ucr_3_pipe22_bF_buf2) );
BUFX4 BUFX4_1879 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe22), .Y(micro_hash_ucr_3_pipe22_bF_buf1) );
BUFX4 BUFX4_1880 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe22), .Y(micro_hash_ucr_3_pipe22_bF_buf0) );
BUFX4 BUFX4_1881 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe24), .Y(micro_hash_ucr_3_pipe24_bF_buf4) );
BUFX4 BUFX4_1882 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe24), .Y(micro_hash_ucr_3_pipe24_bF_buf3) );
BUFX4 BUFX4_1883 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe24), .Y(micro_hash_ucr_3_pipe24_bF_buf2) );
BUFX4 BUFX4_1884 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe24), .Y(micro_hash_ucr_3_pipe24_bF_buf1) );
BUFX4 BUFX4_1885 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe24), .Y(micro_hash_ucr_3_pipe24_bF_buf0) );
BUFX4 BUFX4_1886 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe25), .Y(micro_hash_ucr_3_pipe25_bF_buf3) );
BUFX4 BUFX4_1887 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe25), .Y(micro_hash_ucr_3_pipe25_bF_buf2) );
BUFX4 BUFX4_1888 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe25), .Y(micro_hash_ucr_3_pipe25_bF_buf1) );
BUFX4 BUFX4_1889 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe25), .Y(micro_hash_ucr_3_pipe25_bF_buf0) );
BUFX4 BUFX4_1890 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe26), .Y(micro_hash_ucr_3_pipe26_bF_buf4) );
BUFX4 BUFX4_1891 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe26), .Y(micro_hash_ucr_3_pipe26_bF_buf3) );
BUFX4 BUFX4_1892 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe26), .Y(micro_hash_ucr_3_pipe26_bF_buf2) );
BUFX4 BUFX4_1893 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe26), .Y(micro_hash_ucr_3_pipe26_bF_buf1) );
BUFX4 BUFX4_1894 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe26), .Y(micro_hash_ucr_3_pipe26_bF_buf0) );
BUFX4 BUFX4_1895 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe28), .Y(micro_hash_ucr_3_pipe28_bF_buf4) );
BUFX4 BUFX4_1896 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe28), .Y(micro_hash_ucr_3_pipe28_bF_buf3) );
BUFX4 BUFX4_1897 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe28), .Y(micro_hash_ucr_3_pipe28_bF_buf2) );
BUFX4 BUFX4_1898 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe28), .Y(micro_hash_ucr_3_pipe28_bF_buf1) );
BUFX4 BUFX4_1899 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe28), .Y(micro_hash_ucr_3_pipe28_bF_buf0) );
BUFX4 BUFX4_1900 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe29), .Y(micro_hash_ucr_3_pipe29_bF_buf3) );
BUFX4 BUFX4_1901 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe29), .Y(micro_hash_ucr_3_pipe29_bF_buf2) );
BUFX4 BUFX4_1902 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe29), .Y(micro_hash_ucr_3_pipe29_bF_buf1) );
BUFX4 BUFX4_1903 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe29), .Y(micro_hash_ucr_3_pipe29_bF_buf0) );
BUFX4 BUFX4_1904 ( .gnd(gnd), .vdd(vdd), .A(_9323_), .Y(_9323__bF_buf3) );
BUFX4 BUFX4_1905 ( .gnd(gnd), .vdd(vdd), .A(_9323_), .Y(_9323__bF_buf2) );
BUFX4 BUFX4_1906 ( .gnd(gnd), .vdd(vdd), .A(_9323_), .Y(_9323__bF_buf1) );
BUFX4 BUFX4_1907 ( .gnd(gnd), .vdd(vdd), .A(_9323_), .Y(_9323__bF_buf0) );
BUFX4 BUFX4_1908 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_5_), .Y(micro_hash_ucr_2_a_5_bF_buf3_) );
BUFX4 BUFX4_1909 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_5_), .Y(micro_hash_ucr_2_a_5_bF_buf2_) );
BUFX4 BUFX4_1910 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_5_), .Y(micro_hash_ucr_2_a_5_bF_buf1_) );
BUFX4 BUFX4_1911 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_5_), .Y(micro_hash_ucr_2_a_5_bF_buf0_) );
BUFX4 BUFX4_1912 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_3_), .Y(micro_hash_ucr_3_b_3_bF_buf3_) );
BUFX4 BUFX4_1913 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_3_), .Y(micro_hash_ucr_3_b_3_bF_buf2_) );
BUFX4 BUFX4_1914 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_3_), .Y(micro_hash_ucr_3_b_3_bF_buf1_) );
BUFX4 BUFX4_1915 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_3_), .Y(micro_hash_ucr_3_b_3_bF_buf0_) );
BUFX4 BUFX4_1916 ( .gnd(gnd), .vdd(vdd), .A(_5108_), .Y(_5108__bF_buf3) );
BUFX4 BUFX4_1917 ( .gnd(gnd), .vdd(vdd), .A(_5108_), .Y(_5108__bF_buf2) );
BUFX4 BUFX4_1918 ( .gnd(gnd), .vdd(vdd), .A(_5108_), .Y(_5108__bF_buf1) );
BUFX4 BUFX4_1919 ( .gnd(gnd), .vdd(vdd), .A(_5108_), .Y(_5108__bF_buf0) );
BUFX4 BUFX4_1920 ( .gnd(gnd), .vdd(vdd), .A(_8632_), .Y(_8632__bF_buf3) );
BUFX4 BUFX4_1921 ( .gnd(gnd), .vdd(vdd), .A(_8632_), .Y(_8632__bF_buf2) );
BUFX4 BUFX4_1922 ( .gnd(gnd), .vdd(vdd), .A(_8632_), .Y(_8632__bF_buf1) );
BUFX4 BUFX4_1923 ( .gnd(gnd), .vdd(vdd), .A(_8632_), .Y(_8632__bF_buf0) );
BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(_0__bF_buf9), .Y(finished) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(_1__0_), .Y(nonce_out[0]) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(_1__1_), .Y(nonce_out[1]) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(_1__2_), .Y(nonce_out[2]) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(_1__3_), .Y(nonce_out[3]) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(_1__4_), .Y(nonce_out[4]) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_1__5_), .Y(nonce_out[5]) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_1__6_), .Y(nonce_out[6]) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(_1__7_), .Y(nonce_out[7]) );
BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(_1__8_), .Y(nonce_out[8]) );
BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(_1__9_), .Y(nonce_out[9]) );
BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(_1__10_), .Y(nonce_out[10]) );
BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(_1__11_), .Y(nonce_out[11]) );
BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(_1__12_), .Y(nonce_out[12]) );
BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(_1__13_), .Y(nonce_out[13]) );
BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(_1__14_), .Y(nonce_out[14]) );
BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(_1__15_), .Y(nonce_out[15]) );
BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(_1__16_), .Y(nonce_out[16]) );
BUFX2 BUFX2_19 ( .gnd(gnd), .vdd(vdd), .A(_1__17_), .Y(nonce_out[17]) );
BUFX2 BUFX2_20 ( .gnd(gnd), .vdd(vdd), .A(_1__18_), .Y(nonce_out[18]) );
BUFX2 BUFX2_21 ( .gnd(gnd), .vdd(vdd), .A(_1__19_), .Y(nonce_out[19]) );
BUFX2 BUFX2_22 ( .gnd(gnd), .vdd(vdd), .A(_1__20_), .Y(nonce_out[20]) );
BUFX2 BUFX2_23 ( .gnd(gnd), .vdd(vdd), .A(_1__21_), .Y(nonce_out[21]) );
BUFX2 BUFX2_24 ( .gnd(gnd), .vdd(vdd), .A(_1__22_), .Y(nonce_out[22]) );
BUFX2 BUFX2_25 ( .gnd(gnd), .vdd(vdd), .A(_1__23_), .Y(nonce_out[23]) );
BUFX2 BUFX2_26 ( .gnd(gnd), .vdd(vdd), .A(_1__24_), .Y(nonce_out[24]) );
BUFX2 BUFX2_27 ( .gnd(gnd), .vdd(vdd), .A(_1__25_), .Y(nonce_out[25]) );
BUFX2 BUFX2_28 ( .gnd(gnd), .vdd(vdd), .A(_1__26_), .Y(nonce_out[26]) );
BUFX2 BUFX2_29 ( .gnd(gnd), .vdd(vdd), .A(_1__27_), .Y(nonce_out[27]) );
BUFX2 BUFX2_30 ( .gnd(gnd), .vdd(vdd), .A(_1__28_), .Y(nonce_out[28]) );
BUFX2 BUFX2_31 ( .gnd(gnd), .vdd(vdd), .A(_1__29_), .Y(nonce_out[29]) );
BUFX2 BUFX2_32 ( .gnd(gnd), .vdd(vdd), .A(_1__30_), .Y(nonce_out[30]) );
BUFX2 BUFX2_33 ( .gnd(gnd), .vdd(vdd), .A(_1__31_), .Y(nonce_out[31]) );
INVX2 INVX2_1 ( .gnd(gnd), .vdd(vdd), .A(target[1]), .Y(_30_) );
NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(H_9_), .B(_30_), .Y(_31_) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(target[0]), .Y(_32_) );
OAI22X1 OAI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_30_), .B(H_9_), .C(_32_), .D(H_8_), .Y(_33_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_31_), .B(_33_), .Y(_34_) );
XOR2X1 XOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(target[3]), .B(H_11_), .Y(_35_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(target[2]), .B(H_10_), .Y(_36_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(target[2]), .B(H_10_), .Y(_37_) );
AOI21X1 AOI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_36_), .B(_37_), .C(_35_), .Y(_38_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(target[3]), .Y(_39_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(H_11_), .B(_39_), .Y(_40_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(target[2]), .Y(_41_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(H_10_), .B(_41_), .Y(_42_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_35_), .B(_42_), .C(_40_), .Y(_43_) );
AOI21X1 AOI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_34_), .B(_38_), .C(_43_), .Y(_44_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(H_15_), .Y(_45_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(H_14_), .Y(_46_) );
OAI22X1 OAI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_45_), .B(target_7_bF_buf3_), .C(target[6]), .D(_46_), .Y(_47_) );
INVX2 INVX2_2 ( .gnd(gnd), .vdd(vdd), .A(target_7_bF_buf2_), .Y(_48_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(target[6]), .Y(_49_) );
OAI22X1 OAI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(_48_), .B(H_15_), .C(_49_), .D(H_14_), .Y(_50_) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_47_), .B(_50_), .Y(_51_) );
INVX2 INVX2_3 ( .gnd(gnd), .vdd(vdd), .A(target[5]), .Y(_52_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(target[4]), .Y(_53_) );
AOI22X1 AOI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_52_), .B(H_13_), .C(_53_), .D(H_12_), .Y(_54_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(H_13_), .Y(_55_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(H_12_), .Y(_56_) );
AOI22X1 AOI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_55_), .B(target[5]), .C(target[4]), .D(_56_), .Y(_57_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_54_), .B(_57_), .C(_51_), .Y(_58_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(target_7_bF_buf1_), .B(_45_), .Y(_59_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(H_13_), .B(_52_), .Y(_60_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_60_), .B(_54_), .Y(_61_) );
AOI22X1 AOI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(_47_), .B(_59_), .C(_51_), .D(_61_), .Y(_62_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_44_), .B(_58_), .C(_62_), .Y(_63_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(H_17_), .B(_30_), .Y(_64_) );
OAI22X1 OAI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(_30_), .B(H_17_), .C(_32_), .D(H_16_), .Y(_65_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_64_), .B(_65_), .Y(_66_) );
XOR2X1 XOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(target[3]), .B(H_19_), .Y(_67_) );
OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(target[2]), .B(H_18_), .Y(_68_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(target[2]), .B(H_18_), .Y(_69_) );
AOI21X1 AOI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_68_), .B(_69_), .C(_67_), .Y(_70_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(H_19_), .B(_39_), .Y(_71_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(H_18_), .B(_41_), .Y(_72_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_67_), .B(_72_), .C(_71_), .Y(_73_) );
AOI21X1 AOI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_66_), .B(_70_), .C(_73_), .Y(_74_) );
INVX2 INVX2_4 ( .gnd(gnd), .vdd(vdd), .A(H_23_), .Y(_75_) );
OAI22X1 OAI22X1_5 ( .gnd(gnd), .vdd(vdd), .A(_75_), .B(target_7_bF_buf0_), .C(_49_), .D(H_22_), .Y(_76_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(H_22_), .Y(_77_) );
OAI22X1 OAI22X1_6 ( .gnd(gnd), .vdd(vdd), .A(_48_), .B(H_23_), .C(target[6]), .D(_77_), .Y(_78_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_76_), .B(_78_), .Y(_79_) );
AOI22X1 AOI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(_52_), .B(H_21_), .C(_53_), .D(H_20_), .Y(_80_) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(H_20_), .Y(_81_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(H_21_), .B(_52_), .Y(_82_) );
AOI21X1 AOI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(target[4]), .B(_81_), .C(_82_), .Y(_83_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_80_), .B(_83_), .C(_79_), .Y(_84_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_82_), .B(_80_), .Y(_85_) );
NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(target[6]), .B(_77_), .Y(_86_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_48_), .B(H_23_), .C(_86_), .Y(_87_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(target_7_bF_buf3_), .B(_75_), .C(_87_), .Y(_88_) );
AOI21X1 AOI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_85_), .B(_79_), .C(_88_), .Y(_89_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_74_), .B(_84_), .C(_89_), .Y(_90_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(comparador_valid_hash), .B(reset_bF_buf10), .Y(_91_) );
NOR3X1 NOR3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_63_), .B(_91_), .C(_90_), .Y(_3_) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_33_), .B(_31_), .Y(_92_) );
XNOR2X1 XNOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(target[3]), .B(H_11_), .Y(_93_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_37_), .B(_36_), .Y(_94_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_93_), .B(_94_), .Y(_95_) );
INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(_40_), .Y(_96_) );
INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(_42_), .Y(_97_) );
AOI21X1 AOI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_93_), .B(_97_), .C(_96_), .Y(_98_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_95_), .B(_92_), .C(_98_), .Y(_99_) );
OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(_47_), .B(_50_), .Y(_4_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_54_), .B(_57_), .Y(_5_) );
NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_5_), .B(_4_), .Y(_6_) );
OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(_54_), .B(_60_), .Y(_7_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_48_), .B(H_15_), .C(_47_), .Y(_8_) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_4_), .B(_7_), .C(_8_), .Y(_9_) );
AOI21X1 AOI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_6_), .B(_99_), .C(_9_), .Y(_10_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(_65_), .B(_64_), .Y(_11_) );
XNOR2X1 XNOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(target[3]), .B(H_19_), .Y(_12_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_69_), .B(_68_), .Y(_13_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_12_), .B(_13_), .Y(_14_) );
INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(_71_), .Y(_15_) );
INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(_72_), .Y(_16_) );
AOI21X1 AOI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_12_), .B(_16_), .C(_15_), .Y(_17_) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_14_), .B(_11_), .C(_17_), .Y(_18_) );
OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(_76_), .B(_78_), .Y(_19_) );
OR2X2 OR2X2_6 ( .gnd(gnd), .vdd(vdd), .A(_52_), .B(H_21_), .Y(_20_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(target[4]), .B(_81_), .Y(_21_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_21_), .B(_80_), .C(_20_), .Y(_22_) );
NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_22_), .B(_19_), .Y(_23_) );
OR2X2 OR2X2_7 ( .gnd(gnd), .vdd(vdd), .A(_80_), .B(_82_), .Y(_24_) );
NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(target_7_bF_buf2_), .B(_75_), .Y(_25_) );
NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(target_7_bF_buf1_), .B(_75_), .Y(_26_) );
AOI21X1 AOI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_26_), .B(_86_), .C(_25_), .Y(_27_) );
OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_19_), .B(_24_), .C(_27_), .Y(_28_) );
AOI21X1 AOI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_23_), .B(_18_), .C(_28_), .Y(_29_) );
AOI21X1 AOI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_10_), .B(_29_), .C(_91_), .Y(_2_) );
DFFPOSX1 DFFPOSX1_1 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf157), .D(_2_), .Q(comparador_next) );
DFFPOSX1 DFFPOSX1_2 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf156), .D(_3_), .Q(comparador_valid) );
INVX2 INVX2_5 ( .gnd(gnd), .vdd(vdd), .A(target[1]), .Y(_128_) );
NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(H_2_9_), .B(_128_), .Y(_129_) );
INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(target[0]), .Y(_130_) );
OAI22X1 OAI22X1_7 ( .gnd(gnd), .vdd(vdd), .A(_128_), .B(H_2_9_), .C(_130_), .D(H_2_8_), .Y(_131_) );
NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_129_), .B(_131_), .Y(_132_) );
XOR2X1 XOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(target[3]), .B(H_2_11_), .Y(_133_) );
OR2X2 OR2X2_8 ( .gnd(gnd), .vdd(vdd), .A(target[2]), .B(H_2_10_), .Y(_134_) );
NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(target[2]), .B(H_2_10_), .Y(_135_) );
AOI21X1 AOI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_134_), .B(_135_), .C(_133_), .Y(_136_) );
INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(target[3]), .Y(_137_) );
NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(H_2_11_), .B(_137_), .Y(_138_) );
INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(target[2]), .Y(_139_) );
NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(H_2_10_), .B(_139_), .Y(_140_) );
OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_133_), .B(_140_), .C(_138_), .Y(_141_) );
AOI21X1 AOI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_132_), .B(_136_), .C(_141_), .Y(_142_) );
INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(H_2_15_), .Y(_143_) );
INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(H_2_14_), .Y(_144_) );
OAI22X1 OAI22X1_8 ( .gnd(gnd), .vdd(vdd), .A(_143_), .B(target_7_bF_buf0_), .C(target[6]), .D(_144_), .Y(_145_) );
INVX2 INVX2_6 ( .gnd(gnd), .vdd(vdd), .A(target_7_bF_buf3_), .Y(_146_) );
INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(target[6]), .Y(_147_) );
OAI22X1 OAI22X1_9 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(H_2_15_), .C(_147_), .D(H_2_14_), .Y(_148_) );
NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_145_), .B(_148_), .Y(_149_) );
INVX2 INVX2_7 ( .gnd(gnd), .vdd(vdd), .A(target[5]), .Y(_150_) );
INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(target[4]), .Y(_151_) );
AOI22X1 AOI22X1_5 ( .gnd(gnd), .vdd(vdd), .A(_150_), .B(H_2_13_), .C(_151_), .D(H_2_12_), .Y(_152_) );
INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(H_2_13_), .Y(_153_) );
INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(H_2_12_), .Y(_154_) );
AOI22X1 AOI22X1_6 ( .gnd(gnd), .vdd(vdd), .A(_153_), .B(target[5]), .C(target[4]), .D(_154_), .Y(_155_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_152_), .B(_155_), .C(_149_), .Y(_156_) );
NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(target_7_bF_buf2_), .B(_143_), .Y(_157_) );
NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(H_2_13_), .B(_150_), .Y(_158_) );
NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_158_), .B(_152_), .Y(_159_) );
AOI22X1 AOI22X1_7 ( .gnd(gnd), .vdd(vdd), .A(_145_), .B(_157_), .C(_149_), .D(_159_), .Y(_160_) );
OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_142_), .B(_156_), .C(_160_), .Y(_161_) );
NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(H_2_17_), .B(_128_), .Y(_162_) );
OAI22X1 OAI22X1_10 ( .gnd(gnd), .vdd(vdd), .A(_128_), .B(H_2_17_), .C(_130_), .D(H_2_16_), .Y(_163_) );
NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_162_), .B(_163_), .Y(_164_) );
XOR2X1 XOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(target[3]), .B(H_2_19_), .Y(_165_) );
OR2X2 OR2X2_9 ( .gnd(gnd), .vdd(vdd), .A(target[2]), .B(H_2_18_), .Y(_166_) );
NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(target[2]), .B(H_2_18_), .Y(_167_) );
AOI21X1 AOI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_166_), .B(_167_), .C(_165_), .Y(_168_) );
NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(H_2_19_), .B(_137_), .Y(_169_) );
NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(H_2_18_), .B(_139_), .Y(_170_) );
OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_165_), .B(_170_), .C(_169_), .Y(_171_) );
AOI21X1 AOI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_164_), .B(_168_), .C(_171_), .Y(_172_) );
INVX2 INVX2_8 ( .gnd(gnd), .vdd(vdd), .A(H_2_23_), .Y(_173_) );
OAI22X1 OAI22X1_11 ( .gnd(gnd), .vdd(vdd), .A(_173_), .B(target_7_bF_buf1_), .C(_147_), .D(H_2_22_), .Y(_174_) );
INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(H_2_22_), .Y(_175_) );
OAI22X1 OAI22X1_12 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(H_2_23_), .C(target[6]), .D(_175_), .Y(_176_) );
NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_174_), .B(_176_), .Y(_177_) );
AOI22X1 AOI22X1_8 ( .gnd(gnd), .vdd(vdd), .A(_150_), .B(H_2_21_), .C(_151_), .D(H_2_20_), .Y(_178_) );
INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(H_2_20_), .Y(_179_) );
NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(H_2_21_), .B(_150_), .Y(_180_) );
AOI21X1 AOI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(target[4]), .B(_179_), .C(_180_), .Y(_181_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_178_), .B(_181_), .C(_177_), .Y(_182_) );
NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_180_), .B(_178_), .Y(_183_) );
NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(target[6]), .B(_175_), .Y(_184_) );
OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(H_2_23_), .C(_184_), .Y(_185_) );
OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(target_7_bF_buf0_), .B(_173_), .C(_185_), .Y(_186_) );
AOI21X1 AOI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_183_), .B(_177_), .C(_186_), .Y(_187_) );
OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_172_), .B(_182_), .C(_187_), .Y(_188_) );
NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(comparador_2_valid_hash), .B(reset_bF_buf9), .Y(_189_) );
NOR3X1 NOR3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_161_), .B(_189_), .C(_188_), .Y(_101_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(_131_), .B(_129_), .Y(_190_) );
XNOR2X1 XNOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(target[3]), .B(H_2_11_), .Y(_191_) );
NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_135_), .B(_134_), .Y(_192_) );
NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(_191_), .B(_192_), .Y(_193_) );
INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(_138_), .Y(_194_) );
INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(_140_), .Y(_195_) );
AOI21X1 AOI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_191_), .B(_195_), .C(_194_), .Y(_196_) );
OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_193_), .B(_190_), .C(_196_), .Y(_197_) );
OR2X2 OR2X2_10 ( .gnd(gnd), .vdd(vdd), .A(_145_), .B(_148_), .Y(_102_) );
NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_152_), .B(_155_), .Y(_103_) );
NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_103_), .B(_102_), .Y(_104_) );
OR2X2 OR2X2_11 ( .gnd(gnd), .vdd(vdd), .A(_152_), .B(_158_), .Y(_105_) );
OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(H_2_15_), .C(_145_), .Y(_106_) );
OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_102_), .B(_105_), .C(_106_), .Y(_107_) );
AOI21X1 AOI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_104_), .B(_197_), .C(_107_), .Y(_108_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(_163_), .B(_162_), .Y(_109_) );
XNOR2X1 XNOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(target[3]), .B(H_2_19_), .Y(_110_) );
NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_167_), .B(_166_), .Y(_111_) );
NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_110_), .B(_111_), .Y(_112_) );
INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(_169_), .Y(_113_) );
INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(_170_), .Y(_114_) );
AOI21X1 AOI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_110_), .B(_114_), .C(_113_), .Y(_115_) );
OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_112_), .B(_109_), .C(_115_), .Y(_116_) );
OR2X2 OR2X2_12 ( .gnd(gnd), .vdd(vdd), .A(_174_), .B(_176_), .Y(_117_) );
OR2X2 OR2X2_13 ( .gnd(gnd), .vdd(vdd), .A(_150_), .B(H_2_21_), .Y(_118_) );
NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(target[4]), .B(_179_), .Y(_119_) );
NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_119_), .B(_178_), .C(_118_), .Y(_120_) );
NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_120_), .B(_117_), .Y(_121_) );
OR2X2 OR2X2_14 ( .gnd(gnd), .vdd(vdd), .A(_178_), .B(_180_), .Y(_122_) );
NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(target_7_bF_buf3_), .B(_173_), .Y(_123_) );
NAND2X1 NAND2X1_38 ( .gnd(gnd), .vdd(vdd), .A(target_7_bF_buf2_), .B(_173_), .Y(_124_) );
AOI21X1 AOI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_124_), .B(_184_), .C(_123_), .Y(_125_) );
OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_117_), .B(_122_), .C(_125_), .Y(_126_) );
AOI21X1 AOI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_121_), .B(_116_), .C(_126_), .Y(_127_) );
AOI21X1 AOI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_108_), .B(_127_), .C(_189_), .Y(_100_) );
DFFPOSX1 DFFPOSX1_3 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf155), .D(_100_), .Q(comparador_next) );
DFFPOSX1 DFFPOSX1_4 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf154), .D(_101_), .Q(comparador_2_valid) );
INVX2 INVX2_9 ( .gnd(gnd), .vdd(vdd), .A(target[1]), .Y(_226_) );
NAND2X1 NAND2X1_39 ( .gnd(gnd), .vdd(vdd), .A(H_3_9_), .B(_226_), .Y(_227_) );
INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(target[0]), .Y(_228_) );
OAI22X1 OAI22X1_13 ( .gnd(gnd), .vdd(vdd), .A(_226_), .B(H_3_9_), .C(_228_), .D(H_3_8_), .Y(_229_) );
NAND2X1 NAND2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_227_), .B(_229_), .Y(_230_) );
XOR2X1 XOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(target[3]), .B(H_3_11_), .Y(_231_) );
OR2X2 OR2X2_15 ( .gnd(gnd), .vdd(vdd), .A(target[2]), .B(H_3_10_), .Y(_232_) );
NAND2X1 NAND2X1_41 ( .gnd(gnd), .vdd(vdd), .A(target[2]), .B(H_3_10_), .Y(_233_) );
AOI21X1 AOI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_232_), .B(_233_), .C(_231_), .Y(_234_) );
INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(target[3]), .Y(_235_) );
NAND2X1 NAND2X1_42 ( .gnd(gnd), .vdd(vdd), .A(H_3_11_), .B(_235_), .Y(_236_) );
INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(target[2]), .Y(_237_) );
NAND2X1 NAND2X1_43 ( .gnd(gnd), .vdd(vdd), .A(H_3_10_), .B(_237_), .Y(_238_) );
OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_231_), .B(_238_), .C(_236_), .Y(_239_) );
AOI21X1 AOI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_230_), .B(_234_), .C(_239_), .Y(_240_) );
INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(H_3_15_), .Y(_241_) );
INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(H_3_14_), .Y(_242_) );
OAI22X1 OAI22X1_14 ( .gnd(gnd), .vdd(vdd), .A(_241_), .B(target_7_bF_buf1_), .C(target[6]), .D(_242_), .Y(_243_) );
INVX2 INVX2_10 ( .gnd(gnd), .vdd(vdd), .A(target_7_bF_buf0_), .Y(_244_) );
INVX1 INVX1_36 ( .gnd(gnd), .vdd(vdd), .A(target[6]), .Y(_245_) );
OAI22X1 OAI22X1_15 ( .gnd(gnd), .vdd(vdd), .A(_244_), .B(H_3_15_), .C(_245_), .D(H_3_14_), .Y(_246_) );
NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_243_), .B(_246_), .Y(_247_) );
INVX2 INVX2_11 ( .gnd(gnd), .vdd(vdd), .A(target[5]), .Y(_248_) );
INVX1 INVX1_37 ( .gnd(gnd), .vdd(vdd), .A(target[4]), .Y(_249_) );
AOI22X1 AOI22X1_9 ( .gnd(gnd), .vdd(vdd), .A(_248_), .B(H_3_13_), .C(_249_), .D(H_3_12_), .Y(_250_) );
INVX1 INVX1_38 ( .gnd(gnd), .vdd(vdd), .A(H_3_13_), .Y(_251_) );
INVX1 INVX1_39 ( .gnd(gnd), .vdd(vdd), .A(H_3_12_), .Y(_252_) );
AOI22X1 AOI22X1_10 ( .gnd(gnd), .vdd(vdd), .A(_251_), .B(target[5]), .C(target[4]), .D(_252_), .Y(_253_) );
NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_250_), .B(_253_), .C(_247_), .Y(_254_) );
NAND2X1 NAND2X1_44 ( .gnd(gnd), .vdd(vdd), .A(target_7_bF_buf3_), .B(_241_), .Y(_255_) );
NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(H_3_13_), .B(_248_), .Y(_256_) );
NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_256_), .B(_250_), .Y(_257_) );
AOI22X1 AOI22X1_11 ( .gnd(gnd), .vdd(vdd), .A(_243_), .B(_255_), .C(_247_), .D(_257_), .Y(_258_) );
OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_240_), .B(_254_), .C(_258_), .Y(_259_) );
NAND2X1 NAND2X1_45 ( .gnd(gnd), .vdd(vdd), .A(H_3_17_), .B(_226_), .Y(_260_) );
OAI22X1 OAI22X1_16 ( .gnd(gnd), .vdd(vdd), .A(_226_), .B(H_3_17_), .C(_228_), .D(H_3_16_), .Y(_261_) );
NAND2X1 NAND2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_260_), .B(_261_), .Y(_262_) );
XOR2X1 XOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(target[3]), .B(H_3_19_), .Y(_263_) );
OR2X2 OR2X2_16 ( .gnd(gnd), .vdd(vdd), .A(target[2]), .B(H_3_18_), .Y(_264_) );
NAND2X1 NAND2X1_47 ( .gnd(gnd), .vdd(vdd), .A(target[2]), .B(H_3_18_), .Y(_265_) );
AOI21X1 AOI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_264_), .B(_265_), .C(_263_), .Y(_266_) );
NAND2X1 NAND2X1_48 ( .gnd(gnd), .vdd(vdd), .A(H_3_19_), .B(_235_), .Y(_267_) );
NAND2X1 NAND2X1_49 ( .gnd(gnd), .vdd(vdd), .A(H_3_18_), .B(_237_), .Y(_268_) );
OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_263_), .B(_268_), .C(_267_), .Y(_269_) );
AOI21X1 AOI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_262_), .B(_266_), .C(_269_), .Y(_270_) );
INVX2 INVX2_12 ( .gnd(gnd), .vdd(vdd), .A(H_3_23_), .Y(_271_) );
OAI22X1 OAI22X1_17 ( .gnd(gnd), .vdd(vdd), .A(_271_), .B(target_7_bF_buf2_), .C(_245_), .D(H_3_22_), .Y(_272_) );
INVX1 INVX1_40 ( .gnd(gnd), .vdd(vdd), .A(H_3_22_), .Y(_273_) );
OAI22X1 OAI22X1_18 ( .gnd(gnd), .vdd(vdd), .A(_244_), .B(H_3_23_), .C(target[6]), .D(_273_), .Y(_274_) );
NOR2X1 NOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_272_), .B(_274_), .Y(_275_) );
AOI22X1 AOI22X1_12 ( .gnd(gnd), .vdd(vdd), .A(_248_), .B(H_3_21_), .C(_249_), .D(H_3_20_), .Y(_276_) );
INVX1 INVX1_41 ( .gnd(gnd), .vdd(vdd), .A(H_3_20_), .Y(_277_) );
NOR2X1 NOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(H_3_21_), .B(_248_), .Y(_278_) );
AOI21X1 AOI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(target[4]), .B(_277_), .C(_278_), .Y(_279_) );
NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_276_), .B(_279_), .C(_275_), .Y(_280_) );
NOR2X1 NOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_278_), .B(_276_), .Y(_281_) );
NOR2X1 NOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(target[6]), .B(_273_), .Y(_282_) );
OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_244_), .B(H_3_23_), .C(_282_), .Y(_283_) );
OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(target_7_bF_buf1_), .B(_271_), .C(_283_), .Y(_284_) );
AOI21X1 AOI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_281_), .B(_275_), .C(_284_), .Y(_285_) );
OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_270_), .B(_280_), .C(_285_), .Y(_286_) );
NAND2X1 NAND2X1_50 ( .gnd(gnd), .vdd(vdd), .A(comparador_3_valid_hash), .B(reset_bF_buf8), .Y(_287_) );
NOR3X1 NOR3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_259_), .B(_287_), .C(_286_), .Y(_199_) );
AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(_229_), .B(_227_), .Y(_288_) );
XNOR2X1 XNOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(target[3]), .B(H_3_11_), .Y(_289_) );
NAND2X1 NAND2X1_51 ( .gnd(gnd), .vdd(vdd), .A(_233_), .B(_232_), .Y(_290_) );
NAND2X1 NAND2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_289_), .B(_290_), .Y(_291_) );
INVX1 INVX1_42 ( .gnd(gnd), .vdd(vdd), .A(_236_), .Y(_292_) );
INVX1 INVX1_43 ( .gnd(gnd), .vdd(vdd), .A(_238_), .Y(_293_) );
AOI21X1 AOI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_289_), .B(_293_), .C(_292_), .Y(_294_) );
OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_291_), .B(_288_), .C(_294_), .Y(_295_) );
OR2X2 OR2X2_17 ( .gnd(gnd), .vdd(vdd), .A(_243_), .B(_246_), .Y(_200_) );
NAND2X1 NAND2X1_53 ( .gnd(gnd), .vdd(vdd), .A(_250_), .B(_253_), .Y(_201_) );
NOR2X1 NOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_201_), .B(_200_), .Y(_202_) );
OR2X2 OR2X2_18 ( .gnd(gnd), .vdd(vdd), .A(_250_), .B(_256_), .Y(_203_) );
OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_244_), .B(H_3_15_), .C(_243_), .Y(_204_) );
OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_200_), .B(_203_), .C(_204_), .Y(_205_) );
AOI21X1 AOI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_202_), .B(_295_), .C(_205_), .Y(_206_) );
AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(_261_), .B(_260_), .Y(_207_) );
XNOR2X1 XNOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(target[3]), .B(H_3_19_), .Y(_208_) );
NAND2X1 NAND2X1_54 ( .gnd(gnd), .vdd(vdd), .A(_265_), .B(_264_), .Y(_209_) );
NAND2X1 NAND2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_208_), .B(_209_), .Y(_210_) );
INVX1 INVX1_44 ( .gnd(gnd), .vdd(vdd), .A(_267_), .Y(_211_) );
INVX1 INVX1_45 ( .gnd(gnd), .vdd(vdd), .A(_268_), .Y(_212_) );
AOI21X1 AOI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_208_), .B(_212_), .C(_211_), .Y(_213_) );
OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_210_), .B(_207_), .C(_213_), .Y(_214_) );
OR2X2 OR2X2_19 ( .gnd(gnd), .vdd(vdd), .A(_272_), .B(_274_), .Y(_215_) );
OR2X2 OR2X2_20 ( .gnd(gnd), .vdd(vdd), .A(_248_), .B(H_3_21_), .Y(_216_) );
NAND2X1 NAND2X1_56 ( .gnd(gnd), .vdd(vdd), .A(target[4]), .B(_277_), .Y(_217_) );
NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_217_), .B(_276_), .C(_216_), .Y(_218_) );
NOR2X1 NOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_218_), .B(_215_), .Y(_219_) );
OR2X2 OR2X2_21 ( .gnd(gnd), .vdd(vdd), .A(_276_), .B(_278_), .Y(_220_) );
NOR2X1 NOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(target_7_bF_buf0_), .B(_271_), .Y(_221_) );
NAND2X1 NAND2X1_57 ( .gnd(gnd), .vdd(vdd), .A(target_7_bF_buf3_), .B(_271_), .Y(_222_) );
AOI21X1 AOI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_222_), .B(_282_), .C(_221_), .Y(_223_) );
OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_215_), .B(_220_), .C(_223_), .Y(_224_) );
AOI21X1 AOI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_219_), .B(_214_), .C(_224_), .Y(_225_) );
AOI21X1 AOI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_206_), .B(_225_), .C(_287_), .Y(_198_) );
DFFPOSX1 DFFPOSX1_5 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf153), .D(_198_), .Q(comparador_next) );
DFFPOSX1 DFFPOSX1_6 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf152), .D(_199_), .Q(comparador_3_valid) );
DFFPOSX1 DFFPOSX1_7 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf151), .D(concatenador_nonce_0_), .Q(concatenador_data_out_0_) );
DFFPOSX1 DFFPOSX1_8 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf150), .D(concatenador_nonce_1_), .Q(concatenador_data_out_1_) );
DFFPOSX1 DFFPOSX1_9 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf149), .D(concatenador_nonce_2_), .Q(concatenador_data_out_2_) );
DFFPOSX1 DFFPOSX1_10 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf148), .D(concatenador_nonce_3_), .Q(concatenador_data_out_3_) );
DFFPOSX1 DFFPOSX1_11 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf147), .D(concatenador_nonce_4_), .Q(concatenador_data_out_4_) );
DFFPOSX1 DFFPOSX1_12 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf146), .D(concatenador_nonce_5_), .Q(concatenador_data_out_5_) );
DFFPOSX1 DFFPOSX1_13 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf145), .D(concatenador_nonce_6_), .Q(concatenador_data_out_6_) );
DFFPOSX1 DFFPOSX1_14 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf144), .D(concatenador_nonce_7_), .Q(concatenador_data_out_7_) );
DFFPOSX1 DFFPOSX1_15 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf143), .D(concatenador_nonce_8_), .Q(concatenador_data_out_8_) );
DFFPOSX1 DFFPOSX1_16 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf142), .D(concatenador_nonce_9_), .Q(concatenador_data_out_9_) );
DFFPOSX1 DFFPOSX1_17 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf141), .D(concatenador_nonce_10_), .Q(concatenador_data_out_10_) );
DFFPOSX1 DFFPOSX1_18 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf140), .D(concatenador_nonce_11_), .Q(concatenador_data_out_11_) );
DFFPOSX1 DFFPOSX1_19 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf139), .D(concatenador_nonce_12_), .Q(concatenador_data_out_12_) );
DFFPOSX1 DFFPOSX1_20 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf138), .D(concatenador_nonce_13_), .Q(concatenador_data_out_13_) );
DFFPOSX1 DFFPOSX1_21 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf137), .D(concatenador_nonce_14_), .Q(concatenador_data_out_14_) );
DFFPOSX1 DFFPOSX1_22 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf136), .D(concatenador_nonce_15_), .Q(concatenador_data_out_15_) );
DFFPOSX1 DFFPOSX1_23 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf135), .D(concatenador_nonce_16_), .Q(concatenador_data_out_16_) );
DFFPOSX1 DFFPOSX1_24 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf134), .D(concatenador_nonce_17_), .Q(concatenador_data_out_17_) );
DFFPOSX1 DFFPOSX1_25 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf133), .D(concatenador_nonce_18_), .Q(concatenador_data_out_18_) );
DFFPOSX1 DFFPOSX1_26 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf132), .D(concatenador_nonce_19_), .Q(concatenador_data_out_19_) );
DFFPOSX1 DFFPOSX1_27 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf131), .D(concatenador_nonce_20_), .Q(concatenador_data_out_20_) );
DFFPOSX1 DFFPOSX1_28 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf130), .D(concatenador_nonce_21_), .Q(concatenador_data_out_21_) );
DFFPOSX1 DFFPOSX1_29 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf129), .D(concatenador_nonce_22_), .Q(concatenador_data_out_22_) );
DFFPOSX1 DFFPOSX1_30 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf128), .D(concatenador_nonce_23_), .Q(concatenador_data_out_23_) );
DFFPOSX1 DFFPOSX1_31 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf127), .D(concatenador_nonce_24_), .Q(concatenador_data_out_24_) );
DFFPOSX1 DFFPOSX1_32 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf126), .D(concatenador_nonce_25_), .Q(concatenador_data_out_25_) );
DFFPOSX1 DFFPOSX1_33 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf125), .D(concatenador_nonce_26_), .Q(concatenador_data_out_26_) );
DFFPOSX1 DFFPOSX1_34 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf124), .D(concatenador_nonce_27_), .Q(concatenador_data_out_27_) );
DFFPOSX1 DFFPOSX1_35 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf123), .D(concatenador_nonce_28_), .Q(concatenador_data_out_28_) );
DFFPOSX1 DFFPOSX1_36 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf122), .D(concatenador_nonce_29_), .Q(concatenador_data_out_29_) );
DFFPOSX1 DFFPOSX1_37 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf121), .D(concatenador_nonce_30_), .Q(concatenador_data_out_30_) );
DFFPOSX1 DFFPOSX1_38 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf120), .D(concatenador_nonce_31_), .Q(concatenador_data_out_31_) );
DFFPOSX1 DFFPOSX1_39 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf119), .D(concatenador_bloque_0_), .Q(concatenador_data_out_32_) );
DFFPOSX1 DFFPOSX1_40 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf118), .D(concatenador_bloque_1_), .Q(concatenador_data_out_33_) );
DFFPOSX1 DFFPOSX1_41 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf117), .D(concatenador_bloque_2_), .Q(concatenador_data_out_34_) );
DFFPOSX1 DFFPOSX1_42 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf116), .D(concatenador_bloque_3_), .Q(concatenador_data_out_35_) );
DFFPOSX1 DFFPOSX1_43 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf115), .D(concatenador_bloque_4_), .Q(concatenador_data_out_36_) );
DFFPOSX1 DFFPOSX1_44 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf114), .D(concatenador_bloque_5_), .Q(concatenador_data_out_37_) );
DFFPOSX1 DFFPOSX1_45 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf113), .D(concatenador_bloque_6_), .Q(concatenador_data_out_38_) );
DFFPOSX1 DFFPOSX1_46 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf112), .D(concatenador_bloque_7_), .Q(concatenador_data_out_39_) );
DFFPOSX1 DFFPOSX1_47 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf111), .D(concatenador_bloque_8_), .Q(concatenador_data_out_40_) );
DFFPOSX1 DFFPOSX1_48 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf110), .D(concatenador_bloque_9_), .Q(concatenador_data_out_41_) );
DFFPOSX1 DFFPOSX1_49 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf109), .D(concatenador_bloque_10_), .Q(concatenador_data_out_42_) );
DFFPOSX1 DFFPOSX1_50 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf108), .D(concatenador_bloque_11_), .Q(concatenador_data_out_43_) );
DFFPOSX1 DFFPOSX1_51 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf107), .D(concatenador_bloque_12_), .Q(concatenador_data_out_44_) );
DFFPOSX1 DFFPOSX1_52 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(concatenador_bloque_13_), .Q(concatenador_data_out_45_) );
DFFPOSX1 DFFPOSX1_53 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(concatenador_bloque_14_), .Q(concatenador_data_out_46_) );
DFFPOSX1 DFFPOSX1_54 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(concatenador_bloque_15_), .Q(concatenador_data_out_47_) );
DFFPOSX1 DFFPOSX1_55 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(concatenador_bloque_16_), .Q(concatenador_data_out_48_) );
DFFPOSX1 DFFPOSX1_56 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(concatenador_bloque_17_), .Q(concatenador_data_out_49_) );
DFFPOSX1 DFFPOSX1_57 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(concatenador_bloque_18_), .Q(concatenador_data_out_50_) );
DFFPOSX1 DFFPOSX1_58 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(concatenador_bloque_19_), .Q(concatenador_data_out_51_) );
DFFPOSX1 DFFPOSX1_59 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(concatenador_bloque_20_), .Q(concatenador_data_out_52_) );
DFFPOSX1 DFFPOSX1_60 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(concatenador_bloque_21_), .Q(concatenador_data_out_53_) );
DFFPOSX1 DFFPOSX1_61 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(concatenador_bloque_22_), .Q(concatenador_data_out_54_) );
DFFPOSX1 DFFPOSX1_62 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(concatenador_bloque_23_), .Q(concatenador_data_out_55_) );
DFFPOSX1 DFFPOSX1_63 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(concatenador_bloque_24_), .Q(concatenador_data_out_56_) );
DFFPOSX1 DFFPOSX1_64 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(concatenador_bloque_25_), .Q(concatenador_data_out_57_) );
DFFPOSX1 DFFPOSX1_65 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(concatenador_bloque_26_), .Q(concatenador_data_out_58_) );
DFFPOSX1 DFFPOSX1_66 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(concatenador_bloque_27_), .Q(concatenador_data_out_59_) );
DFFPOSX1 DFFPOSX1_67 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(concatenador_bloque_28_), .Q(concatenador_data_out_60_) );
DFFPOSX1 DFFPOSX1_68 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(concatenador_bloque_29_), .Q(concatenador_data_out_61_) );
DFFPOSX1 DFFPOSX1_69 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(concatenador_bloque_30_), .Q(concatenador_data_out_62_) );
DFFPOSX1 DFFPOSX1_70 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(concatenador_bloque_31_), .Q(concatenador_data_out_63_) );
DFFPOSX1 DFFPOSX1_71 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(concatenador_bloque_32_), .Q(concatenador_data_out_64_) );
DFFPOSX1 DFFPOSX1_72 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(concatenador_bloque_33_), .Q(concatenador_data_out_65_) );
DFFPOSX1 DFFPOSX1_73 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(concatenador_bloque_34_), .Q(concatenador_data_out_66_) );
DFFPOSX1 DFFPOSX1_74 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(concatenador_bloque_35_), .Q(concatenador_data_out_67_) );
DFFPOSX1 DFFPOSX1_75 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(concatenador_bloque_36_), .Q(concatenador_data_out_68_) );
DFFPOSX1 DFFPOSX1_76 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(concatenador_bloque_37_), .Q(concatenador_data_out_69_) );
DFFPOSX1 DFFPOSX1_77 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(concatenador_bloque_38_), .Q(concatenador_data_out_70_) );
DFFPOSX1 DFFPOSX1_78 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(concatenador_bloque_39_), .Q(concatenador_data_out_71_) );
DFFPOSX1 DFFPOSX1_79 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(concatenador_bloque_40_), .Q(concatenador_data_out_72_) );
DFFPOSX1 DFFPOSX1_80 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(concatenador_bloque_41_), .Q(concatenador_data_out_73_) );
DFFPOSX1 DFFPOSX1_81 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(concatenador_bloque_42_), .Q(concatenador_data_out_74_) );
DFFPOSX1 DFFPOSX1_82 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(concatenador_bloque_43_), .Q(concatenador_data_out_75_) );
DFFPOSX1 DFFPOSX1_83 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(concatenador_bloque_44_), .Q(concatenador_data_out_76_) );
DFFPOSX1 DFFPOSX1_84 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(concatenador_bloque_45_), .Q(concatenador_data_out_77_) );
DFFPOSX1 DFFPOSX1_85 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(concatenador_bloque_46_), .Q(concatenador_data_out_78_) );
DFFPOSX1 DFFPOSX1_86 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(concatenador_bloque_47_), .Q(concatenador_data_out_79_) );
DFFPOSX1 DFFPOSX1_87 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(concatenador_bloque_48_), .Q(concatenador_data_out_80_) );
DFFPOSX1 DFFPOSX1_88 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(concatenador_bloque_49_), .Q(concatenador_data_out_81_) );
DFFPOSX1 DFFPOSX1_89 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(concatenador_bloque_50_), .Q(concatenador_data_out_82_) );
DFFPOSX1 DFFPOSX1_90 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(concatenador_bloque_51_), .Q(concatenador_data_out_83_) );
DFFPOSX1 DFFPOSX1_91 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(concatenador_bloque_52_), .Q(concatenador_data_out_84_) );
DFFPOSX1 DFFPOSX1_92 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(concatenador_bloque_53_), .Q(concatenador_data_out_85_) );
DFFPOSX1 DFFPOSX1_93 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(concatenador_bloque_54_), .Q(concatenador_data_out_86_) );
DFFPOSX1 DFFPOSX1_94 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(concatenador_bloque_55_), .Q(concatenador_data_out_87_) );
DFFPOSX1 DFFPOSX1_95 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(concatenador_bloque_56_), .Q(concatenador_data_out_88_) );
DFFPOSX1 DFFPOSX1_96 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(concatenador_bloque_57_), .Q(concatenador_data_out_89_) );
DFFPOSX1 DFFPOSX1_97 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(concatenador_bloque_58_), .Q(concatenador_data_out_90_) );
DFFPOSX1 DFFPOSX1_98 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(concatenador_bloque_59_), .Q(concatenador_data_out_91_) );
DFFPOSX1 DFFPOSX1_99 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(concatenador_bloque_60_), .Q(concatenador_data_out_92_) );
DFFPOSX1 DFFPOSX1_100 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(concatenador_bloque_61_), .Q(concatenador_data_out_93_) );
DFFPOSX1 DFFPOSX1_101 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(concatenador_bloque_62_), .Q(concatenador_data_out_94_) );
DFFPOSX1 DFFPOSX1_102 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(concatenador_bloque_63_), .Q(concatenador_data_out_95_) );
DFFPOSX1 DFFPOSX1_103 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(concatenador_bloque_64_), .Q(concatenador_data_out_96_) );
DFFPOSX1 DFFPOSX1_104 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(concatenador_bloque_65_), .Q(concatenador_data_out_97_) );
DFFPOSX1 DFFPOSX1_105 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(concatenador_bloque_66_), .Q(concatenador_data_out_98_) );
DFFPOSX1 DFFPOSX1_106 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(concatenador_bloque_67_), .Q(concatenador_data_out_99_) );
DFFPOSX1 DFFPOSX1_107 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(concatenador_bloque_68_), .Q(concatenador_data_out_100_) );
DFFPOSX1 DFFPOSX1_108 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(concatenador_bloque_69_), .Q(concatenador_data_out_101_) );
DFFPOSX1 DFFPOSX1_109 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(concatenador_bloque_70_), .Q(concatenador_data_out_102_) );
DFFPOSX1 DFFPOSX1_110 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(concatenador_bloque_71_), .Q(concatenador_data_out_103_) );
DFFPOSX1 DFFPOSX1_111 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(concatenador_bloque_72_), .Q(concatenador_data_out_104_) );
DFFPOSX1 DFFPOSX1_112 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(concatenador_bloque_73_), .Q(concatenador_data_out_105_) );
DFFPOSX1 DFFPOSX1_113 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(concatenador_bloque_74_), .Q(concatenador_data_out_106_) );
DFFPOSX1 DFFPOSX1_114 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(concatenador_bloque_75_), .Q(concatenador_data_out_107_) );
DFFPOSX1 DFFPOSX1_115 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(concatenador_bloque_76_), .Q(concatenador_data_out_108_) );
DFFPOSX1 DFFPOSX1_116 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(concatenador_bloque_77_), .Q(concatenador_data_out_109_) );
DFFPOSX1 DFFPOSX1_117 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(concatenador_bloque_78_), .Q(concatenador_data_out_110_) );
DFFPOSX1 DFFPOSX1_118 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(concatenador_bloque_79_), .Q(concatenador_data_out_111_) );
DFFPOSX1 DFFPOSX1_119 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(concatenador_bloque_80_), .Q(concatenador_data_out_112_) );
DFFPOSX1 DFFPOSX1_120 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(concatenador_bloque_81_), .Q(concatenador_data_out_113_) );
DFFPOSX1 DFFPOSX1_121 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(concatenador_bloque_82_), .Q(concatenador_data_out_114_) );
DFFPOSX1 DFFPOSX1_122 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(concatenador_bloque_83_), .Q(concatenador_data_out_115_) );
DFFPOSX1 DFFPOSX1_123 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(concatenador_bloque_84_), .Q(concatenador_data_out_116_) );
DFFPOSX1 DFFPOSX1_124 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(concatenador_bloque_85_), .Q(concatenador_data_out_117_) );
DFFPOSX1 DFFPOSX1_125 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(concatenador_bloque_86_), .Q(concatenador_data_out_118_) );
DFFPOSX1 DFFPOSX1_126 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(concatenador_bloque_87_), .Q(concatenador_data_out_119_) );
DFFPOSX1 DFFPOSX1_127 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(concatenador_bloque_88_), .Q(concatenador_data_out_120_) );
DFFPOSX1 DFFPOSX1_128 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(concatenador_bloque_89_), .Q(concatenador_data_out_121_) );
DFFPOSX1 DFFPOSX1_129 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(concatenador_bloque_90_), .Q(concatenador_data_out_122_) );
DFFPOSX1 DFFPOSX1_130 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(concatenador_bloque_91_), .Q(concatenador_data_out_123_) );
DFFPOSX1 DFFPOSX1_131 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(concatenador_bloque_92_), .Q(concatenador_data_out_124_) );
DFFPOSX1 DFFPOSX1_132 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(concatenador_bloque_93_), .Q(concatenador_data_out_125_) );
DFFPOSX1 DFFPOSX1_133 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(concatenador_bloque_94_), .Q(concatenador_data_out_126_) );
DFFPOSX1 DFFPOSX1_134 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(concatenador_bloque_95_), .Q(concatenador_data_out_127_) );
DFFPOSX1 DFFPOSX1_135 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(concatenador_2_nonce_0_), .Q(concatenador_2_data_out_0_) );
DFFPOSX1 DFFPOSX1_136 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(concatenador_2_nonce_1_), .Q(concatenador_2_data_out_1_) );
DFFPOSX1 DFFPOSX1_137 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(concatenador_2_nonce_2_), .Q(concatenador_2_data_out_2_) );
DFFPOSX1 DFFPOSX1_138 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(concatenador_2_nonce_3_), .Q(concatenador_2_data_out_3_) );
DFFPOSX1 DFFPOSX1_139 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(concatenador_2_nonce_4_), .Q(concatenador_2_data_out_4_) );
DFFPOSX1 DFFPOSX1_140 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(concatenador_2_nonce_5_), .Q(concatenador_2_data_out_5_) );
DFFPOSX1 DFFPOSX1_141 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(concatenador_2_nonce_6_), .Q(concatenador_2_data_out_6_) );
DFFPOSX1 DFFPOSX1_142 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(concatenador_2_nonce_7_), .Q(concatenador_2_data_out_7_) );
DFFPOSX1 DFFPOSX1_143 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(concatenador_2_nonce_8_), .Q(concatenador_2_data_out_8_) );
DFFPOSX1 DFFPOSX1_144 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(concatenador_2_nonce_9_), .Q(concatenador_2_data_out_9_) );
DFFPOSX1 DFFPOSX1_145 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(concatenador_2_nonce_10_), .Q(concatenador_2_data_out_10_) );
DFFPOSX1 DFFPOSX1_146 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(concatenador_2_nonce_11_), .Q(concatenador_2_data_out_11_) );
DFFPOSX1 DFFPOSX1_147 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(concatenador_2_nonce_12_), .Q(concatenador_2_data_out_12_) );
DFFPOSX1 DFFPOSX1_148 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(concatenador_2_nonce_13_), .Q(concatenador_2_data_out_13_) );
DFFPOSX1 DFFPOSX1_149 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(concatenador_2_nonce_14_), .Q(concatenador_2_data_out_14_) );
DFFPOSX1 DFFPOSX1_150 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(concatenador_2_nonce_15_), .Q(concatenador_2_data_out_15_) );
DFFPOSX1 DFFPOSX1_151 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(concatenador_2_nonce_16_), .Q(concatenador_2_data_out_16_) );
DFFPOSX1 DFFPOSX1_152 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(concatenador_2_nonce_17_), .Q(concatenador_2_data_out_17_) );
DFFPOSX1 DFFPOSX1_153 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(concatenador_2_nonce_18_), .Q(concatenador_2_data_out_18_) );
DFFPOSX1 DFFPOSX1_154 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(concatenador_2_nonce_19_), .Q(concatenador_2_data_out_19_) );
DFFPOSX1 DFFPOSX1_155 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(concatenador_2_nonce_20_), .Q(concatenador_2_data_out_20_) );
DFFPOSX1 DFFPOSX1_156 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(concatenador_2_nonce_21_), .Q(concatenador_2_data_out_21_) );
DFFPOSX1 DFFPOSX1_157 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(concatenador_2_nonce_22_), .Q(concatenador_2_data_out_22_) );
DFFPOSX1 DFFPOSX1_158 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(concatenador_2_nonce_23_), .Q(concatenador_2_data_out_23_) );
DFFPOSX1 DFFPOSX1_159 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf157), .D(concatenador_2_nonce_24_), .Q(concatenador_2_data_out_24_) );
DFFPOSX1 DFFPOSX1_160 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf156), .D(concatenador_2_nonce_25_), .Q(concatenador_2_data_out_25_) );
DFFPOSX1 DFFPOSX1_161 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf155), .D(concatenador_2_nonce_26_), .Q(concatenador_2_data_out_26_) );
DFFPOSX1 DFFPOSX1_162 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf154), .D(concatenador_2_nonce_27_), .Q(concatenador_2_data_out_27_) );
DFFPOSX1 DFFPOSX1_163 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf153), .D(concatenador_2_nonce_28_), .Q(concatenador_2_data_out_28_) );
DFFPOSX1 DFFPOSX1_164 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf152), .D(concatenador_2_nonce_29_), .Q(concatenador_2_data_out_29_) );
DFFPOSX1 DFFPOSX1_165 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf151), .D(concatenador_2_nonce_30_), .Q(concatenador_2_data_out_30_) );
DFFPOSX1 DFFPOSX1_166 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf150), .D(concatenador_2_nonce_31_), .Q(concatenador_2_data_out_31_) );
DFFPOSX1 DFFPOSX1_167 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf149), .D(concatenador_bloque_0_), .Q(concatenador_2_data_out_32_) );
DFFPOSX1 DFFPOSX1_168 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf148), .D(concatenador_bloque_1_), .Q(concatenador_2_data_out_33_) );
DFFPOSX1 DFFPOSX1_169 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf147), .D(concatenador_bloque_2_), .Q(concatenador_2_data_out_34_) );
DFFPOSX1 DFFPOSX1_170 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf146), .D(concatenador_bloque_3_), .Q(concatenador_2_data_out_35_) );
DFFPOSX1 DFFPOSX1_171 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf145), .D(concatenador_bloque_4_), .Q(concatenador_2_data_out_36_) );
DFFPOSX1 DFFPOSX1_172 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf144), .D(concatenador_bloque_5_), .Q(concatenador_2_data_out_37_) );
DFFPOSX1 DFFPOSX1_173 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf143), .D(concatenador_bloque_6_), .Q(concatenador_2_data_out_38_) );
DFFPOSX1 DFFPOSX1_174 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf142), .D(concatenador_bloque_7_), .Q(concatenador_2_data_out_39_) );
DFFPOSX1 DFFPOSX1_175 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf141), .D(concatenador_bloque_8_), .Q(concatenador_2_data_out_40_) );
DFFPOSX1 DFFPOSX1_176 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf140), .D(concatenador_bloque_9_), .Q(concatenador_2_data_out_41_) );
DFFPOSX1 DFFPOSX1_177 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf139), .D(concatenador_bloque_10_), .Q(concatenador_2_data_out_42_) );
DFFPOSX1 DFFPOSX1_178 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf138), .D(concatenador_bloque_11_), .Q(concatenador_2_data_out_43_) );
DFFPOSX1 DFFPOSX1_179 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf137), .D(concatenador_bloque_12_), .Q(concatenador_2_data_out_44_) );
DFFPOSX1 DFFPOSX1_180 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf136), .D(concatenador_bloque_13_), .Q(concatenador_2_data_out_45_) );
DFFPOSX1 DFFPOSX1_181 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf135), .D(concatenador_bloque_14_), .Q(concatenador_2_data_out_46_) );
DFFPOSX1 DFFPOSX1_182 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf134), .D(concatenador_bloque_15_), .Q(concatenador_2_data_out_47_) );
DFFPOSX1 DFFPOSX1_183 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf133), .D(concatenador_bloque_16_), .Q(concatenador_2_data_out_48_) );
DFFPOSX1 DFFPOSX1_184 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf132), .D(concatenador_bloque_17_), .Q(concatenador_2_data_out_49_) );
DFFPOSX1 DFFPOSX1_185 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf131), .D(concatenador_bloque_18_), .Q(concatenador_2_data_out_50_) );
DFFPOSX1 DFFPOSX1_186 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf130), .D(concatenador_bloque_19_), .Q(concatenador_2_data_out_51_) );
DFFPOSX1 DFFPOSX1_187 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf129), .D(concatenador_bloque_20_), .Q(concatenador_2_data_out_52_) );
DFFPOSX1 DFFPOSX1_188 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf128), .D(concatenador_bloque_21_), .Q(concatenador_2_data_out_53_) );
DFFPOSX1 DFFPOSX1_189 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf127), .D(concatenador_bloque_22_), .Q(concatenador_2_data_out_54_) );
DFFPOSX1 DFFPOSX1_190 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf126), .D(concatenador_bloque_23_), .Q(concatenador_2_data_out_55_) );
DFFPOSX1 DFFPOSX1_191 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf125), .D(concatenador_bloque_24_), .Q(concatenador_2_data_out_56_) );
DFFPOSX1 DFFPOSX1_192 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf124), .D(concatenador_bloque_25_), .Q(concatenador_2_data_out_57_) );
DFFPOSX1 DFFPOSX1_193 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf123), .D(concatenador_bloque_26_), .Q(concatenador_2_data_out_58_) );
DFFPOSX1 DFFPOSX1_194 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf122), .D(concatenador_bloque_27_), .Q(concatenador_2_data_out_59_) );
DFFPOSX1 DFFPOSX1_195 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf121), .D(concatenador_bloque_28_), .Q(concatenador_2_data_out_60_) );
DFFPOSX1 DFFPOSX1_196 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf120), .D(concatenador_bloque_29_), .Q(concatenador_2_data_out_61_) );
DFFPOSX1 DFFPOSX1_197 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf119), .D(concatenador_bloque_30_), .Q(concatenador_2_data_out_62_) );
DFFPOSX1 DFFPOSX1_198 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf118), .D(concatenador_bloque_31_), .Q(concatenador_2_data_out_63_) );
DFFPOSX1 DFFPOSX1_199 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf117), .D(concatenador_bloque_32_), .Q(concatenador_2_data_out_64_) );
DFFPOSX1 DFFPOSX1_200 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf116), .D(concatenador_bloque_33_), .Q(concatenador_2_data_out_65_) );
DFFPOSX1 DFFPOSX1_201 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf115), .D(concatenador_bloque_34_), .Q(concatenador_2_data_out_66_) );
DFFPOSX1 DFFPOSX1_202 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf114), .D(concatenador_bloque_35_), .Q(concatenador_2_data_out_67_) );
DFFPOSX1 DFFPOSX1_203 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf113), .D(concatenador_bloque_36_), .Q(concatenador_2_data_out_68_) );
DFFPOSX1 DFFPOSX1_204 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf112), .D(concatenador_bloque_37_), .Q(concatenador_2_data_out_69_) );
DFFPOSX1 DFFPOSX1_205 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf111), .D(concatenador_bloque_38_), .Q(concatenador_2_data_out_70_) );
DFFPOSX1 DFFPOSX1_206 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf110), .D(concatenador_bloque_39_), .Q(concatenador_2_data_out_71_) );
DFFPOSX1 DFFPOSX1_207 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf109), .D(concatenador_bloque_40_), .Q(concatenador_2_data_out_72_) );
DFFPOSX1 DFFPOSX1_208 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf108), .D(concatenador_bloque_41_), .Q(concatenador_2_data_out_73_) );
DFFPOSX1 DFFPOSX1_209 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf107), .D(concatenador_bloque_42_), .Q(concatenador_2_data_out_74_) );
DFFPOSX1 DFFPOSX1_210 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(concatenador_bloque_43_), .Q(concatenador_2_data_out_75_) );
DFFPOSX1 DFFPOSX1_211 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(concatenador_bloque_44_), .Q(concatenador_2_data_out_76_) );
DFFPOSX1 DFFPOSX1_212 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(concatenador_bloque_45_), .Q(concatenador_2_data_out_77_) );
DFFPOSX1 DFFPOSX1_213 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(concatenador_bloque_46_), .Q(concatenador_2_data_out_78_) );
DFFPOSX1 DFFPOSX1_214 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(concatenador_bloque_47_), .Q(concatenador_2_data_out_79_) );
DFFPOSX1 DFFPOSX1_215 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(concatenador_bloque_48_), .Q(concatenador_2_data_out_80_) );
DFFPOSX1 DFFPOSX1_216 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(concatenador_bloque_49_), .Q(concatenador_2_data_out_81_) );
DFFPOSX1 DFFPOSX1_217 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(concatenador_bloque_50_), .Q(concatenador_2_data_out_82_) );
DFFPOSX1 DFFPOSX1_218 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(concatenador_bloque_51_), .Q(concatenador_2_data_out_83_) );
DFFPOSX1 DFFPOSX1_219 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(concatenador_bloque_52_), .Q(concatenador_2_data_out_84_) );
DFFPOSX1 DFFPOSX1_220 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(concatenador_bloque_53_), .Q(concatenador_2_data_out_85_) );
DFFPOSX1 DFFPOSX1_221 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(concatenador_bloque_54_), .Q(concatenador_2_data_out_86_) );
DFFPOSX1 DFFPOSX1_222 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(concatenador_bloque_55_), .Q(concatenador_2_data_out_87_) );
DFFPOSX1 DFFPOSX1_223 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(concatenador_bloque_56_), .Q(concatenador_2_data_out_88_) );
DFFPOSX1 DFFPOSX1_224 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(concatenador_bloque_57_), .Q(concatenador_2_data_out_89_) );
DFFPOSX1 DFFPOSX1_225 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(concatenador_bloque_58_), .Q(concatenador_2_data_out_90_) );
DFFPOSX1 DFFPOSX1_226 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(concatenador_bloque_59_), .Q(concatenador_2_data_out_91_) );
DFFPOSX1 DFFPOSX1_227 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(concatenador_bloque_60_), .Q(concatenador_2_data_out_92_) );
DFFPOSX1 DFFPOSX1_228 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(concatenador_bloque_61_), .Q(concatenador_2_data_out_93_) );
DFFPOSX1 DFFPOSX1_229 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(concatenador_bloque_62_), .Q(concatenador_2_data_out_94_) );
DFFPOSX1 DFFPOSX1_230 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(concatenador_bloque_63_), .Q(concatenador_2_data_out_95_) );
DFFPOSX1 DFFPOSX1_231 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(concatenador_bloque_64_), .Q(concatenador_2_data_out_96_) );
DFFPOSX1 DFFPOSX1_232 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(concatenador_bloque_65_), .Q(concatenador_2_data_out_97_) );
DFFPOSX1 DFFPOSX1_233 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(concatenador_bloque_66_), .Q(concatenador_2_data_out_98_) );
DFFPOSX1 DFFPOSX1_234 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(concatenador_bloque_67_), .Q(concatenador_2_data_out_99_) );
DFFPOSX1 DFFPOSX1_235 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(concatenador_bloque_68_), .Q(concatenador_2_data_out_100_) );
DFFPOSX1 DFFPOSX1_236 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(concatenador_bloque_69_), .Q(concatenador_2_data_out_101_) );
DFFPOSX1 DFFPOSX1_237 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(concatenador_bloque_70_), .Q(concatenador_2_data_out_102_) );
DFFPOSX1 DFFPOSX1_238 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(concatenador_bloque_71_), .Q(concatenador_2_data_out_103_) );
DFFPOSX1 DFFPOSX1_239 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(concatenador_bloque_72_), .Q(concatenador_2_data_out_104_) );
DFFPOSX1 DFFPOSX1_240 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(concatenador_bloque_73_), .Q(concatenador_2_data_out_105_) );
DFFPOSX1 DFFPOSX1_241 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(concatenador_bloque_74_), .Q(concatenador_2_data_out_106_) );
DFFPOSX1 DFFPOSX1_242 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(concatenador_bloque_75_), .Q(concatenador_2_data_out_107_) );
DFFPOSX1 DFFPOSX1_243 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(concatenador_bloque_76_), .Q(concatenador_2_data_out_108_) );
DFFPOSX1 DFFPOSX1_244 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(concatenador_bloque_77_), .Q(concatenador_2_data_out_109_) );
DFFPOSX1 DFFPOSX1_245 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(concatenador_bloque_78_), .Q(concatenador_2_data_out_110_) );
DFFPOSX1 DFFPOSX1_246 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(concatenador_bloque_79_), .Q(concatenador_2_data_out_111_) );
DFFPOSX1 DFFPOSX1_247 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(concatenador_bloque_80_), .Q(concatenador_2_data_out_112_) );
DFFPOSX1 DFFPOSX1_248 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(concatenador_bloque_81_), .Q(concatenador_2_data_out_113_) );
DFFPOSX1 DFFPOSX1_249 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(concatenador_bloque_82_), .Q(concatenador_2_data_out_114_) );
DFFPOSX1 DFFPOSX1_250 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(concatenador_bloque_83_), .Q(concatenador_2_data_out_115_) );
DFFPOSX1 DFFPOSX1_251 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(concatenador_bloque_84_), .Q(concatenador_2_data_out_116_) );
DFFPOSX1 DFFPOSX1_252 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(concatenador_bloque_85_), .Q(concatenador_2_data_out_117_) );
DFFPOSX1 DFFPOSX1_253 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(concatenador_bloque_86_), .Q(concatenador_2_data_out_118_) );
DFFPOSX1 DFFPOSX1_254 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(concatenador_bloque_87_), .Q(concatenador_2_data_out_119_) );
DFFPOSX1 DFFPOSX1_255 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(concatenador_bloque_88_), .Q(concatenador_2_data_out_120_) );
DFFPOSX1 DFFPOSX1_256 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(concatenador_bloque_89_), .Q(concatenador_2_data_out_121_) );
DFFPOSX1 DFFPOSX1_257 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(concatenador_bloque_90_), .Q(concatenador_2_data_out_122_) );
DFFPOSX1 DFFPOSX1_258 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(concatenador_bloque_91_), .Q(concatenador_2_data_out_123_) );
DFFPOSX1 DFFPOSX1_259 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(concatenador_bloque_92_), .Q(concatenador_2_data_out_124_) );
DFFPOSX1 DFFPOSX1_260 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(concatenador_bloque_93_), .Q(concatenador_2_data_out_125_) );
DFFPOSX1 DFFPOSX1_261 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(concatenador_bloque_94_), .Q(concatenador_2_data_out_126_) );
DFFPOSX1 DFFPOSX1_262 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(concatenador_bloque_95_), .Q(concatenador_2_data_out_127_) );
DFFPOSX1 DFFPOSX1_263 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(concatenador_3_nonce_0_), .Q(concatenador_3_data_out_0_) );
DFFPOSX1 DFFPOSX1_264 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(concatenador_3_nonce_1_), .Q(concatenador_3_data_out_1_) );
DFFPOSX1 DFFPOSX1_265 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(concatenador_3_nonce_2_), .Q(concatenador_3_data_out_2_) );
DFFPOSX1 DFFPOSX1_266 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(concatenador_3_nonce_3_), .Q(concatenador_3_data_out_3_) );
DFFPOSX1 DFFPOSX1_267 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(concatenador_3_nonce_4_), .Q(concatenador_3_data_out_4_) );
DFFPOSX1 DFFPOSX1_268 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(concatenador_3_nonce_5_), .Q(concatenador_3_data_out_5_) );
DFFPOSX1 DFFPOSX1_269 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(concatenador_3_nonce_6_), .Q(concatenador_3_data_out_6_) );
DFFPOSX1 DFFPOSX1_270 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(concatenador_3_nonce_7_), .Q(concatenador_3_data_out_7_) );
DFFPOSX1 DFFPOSX1_271 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(concatenador_3_nonce_8_), .Q(concatenador_3_data_out_8_) );
DFFPOSX1 DFFPOSX1_272 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(concatenador_3_nonce_9_), .Q(concatenador_3_data_out_9_) );
DFFPOSX1 DFFPOSX1_273 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(concatenador_3_nonce_10_), .Q(concatenador_3_data_out_10_) );
DFFPOSX1 DFFPOSX1_274 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(concatenador_3_nonce_11_), .Q(concatenador_3_data_out_11_) );
DFFPOSX1 DFFPOSX1_275 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(concatenador_3_nonce_12_), .Q(concatenador_3_data_out_12_) );
DFFPOSX1 DFFPOSX1_276 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(concatenador_3_nonce_13_), .Q(concatenador_3_data_out_13_) );
DFFPOSX1 DFFPOSX1_277 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(concatenador_3_nonce_14_), .Q(concatenador_3_data_out_14_) );
DFFPOSX1 DFFPOSX1_278 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(concatenador_3_nonce_15_), .Q(concatenador_3_data_out_15_) );
DFFPOSX1 DFFPOSX1_279 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(concatenador_3_nonce_16_), .Q(concatenador_3_data_out_16_) );
DFFPOSX1 DFFPOSX1_280 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(concatenador_3_nonce_17_), .Q(concatenador_3_data_out_17_) );
DFFPOSX1 DFFPOSX1_281 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(concatenador_3_nonce_18_), .Q(concatenador_3_data_out_18_) );
DFFPOSX1 DFFPOSX1_282 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(concatenador_3_nonce_19_), .Q(concatenador_3_data_out_19_) );
DFFPOSX1 DFFPOSX1_283 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(concatenador_3_nonce_20_), .Q(concatenador_3_data_out_20_) );
DFFPOSX1 DFFPOSX1_284 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(concatenador_3_nonce_21_), .Q(concatenador_3_data_out_21_) );
DFFPOSX1 DFFPOSX1_285 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(concatenador_3_nonce_22_), .Q(concatenador_3_data_out_22_) );
DFFPOSX1 DFFPOSX1_286 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(concatenador_3_nonce_23_), .Q(concatenador_3_data_out_23_) );
DFFPOSX1 DFFPOSX1_287 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(concatenador_3_nonce_24_), .Q(concatenador_3_data_out_24_) );
DFFPOSX1 DFFPOSX1_288 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(concatenador_3_nonce_25_), .Q(concatenador_3_data_out_25_) );
DFFPOSX1 DFFPOSX1_289 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(concatenador_3_nonce_26_), .Q(concatenador_3_data_out_26_) );
DFFPOSX1 DFFPOSX1_290 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(concatenador_3_nonce_27_), .Q(concatenador_3_data_out_27_) );
DFFPOSX1 DFFPOSX1_291 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(concatenador_3_nonce_28_), .Q(concatenador_3_data_out_28_) );
DFFPOSX1 DFFPOSX1_292 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(concatenador_3_nonce_29_), .Q(concatenador_3_data_out_29_) );
DFFPOSX1 DFFPOSX1_293 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(concatenador_3_nonce_30_), .Q(concatenador_3_data_out_30_) );
DFFPOSX1 DFFPOSX1_294 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(concatenador_3_nonce_31_), .Q(concatenador_3_data_out_31_) );
DFFPOSX1 DFFPOSX1_295 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(concatenador_bloque_0_), .Q(concatenador_3_data_out_32_) );
DFFPOSX1 DFFPOSX1_296 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(concatenador_bloque_1_), .Q(concatenador_3_data_out_33_) );
DFFPOSX1 DFFPOSX1_297 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(concatenador_bloque_2_), .Q(concatenador_3_data_out_34_) );
DFFPOSX1 DFFPOSX1_298 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(concatenador_bloque_3_), .Q(concatenador_3_data_out_35_) );
DFFPOSX1 DFFPOSX1_299 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(concatenador_bloque_4_), .Q(concatenador_3_data_out_36_) );
DFFPOSX1 DFFPOSX1_300 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(concatenador_bloque_5_), .Q(concatenador_3_data_out_37_) );
DFFPOSX1 DFFPOSX1_301 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(concatenador_bloque_6_), .Q(concatenador_3_data_out_38_) );
DFFPOSX1 DFFPOSX1_302 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(concatenador_bloque_7_), .Q(concatenador_3_data_out_39_) );
DFFPOSX1 DFFPOSX1_303 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(concatenador_bloque_8_), .Q(concatenador_3_data_out_40_) );
DFFPOSX1 DFFPOSX1_304 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(concatenador_bloque_9_), .Q(concatenador_3_data_out_41_) );
DFFPOSX1 DFFPOSX1_305 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(concatenador_bloque_10_), .Q(concatenador_3_data_out_42_) );
DFFPOSX1 DFFPOSX1_306 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(concatenador_bloque_11_), .Q(concatenador_3_data_out_43_) );
DFFPOSX1 DFFPOSX1_307 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(concatenador_bloque_12_), .Q(concatenador_3_data_out_44_) );
DFFPOSX1 DFFPOSX1_308 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(concatenador_bloque_13_), .Q(concatenador_3_data_out_45_) );
DFFPOSX1 DFFPOSX1_309 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(concatenador_bloque_14_), .Q(concatenador_3_data_out_46_) );
DFFPOSX1 DFFPOSX1_310 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(concatenador_bloque_15_), .Q(concatenador_3_data_out_47_) );
DFFPOSX1 DFFPOSX1_311 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(concatenador_bloque_16_), .Q(concatenador_3_data_out_48_) );
DFFPOSX1 DFFPOSX1_312 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(concatenador_bloque_17_), .Q(concatenador_3_data_out_49_) );
DFFPOSX1 DFFPOSX1_313 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(concatenador_bloque_18_), .Q(concatenador_3_data_out_50_) );
DFFPOSX1 DFFPOSX1_314 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(concatenador_bloque_19_), .Q(concatenador_3_data_out_51_) );
DFFPOSX1 DFFPOSX1_315 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(concatenador_bloque_20_), .Q(concatenador_3_data_out_52_) );
DFFPOSX1 DFFPOSX1_316 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(concatenador_bloque_21_), .Q(concatenador_3_data_out_53_) );
DFFPOSX1 DFFPOSX1_317 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf157), .D(concatenador_bloque_22_), .Q(concatenador_3_data_out_54_) );
DFFPOSX1 DFFPOSX1_318 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf156), .D(concatenador_bloque_23_), .Q(concatenador_3_data_out_55_) );
DFFPOSX1 DFFPOSX1_319 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf155), .D(concatenador_bloque_24_), .Q(concatenador_3_data_out_56_) );
DFFPOSX1 DFFPOSX1_320 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf154), .D(concatenador_bloque_25_), .Q(concatenador_3_data_out_57_) );
DFFPOSX1 DFFPOSX1_321 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf153), .D(concatenador_bloque_26_), .Q(concatenador_3_data_out_58_) );
DFFPOSX1 DFFPOSX1_322 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf152), .D(concatenador_bloque_27_), .Q(concatenador_3_data_out_59_) );
DFFPOSX1 DFFPOSX1_323 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf151), .D(concatenador_bloque_28_), .Q(concatenador_3_data_out_60_) );
DFFPOSX1 DFFPOSX1_324 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf150), .D(concatenador_bloque_29_), .Q(concatenador_3_data_out_61_) );
DFFPOSX1 DFFPOSX1_325 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf149), .D(concatenador_bloque_30_), .Q(concatenador_3_data_out_62_) );
DFFPOSX1 DFFPOSX1_326 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf148), .D(concatenador_bloque_31_), .Q(concatenador_3_data_out_63_) );
DFFPOSX1 DFFPOSX1_327 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf147), .D(concatenador_bloque_32_), .Q(concatenador_3_data_out_64_) );
DFFPOSX1 DFFPOSX1_328 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf146), .D(concatenador_bloque_33_), .Q(concatenador_3_data_out_65_) );
DFFPOSX1 DFFPOSX1_329 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf145), .D(concatenador_bloque_34_), .Q(concatenador_3_data_out_66_) );
DFFPOSX1 DFFPOSX1_330 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf144), .D(concatenador_bloque_35_), .Q(concatenador_3_data_out_67_) );
DFFPOSX1 DFFPOSX1_331 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf143), .D(concatenador_bloque_36_), .Q(concatenador_3_data_out_68_) );
DFFPOSX1 DFFPOSX1_332 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf142), .D(concatenador_bloque_37_), .Q(concatenador_3_data_out_69_) );
DFFPOSX1 DFFPOSX1_333 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf141), .D(concatenador_bloque_38_), .Q(concatenador_3_data_out_70_) );
DFFPOSX1 DFFPOSX1_334 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf140), .D(concatenador_bloque_39_), .Q(concatenador_3_data_out_71_) );
DFFPOSX1 DFFPOSX1_335 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf139), .D(concatenador_bloque_40_), .Q(concatenador_3_data_out_72_) );
DFFPOSX1 DFFPOSX1_336 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf138), .D(concatenador_bloque_41_), .Q(concatenador_3_data_out_73_) );
DFFPOSX1 DFFPOSX1_337 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf137), .D(concatenador_bloque_42_), .Q(concatenador_3_data_out_74_) );
DFFPOSX1 DFFPOSX1_338 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf136), .D(concatenador_bloque_43_), .Q(concatenador_3_data_out_75_) );
DFFPOSX1 DFFPOSX1_339 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf135), .D(concatenador_bloque_44_), .Q(concatenador_3_data_out_76_) );
DFFPOSX1 DFFPOSX1_340 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf134), .D(concatenador_bloque_45_), .Q(concatenador_3_data_out_77_) );
DFFPOSX1 DFFPOSX1_341 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf133), .D(concatenador_bloque_46_), .Q(concatenador_3_data_out_78_) );
DFFPOSX1 DFFPOSX1_342 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf132), .D(concatenador_bloque_47_), .Q(concatenador_3_data_out_79_) );
DFFPOSX1 DFFPOSX1_343 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf131), .D(concatenador_bloque_48_), .Q(concatenador_3_data_out_80_) );
DFFPOSX1 DFFPOSX1_344 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf130), .D(concatenador_bloque_49_), .Q(concatenador_3_data_out_81_) );
DFFPOSX1 DFFPOSX1_345 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf129), .D(concatenador_bloque_50_), .Q(concatenador_3_data_out_82_) );
DFFPOSX1 DFFPOSX1_346 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf128), .D(concatenador_bloque_51_), .Q(concatenador_3_data_out_83_) );
DFFPOSX1 DFFPOSX1_347 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf127), .D(concatenador_bloque_52_), .Q(concatenador_3_data_out_84_) );
DFFPOSX1 DFFPOSX1_348 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf126), .D(concatenador_bloque_53_), .Q(concatenador_3_data_out_85_) );
DFFPOSX1 DFFPOSX1_349 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf125), .D(concatenador_bloque_54_), .Q(concatenador_3_data_out_86_) );
DFFPOSX1 DFFPOSX1_350 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf124), .D(concatenador_bloque_55_), .Q(concatenador_3_data_out_87_) );
DFFPOSX1 DFFPOSX1_351 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf123), .D(concatenador_bloque_56_), .Q(concatenador_3_data_out_88_) );
DFFPOSX1 DFFPOSX1_352 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf122), .D(concatenador_bloque_57_), .Q(concatenador_3_data_out_89_) );
DFFPOSX1 DFFPOSX1_353 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf121), .D(concatenador_bloque_58_), .Q(concatenador_3_data_out_90_) );
DFFPOSX1 DFFPOSX1_354 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf120), .D(concatenador_bloque_59_), .Q(concatenador_3_data_out_91_) );
DFFPOSX1 DFFPOSX1_355 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf119), .D(concatenador_bloque_60_), .Q(concatenador_3_data_out_92_) );
DFFPOSX1 DFFPOSX1_356 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf118), .D(concatenador_bloque_61_), .Q(concatenador_3_data_out_93_) );
DFFPOSX1 DFFPOSX1_357 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf117), .D(concatenador_bloque_62_), .Q(concatenador_3_data_out_94_) );
DFFPOSX1 DFFPOSX1_358 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf116), .D(concatenador_bloque_63_), .Q(concatenador_3_data_out_95_) );
DFFPOSX1 DFFPOSX1_359 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf115), .D(concatenador_bloque_64_), .Q(concatenador_3_data_out_96_) );
DFFPOSX1 DFFPOSX1_360 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf114), .D(concatenador_bloque_65_), .Q(concatenador_3_data_out_97_) );
DFFPOSX1 DFFPOSX1_361 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf113), .D(concatenador_bloque_66_), .Q(concatenador_3_data_out_98_) );
DFFPOSX1 DFFPOSX1_362 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf112), .D(concatenador_bloque_67_), .Q(concatenador_3_data_out_99_) );
DFFPOSX1 DFFPOSX1_363 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf111), .D(concatenador_bloque_68_), .Q(concatenador_3_data_out_100_) );
DFFPOSX1 DFFPOSX1_364 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf110), .D(concatenador_bloque_69_), .Q(concatenador_3_data_out_101_) );
DFFPOSX1 DFFPOSX1_365 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf109), .D(concatenador_bloque_70_), .Q(concatenador_3_data_out_102_) );
DFFPOSX1 DFFPOSX1_366 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf108), .D(concatenador_bloque_71_), .Q(concatenador_3_data_out_103_) );
DFFPOSX1 DFFPOSX1_367 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf107), .D(concatenador_bloque_72_), .Q(concatenador_3_data_out_104_) );
DFFPOSX1 DFFPOSX1_368 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(concatenador_bloque_73_), .Q(concatenador_3_data_out_105_) );
DFFPOSX1 DFFPOSX1_369 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(concatenador_bloque_74_), .Q(concatenador_3_data_out_106_) );
DFFPOSX1 DFFPOSX1_370 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(concatenador_bloque_75_), .Q(concatenador_3_data_out_107_) );
DFFPOSX1 DFFPOSX1_371 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(concatenador_bloque_76_), .Q(concatenador_3_data_out_108_) );
DFFPOSX1 DFFPOSX1_372 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(concatenador_bloque_77_), .Q(concatenador_3_data_out_109_) );
DFFPOSX1 DFFPOSX1_373 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(concatenador_bloque_78_), .Q(concatenador_3_data_out_110_) );
DFFPOSX1 DFFPOSX1_374 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(concatenador_bloque_79_), .Q(concatenador_3_data_out_111_) );
DFFPOSX1 DFFPOSX1_375 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(concatenador_bloque_80_), .Q(concatenador_3_data_out_112_) );
DFFPOSX1 DFFPOSX1_376 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(concatenador_bloque_81_), .Q(concatenador_3_data_out_113_) );
DFFPOSX1 DFFPOSX1_377 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(concatenador_bloque_82_), .Q(concatenador_3_data_out_114_) );
DFFPOSX1 DFFPOSX1_378 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(concatenador_bloque_83_), .Q(concatenador_3_data_out_115_) );
DFFPOSX1 DFFPOSX1_379 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(concatenador_bloque_84_), .Q(concatenador_3_data_out_116_) );
DFFPOSX1 DFFPOSX1_380 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(concatenador_bloque_85_), .Q(concatenador_3_data_out_117_) );
DFFPOSX1 DFFPOSX1_381 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(concatenador_bloque_86_), .Q(concatenador_3_data_out_118_) );
DFFPOSX1 DFFPOSX1_382 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(concatenador_bloque_87_), .Q(concatenador_3_data_out_119_) );
DFFPOSX1 DFFPOSX1_383 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(concatenador_bloque_88_), .Q(concatenador_3_data_out_120_) );
DFFPOSX1 DFFPOSX1_384 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(concatenador_bloque_89_), .Q(concatenador_3_data_out_121_) );
DFFPOSX1 DFFPOSX1_385 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(concatenador_bloque_90_), .Q(concatenador_3_data_out_122_) );
DFFPOSX1 DFFPOSX1_386 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(concatenador_bloque_91_), .Q(concatenador_3_data_out_123_) );
DFFPOSX1 DFFPOSX1_387 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(concatenador_bloque_92_), .Q(concatenador_3_data_out_124_) );
DFFPOSX1 DFFPOSX1_388 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(concatenador_bloque_93_), .Q(concatenador_3_data_out_125_) );
DFFPOSX1 DFFPOSX1_389 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(concatenador_bloque_94_), .Q(concatenador_3_data_out_126_) );
DFFPOSX1 DFFPOSX1_390 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(concatenador_bloque_95_), .Q(concatenador_3_data_out_127_) );
INVX1 INVX1_46 ( .gnd(gnd), .vdd(vdd), .A(_0__bF_buf8), .Y(_4418_) );
NAND2X1 NAND2X1_58 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf7), .B(_4418_), .Y(_4419_) );
NOR2X1 NOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(comparador_next_bF_buf3), .B(_4419_), .Y(_302_) );
NOR2X1 NOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe70_bF_buf3), .B(micro_hash_ucr_pipe5), .Y(_4420_) );
NAND2X1 NAND2X1_59 ( .gnd(gnd), .vdd(vdd), .A(H_16_), .B(_4420_), .Y(_4421_) );
INVX1 INVX1_47 ( .gnd(gnd), .vdd(vdd), .A(H_16_), .Y(_4422_) );
INVX8 INVX8_1 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_0_bF_buf3_), .Y(_4423_) );
OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_4422_), .B(_4423__bF_buf3), .C(micro_hash_ucr_pipe70_bF_buf2), .Y(_4424_) );
OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(H_16_), .B(micro_hash_ucr_c_0_bF_buf2_), .C(_302__bF_buf13), .Y(_4425_) );
AOI21X1 AOI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_4421_), .B(_4424_), .C(_4425_), .Y(_300__16_) );
NOR2X1 NOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(_4422_), .B(_4423__bF_buf2), .Y(_4426_) );
NOR2X1 NOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(H_17_), .B(micro_hash_ucr_c_1_bF_buf3_), .Y(_4427_) );
NAND2X1 NAND2X1_60 ( .gnd(gnd), .vdd(vdd), .A(H_17_), .B(micro_hash_ucr_c_1_bF_buf2_), .Y(_4428_) );
INVX1 INVX1_48 ( .gnd(gnd), .vdd(vdd), .A(_4428_), .Y(_4429_) );
NOR2X1 NOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_4427_), .B(_4429_), .Y(_4430_) );
XNOR2X1 XNOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_4430_), .B(_4426_), .Y(_4431_) );
INVX8 INVX8_2 ( .gnd(gnd), .vdd(vdd), .A(_4420_), .Y(_4432_) );
OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(H_17_), .B(_4432_), .C(_302__bF_buf12), .Y(_4433_) );
AOI21X1 AOI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe70_bF_buf1), .B(_4431_), .C(_4433_), .Y(_300__17_) );
INVX1 INVX1_49 ( .gnd(gnd), .vdd(vdd), .A(_4426_), .Y(_4434_) );
OAI21X1 OAI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_4434_), .B(_4427_), .C(_4428_), .Y(_4435_) );
XOR2X1 XOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(H_18_), .B(micro_hash_ucr_c_2_bF_buf3_), .Y(_4436_) );
XNOR2X1 XNOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_4435_), .B(_4436_), .Y(_4437_) );
OAI21X1 OAI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(H_18_), .B(_4432_), .C(_302__bF_buf11), .Y(_4438_) );
AOI21X1 AOI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe70_bF_buf0), .B(_4437_), .C(_4438_), .Y(_300__18_) );
INVX1 INVX1_50 ( .gnd(gnd), .vdd(vdd), .A(_4435_), .Y(_4439_) );
INVX1 INVX1_51 ( .gnd(gnd), .vdd(vdd), .A(_4436_), .Y(_4440_) );
NOR2X1 NOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_4440_), .B(_4439_), .Y(_4441_) );
AOI21X1 AOI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(H_18_), .B(micro_hash_ucr_c_2_bF_buf2_), .C(_4441_), .Y(_4442_) );
NOR2X1 NOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(H_19_), .B(micro_hash_ucr_c_3_bF_buf4_), .Y(_4443_) );
INVX1 INVX1_52 ( .gnd(gnd), .vdd(vdd), .A(H_19_), .Y(_4444_) );
INVX4 INVX4_1 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_3_bF_buf3_), .Y(_4445_) );
NOR2X1 NOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_4444_), .B(_4445_), .Y(_4446_) );
OR2X2 OR2X2_22 ( .gnd(gnd), .vdd(vdd), .A(_4446_), .B(_4443_), .Y(_4447_) );
XNOR2X1 XNOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_4442_), .B(_4447_), .Y(_4448_) );
OAI21X1 OAI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(H_19_), .B(_4432_), .C(_302__bF_buf10), .Y(_4449_) );
AOI21X1 AOI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe70_bF_buf3), .B(_4448_), .C(_4449_), .Y(_300__19_) );
NOR2X1 NOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(H_20_), .B(micro_hash_ucr_c_4_), .Y(_4450_) );
AND2X2 AND2X2_7 ( .gnd(gnd), .vdd(vdd), .A(H_20_), .B(micro_hash_ucr_c_4_), .Y(_4451_) );
NOR2X1 NOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_4450_), .B(_4451_), .Y(_4452_) );
INVX1 INVX1_53 ( .gnd(gnd), .vdd(vdd), .A(_4446_), .Y(_4453_) );
OAI21X1 OAI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_4442_), .B(_4443_), .C(_4453_), .Y(_4454_) );
XNOR2X1 XNOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_4454_), .B(_4452_), .Y(_4455_) );
OAI21X1 OAI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(H_20_), .B(_4432_), .C(_302__bF_buf9), .Y(_4456_) );
AOI21X1 AOI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe70_bF_buf2), .B(_4455_), .C(_4456_), .Y(_300__20_) );
AOI21X1 AOI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_4452_), .B(_4454_), .C(_4451_), .Y(_4457_) );
NOR2X1 NOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(H_21_), .B(micro_hash_ucr_c_5_), .Y(_4458_) );
INVX1 INVX1_54 ( .gnd(gnd), .vdd(vdd), .A(H_21_), .Y(_4459_) );
INVX2 INVX2_13 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_5_), .Y(_4460_) );
NOR2X1 NOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_4459_), .B(_4460_), .Y(_4461_) );
NOR2X1 NOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_4458_), .B(_4461_), .Y(_4462_) );
OAI21X1 OAI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_4457_), .B(_4462_), .C(micro_hash_ucr_pipe70_bF_buf1), .Y(_4463_) );
AOI21X1 AOI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(_4457_), .B(_4462_), .C(_4463_), .Y(_4464_) );
OAI21X1 OAI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(H_21_), .B(_4432_), .C(_302__bF_buf8), .Y(_4465_) );
NOR2X1 NOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_4465_), .B(_4464_), .Y(_300__21_) );
XOR2X1 XOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(H_22_), .B(micro_hash_ucr_c_6_), .Y(_4466_) );
INVX1 INVX1_55 ( .gnd(gnd), .vdd(vdd), .A(_4461_), .Y(_4467_) );
OAI21X1 OAI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(_4457_), .B(_4458_), .C(_4467_), .Y(_4468_) );
XNOR2X1 XNOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_4468_), .B(_4466_), .Y(_4469_) );
OAI21X1 OAI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(H_22_), .B(_4432_), .C(_302__bF_buf7), .Y(_4470_) );
AOI21X1 AOI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe70_bF_buf0), .B(_4469_), .C(_4470_), .Y(_300__22_) );
INVX1 INVX1_56 ( .gnd(gnd), .vdd(vdd), .A(H_22_), .Y(_4471_) );
INVX2 INVX2_14 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_6_), .Y(_4472_) );
NAND2X1 NAND2X1_61 ( .gnd(gnd), .vdd(vdd), .A(_4466_), .B(_4468_), .Y(_4473_) );
OAI21X1 OAI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_4471_), .B(_4472_), .C(_4473_), .Y(_4474_) );
XOR2X1 XOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(H_23_), .B(micro_hash_ucr_c_7_), .Y(_4475_) );
XNOR2X1 XNOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_4474_), .B(_4475_), .Y(_4476_) );
OAI21X1 OAI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(H_23_), .B(_4432_), .C(_302__bF_buf6), .Y(_4477_) );
AOI21X1 AOI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe70_bF_buf3), .B(_4476_), .C(_4477_), .Y(_300__23_) );
INVX2 INVX2_15 ( .gnd(gnd), .vdd(vdd), .A(H_8_), .Y(_4478_) );
INVX8 INVX8_3 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe70_bF_buf2), .Y(_4479_) );
OAI21X1 OAI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_4479__bF_buf3), .B(micro_hash_ucr_b_0_bF_buf3_), .C(_4432_), .Y(_4480_) );
INVX8 INVX8_4 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_0_bF_buf2_), .Y(_4481_) );
NOR2X1 NOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(_4478_), .B(_4481_), .Y(_4482_) );
INVX1 INVX1_57 ( .gnd(gnd), .vdd(vdd), .A(_4482_), .Y(_4483_) );
OAI21X1 OAI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_4483_), .B(_4479__bF_buf2), .C(_302__bF_buf5), .Y(_4484_) );
AOI21X1 AOI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_4478_), .B(_4480_), .C(_4484_), .Y(_300__8_) );
INVX2 INVX2_16 ( .gnd(gnd), .vdd(vdd), .A(H_9_), .Y(_4485_) );
NOR2X1 NOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(H_9_), .B(micro_hash_ucr_b_1_bF_buf3_), .Y(_4486_) );
INVX8 INVX8_5 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_1_bF_buf2_), .Y(_4487_) );
NOR2X1 NOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(_4485_), .B(_4487_), .Y(_4488_) );
NOR2X1 NOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_4486_), .B(_4488_), .Y(_4489_) );
AOI21X1 AOI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_4482_), .B(_4489_), .C(_4479__bF_buf1), .Y(_376_) );
OAI21X1 OAI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_4482_), .B(_4489_), .C(_376_), .Y(_377_) );
OAI21X1 OAI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_4485_), .B(_4432_), .C(_377_), .Y(_378_) );
AND2X2 AND2X2_8 ( .gnd(gnd), .vdd(vdd), .A(_378_), .B(_302__bF_buf4), .Y(_300__9_) );
INVX2 INVX2_17 ( .gnd(gnd), .vdd(vdd), .A(H_10_), .Y(_379_) );
INVX1 INVX1_58 ( .gnd(gnd), .vdd(vdd), .A(_4488_), .Y(_380_) );
OAI21X1 OAI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_4483_), .B(_4486_), .C(_380_), .Y(_381_) );
XOR2X1 XOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(H_10_), .B(micro_hash_ucr_b_2_bF_buf3_), .Y(_382_) );
INVX1 INVX1_59 ( .gnd(gnd), .vdd(vdd), .A(_381_), .Y(_383_) );
INVX1 INVX1_60 ( .gnd(gnd), .vdd(vdd), .A(_382_), .Y(_384_) );
NOR2X1 NOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(_384_), .B(_383_), .Y(_385_) );
NOR2X1 NOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(_4479__bF_buf0), .B(_385_), .Y(_386_) );
OAI21X1 OAI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(_381_), .B(_382_), .C(_386_), .Y(_387_) );
OAI21X1 OAI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(_379_), .B(_4432_), .C(_387_), .Y(_388_) );
AND2X2 AND2X2_9 ( .gnd(gnd), .vdd(vdd), .A(_388_), .B(_302__bF_buf3), .Y(_300__10_) );
INVX8 INVX8_6 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_2_bF_buf2_), .Y(_389_) );
INVX1 INVX1_61 ( .gnd(gnd), .vdd(vdd), .A(_385_), .Y(_390_) );
OAI21X1 OAI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(_379_), .B(_389_), .C(_390_), .Y(_391_) );
NOR2X1 NOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(H_11_), .B(micro_hash_ucr_b_3_bF_buf3_), .Y(_392_) );
INVX1 INVX1_62 ( .gnd(gnd), .vdd(vdd), .A(H_11_), .Y(_393_) );
INVX8 INVX8_7 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_3_bF_buf2_), .Y(_394_) );
NOR2X1 NOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_393_), .B(_394_), .Y(_395_) );
OR2X2 OR2X2_23 ( .gnd(gnd), .vdd(vdd), .A(_395_), .B(_392_), .Y(_396_) );
OAI21X1 OAI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_391_), .B(_396_), .C(micro_hash_ucr_pipe70_bF_buf1), .Y(_397_) );
AOI21X1 AOI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_391_), .B(_396_), .C(_397_), .Y(_398_) );
OAI21X1 OAI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(H_11_), .B(_4432_), .C(_302__bF_buf2), .Y(_399_) );
NOR2X1 NOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(_399_), .B(_398_), .Y(_300__11_) );
INVX8 INVX8_8 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf1), .Y(_400_) );
XOR2X1 XOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(H_12_), .B(micro_hash_ucr_b_4_bF_buf3_), .Y(_401_) );
INVX1 INVX1_63 ( .gnd(gnd), .vdd(vdd), .A(_392_), .Y(_402_) );
AOI21X1 AOI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_402_), .B(_391_), .C(_395_), .Y(_403_) );
XNOR2X1 XNOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_403_), .B(_401_), .Y(_404_) );
INVX1 INVX1_64 ( .gnd(gnd), .vdd(vdd), .A(H_12_), .Y(_405_) );
OAI21X1 OAI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(_405_), .B(micro_hash_ucr_pipe5), .C(_4479__bF_buf3), .Y(_406_) );
OAI21X1 OAI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(_404_), .B(_4479__bF_buf2), .C(_406_), .Y(_407_) );
NOR2X1 NOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(_400__bF_buf12), .B(_407_), .Y(_300__12_) );
NAND2X1 NAND2X1_62 ( .gnd(gnd), .vdd(vdd), .A(H_12_), .B(micro_hash_ucr_b_4_bF_buf2_), .Y(_408_) );
INVX1 INVX1_65 ( .gnd(gnd), .vdd(vdd), .A(_401_), .Y(_409_) );
OAI21X1 OAI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(_403_), .B(_409_), .C(_408_), .Y(_410_) );
INVX2 INVX2_18 ( .gnd(gnd), .vdd(vdd), .A(_410_), .Y(_411_) );
NOR2X1 NOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(H_13_), .B(micro_hash_ucr_b_5_bF_buf3_), .Y(_412_) );
INVX1 INVX1_66 ( .gnd(gnd), .vdd(vdd), .A(H_13_), .Y(_413_) );
INVX8 INVX8_9 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_5_bF_buf2_), .Y(_414_) );
NOR2X1 NOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(_413_), .B(_414__bF_buf3), .Y(_415_) );
NOR2X1 NOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(_412_), .B(_415_), .Y(_416_) );
AND2X2 AND2X2_10 ( .gnd(gnd), .vdd(vdd), .A(_411_), .B(_416_), .Y(_417_) );
OAI21X1 OAI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(_411_), .B(_416_), .C(micro_hash_ucr_pipe70_bF_buf0), .Y(_418_) );
OAI21X1 OAI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(_413_), .B(micro_hash_ucr_pipe5), .C(_4479__bF_buf1), .Y(_419_) );
OAI21X1 OAI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(_417_), .B(_418_), .C(_419_), .Y(_420_) );
NOR2X1 NOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(_400__bF_buf11), .B(_420_), .Y(_300__13_) );
XOR2X1 XOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(H_14_), .B(micro_hash_ucr_b_6_bF_buf3_), .Y(_421_) );
INVX1 INVX1_67 ( .gnd(gnd), .vdd(vdd), .A(_415_), .Y(_422_) );
OAI21X1 OAI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(_411_), .B(_412_), .C(_422_), .Y(_423_) );
XNOR2X1 XNOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_423_), .B(_421_), .Y(_424_) );
INVX2 INVX2_19 ( .gnd(gnd), .vdd(vdd), .A(H_14_), .Y(_425_) );
OAI21X1 OAI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(_425_), .B(micro_hash_ucr_pipe5), .C(_4479__bF_buf0), .Y(_426_) );
NAND2X1 NAND2X1_63 ( .gnd(gnd), .vdd(vdd), .A(_426_), .B(_302__bF_buf0), .Y(_427_) );
AOI21X1 AOI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe70_bF_buf3), .B(_424_), .C(_427_), .Y(_300__14_) );
INVX8 INVX8_10 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_6_bF_buf2_), .Y(_428_) );
NAND2X1 NAND2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_421_), .B(_423_), .Y(_429_) );
OAI21X1 OAI21X1_66 ( .gnd(gnd), .vdd(vdd), .A(_425_), .B(_428__bF_buf3), .C(_429_), .Y(_430_) );
XOR2X1 XOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(H_15_), .B(micro_hash_ucr_b_7_), .Y(_431_) );
XNOR2X1 XNOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_430_), .B(_431_), .Y(_432_) );
OAI21X1 OAI21X1_67 ( .gnd(gnd), .vdd(vdd), .A(H_15_), .B(_4432_), .C(_302__bF_buf13), .Y(_433_) );
AOI21X1 AOI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe70_bF_buf2), .B(_432_), .C(_433_), .Y(_300__15_) );
INVX2 INVX2_20 ( .gnd(gnd), .vdd(vdd), .A(H_0_), .Y(_434_) );
OAI21X1 OAI21X1_68 ( .gnd(gnd), .vdd(vdd), .A(_4479__bF_buf3), .B(micro_hash_ucr_a_0_bF_buf3_), .C(_4432_), .Y(_435_) );
INVX4 INVX4_2 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_0_bF_buf2_), .Y(_436_) );
NOR2X1 NOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(_434_), .B(_436_), .Y(_437_) );
INVX1 INVX1_68 ( .gnd(gnd), .vdd(vdd), .A(_437_), .Y(_438_) );
OAI21X1 OAI21X1_69 ( .gnd(gnd), .vdd(vdd), .A(_438_), .B(_4479__bF_buf2), .C(_302__bF_buf12), .Y(_439_) );
AOI21X1 AOI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(_434_), .B(_435_), .C(_439_), .Y(_300__0_) );
INVX1 INVX1_69 ( .gnd(gnd), .vdd(vdd), .A(H_1_), .Y(_440_) );
NOR2X1 NOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(H_1_), .B(micro_hash_ucr_a_1_), .Y(_441_) );
INVX8 INVX8_11 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_1_), .Y(_442_) );
NOR2X1 NOR2X1_61 ( .gnd(gnd), .vdd(vdd), .A(_440_), .B(_442_), .Y(_443_) );
NOR2X1 NOR2X1_62 ( .gnd(gnd), .vdd(vdd), .A(_441_), .B(_443_), .Y(_444_) );
AOI21X1 AOI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(_437_), .B(_444_), .C(_4479__bF_buf1), .Y(_445_) );
OAI21X1 OAI21X1_70 ( .gnd(gnd), .vdd(vdd), .A(_437_), .B(_444_), .C(_445_), .Y(_446_) );
OAI21X1 OAI21X1_71 ( .gnd(gnd), .vdd(vdd), .A(_440_), .B(_4432_), .C(_446_), .Y(_447_) );
AND2X2 AND2X2_11 ( .gnd(gnd), .vdd(vdd), .A(_447_), .B(_302__bF_buf11), .Y(_300__1_) );
INVX1 INVX1_70 ( .gnd(gnd), .vdd(vdd), .A(_443_), .Y(_448_) );
OAI21X1 OAI21X1_72 ( .gnd(gnd), .vdd(vdd), .A(_438_), .B(_441_), .C(_448_), .Y(_449_) );
XOR2X1 XOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(H_2_), .B(micro_hash_ucr_a_2_), .Y(_450_) );
INVX1 INVX1_71 ( .gnd(gnd), .vdd(vdd), .A(_449_), .Y(_451_) );
INVX1 INVX1_72 ( .gnd(gnd), .vdd(vdd), .A(_450_), .Y(_452_) );
NOR2X1 NOR2X1_63 ( .gnd(gnd), .vdd(vdd), .A(_452_), .B(_451_), .Y(_453_) );
NOR2X1 NOR2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_4479__bF_buf0), .B(_453_), .Y(_454_) );
OAI21X1 OAI21X1_73 ( .gnd(gnd), .vdd(vdd), .A(_449_), .B(_450_), .C(_454_), .Y(_455_) );
NAND2X1 NAND2X1_65 ( .gnd(gnd), .vdd(vdd), .A(H_2_), .B(_4420_), .Y(_456_) );
AOI21X1 AOI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(_456_), .B(_455_), .C(_400__bF_buf10), .Y(_300__2_) );
AOI21X1 AOI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(H_2_), .B(micro_hash_ucr_a_2_), .C(_453_), .Y(_457_) );
NOR2X1 NOR2X1_65 ( .gnd(gnd), .vdd(vdd), .A(H_3_), .B(micro_hash_ucr_a_3_), .Y(_458_) );
INVX1 INVX1_73 ( .gnd(gnd), .vdd(vdd), .A(H_3_), .Y(_459_) );
INVX8 INVX8_12 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_3_), .Y(_460_) );
NOR2X1 NOR2X1_66 ( .gnd(gnd), .vdd(vdd), .A(_459_), .B(_460__bF_buf3), .Y(_461_) );
NOR2X1 NOR2X1_67 ( .gnd(gnd), .vdd(vdd), .A(_458_), .B(_461_), .Y(_462_) );
AND2X2 AND2X2_12 ( .gnd(gnd), .vdd(vdd), .A(_457_), .B(_462_), .Y(_463_) );
OAI21X1 OAI21X1_74 ( .gnd(gnd), .vdd(vdd), .A(_457_), .B(_462_), .C(micro_hash_ucr_pipe70_bF_buf1), .Y(_464_) );
OAI21X1 OAI21X1_75 ( .gnd(gnd), .vdd(vdd), .A(_459_), .B(micro_hash_ucr_pipe5), .C(_4479__bF_buf3), .Y(_465_) );
OAI21X1 OAI21X1_76 ( .gnd(gnd), .vdd(vdd), .A(_463_), .B(_464_), .C(_465_), .Y(_466_) );
NOR2X1 NOR2X1_68 ( .gnd(gnd), .vdd(vdd), .A(_400__bF_buf9), .B(_466_), .Y(_300__3_) );
XOR2X1 XOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(H_4_), .B(micro_hash_ucr_a_4_), .Y(_467_) );
INVX1 INVX1_74 ( .gnd(gnd), .vdd(vdd), .A(_461_), .Y(_468_) );
OAI21X1 OAI21X1_77 ( .gnd(gnd), .vdd(vdd), .A(_457_), .B(_458_), .C(_468_), .Y(_469_) );
XNOR2X1 XNOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_469_), .B(_467_), .Y(_470_) );
INVX2 INVX2_21 ( .gnd(gnd), .vdd(vdd), .A(H_4_), .Y(_471_) );
OAI21X1 OAI21X1_78 ( .gnd(gnd), .vdd(vdd), .A(_471_), .B(micro_hash_ucr_pipe5), .C(_4479__bF_buf2), .Y(_472_) );
NAND2X1 NAND2X1_66 ( .gnd(gnd), .vdd(vdd), .A(_472_), .B(_302__bF_buf10), .Y(_473_) );
AOI21X1 AOI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe70_bF_buf0), .B(_470_), .C(_473_), .Y(_300__4_) );
INVX8 INVX8_13 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_4_), .Y(_474_) );
NAND2X1 NAND2X1_67 ( .gnd(gnd), .vdd(vdd), .A(_467_), .B(_469_), .Y(_475_) );
OAI21X1 OAI21X1_79 ( .gnd(gnd), .vdd(vdd), .A(_471_), .B(_474__bF_buf3), .C(_475_), .Y(_476_) );
INVX2 INVX2_22 ( .gnd(gnd), .vdd(vdd), .A(_476_), .Y(_477_) );
NOR2X1 NOR2X1_69 ( .gnd(gnd), .vdd(vdd), .A(H_5_), .B(micro_hash_ucr_a_5_bF_buf3_), .Y(_478_) );
INVX2 INVX2_23 ( .gnd(gnd), .vdd(vdd), .A(H_5_), .Y(_479_) );
INVX8 INVX8_14 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_5_bF_buf2_), .Y(_480_) );
NOR2X1 NOR2X1_70 ( .gnd(gnd), .vdd(vdd), .A(_479_), .B(_480_), .Y(_481_) );
NOR2X1 NOR2X1_71 ( .gnd(gnd), .vdd(vdd), .A(_478_), .B(_481_), .Y(_482_) );
AND2X2 AND2X2_13 ( .gnd(gnd), .vdd(vdd), .A(_477_), .B(_482_), .Y(_483_) );
OAI21X1 OAI21X1_80 ( .gnd(gnd), .vdd(vdd), .A(_477_), .B(_482_), .C(micro_hash_ucr_pipe70_bF_buf3), .Y(_484_) );
OAI21X1 OAI21X1_81 ( .gnd(gnd), .vdd(vdd), .A(_479_), .B(micro_hash_ucr_pipe5), .C(_4479__bF_buf1), .Y(_485_) );
OAI21X1 OAI21X1_82 ( .gnd(gnd), .vdd(vdd), .A(_483_), .B(_484_), .C(_485_), .Y(_486_) );
NOR2X1 NOR2X1_72 ( .gnd(gnd), .vdd(vdd), .A(_400__bF_buf8), .B(_486_), .Y(_300__5_) );
XOR2X1 XOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(H_6_), .B(micro_hash_ucr_a_6_bF_buf3_), .Y(_487_) );
INVX1 INVX1_75 ( .gnd(gnd), .vdd(vdd), .A(_481_), .Y(_488_) );
OAI21X1 OAI21X1_83 ( .gnd(gnd), .vdd(vdd), .A(_477_), .B(_478_), .C(_488_), .Y(_489_) );
XOR2X1 XOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_489_), .B(_487_), .Y(_490_) );
INVX1 INVX1_76 ( .gnd(gnd), .vdd(vdd), .A(H_6_), .Y(_491_) );
OAI21X1 OAI21X1_84 ( .gnd(gnd), .vdd(vdd), .A(_491_), .B(micro_hash_ucr_pipe5), .C(_4479__bF_buf0), .Y(_492_) );
OAI21X1 OAI21X1_85 ( .gnd(gnd), .vdd(vdd), .A(_490_), .B(_4479__bF_buf3), .C(_492_), .Y(_493_) );
NOR2X1 NOR2X1_73 ( .gnd(gnd), .vdd(vdd), .A(_400__bF_buf7), .B(_493_), .Y(_300__6_) );
INVX8 INVX8_15 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_6_bF_buf2_), .Y(_494_) );
NAND2X1 NAND2X1_68 ( .gnd(gnd), .vdd(vdd), .A(_487_), .B(_489_), .Y(_495_) );
OAI21X1 OAI21X1_86 ( .gnd(gnd), .vdd(vdd), .A(_491_), .B(_494_), .C(_495_), .Y(_496_) );
XNOR2X1 XNOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(H_7_), .B(micro_hash_ucr_a_7_), .Y(_497_) );
AND2X2 AND2X2_14 ( .gnd(gnd), .vdd(vdd), .A(_496_), .B(_497_), .Y(_498_) );
OAI21X1 OAI21X1_87 ( .gnd(gnd), .vdd(vdd), .A(_496_), .B(_497_), .C(micro_hash_ucr_pipe70_bF_buf2), .Y(_499_) );
INVX1 INVX1_77 ( .gnd(gnd), .vdd(vdd), .A(H_7_), .Y(_500_) );
OAI21X1 OAI21X1_88 ( .gnd(gnd), .vdd(vdd), .A(_500_), .B(micro_hash_ucr_pipe5), .C(_4479__bF_buf2), .Y(_501_) );
OAI21X1 OAI21X1_89 ( .gnd(gnd), .vdd(vdd), .A(_498_), .B(_499_), .C(_501_), .Y(_502_) );
NOR2X1 NOR2X1_74 ( .gnd(gnd), .vdd(vdd), .A(_400__bF_buf6), .B(_502_), .Y(_300__7_) );
INVX4 INVX4_3 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_112_), .Y(_503_) );
AOI21X1 AOI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_152_), .B(_503_), .C(micro_hash_ucr_Wx_200_), .Y(_504_) );
OAI21X1 OAI21X1_90 ( .gnd(gnd), .vdd(vdd), .A(_503_), .B(micro_hash_ucr_Wx_152_), .C(_504_), .Y(_505_) );
AND2X2 AND2X2_15 ( .gnd(gnd), .vdd(vdd), .A(_505_), .B(_302__bF_buf9), .Y(_296__224_) );
INVX4 INVX4_4 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_113_), .Y(_506_) );
INVX2 INVX2_24 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_201_), .Y(_507_) );
OAI21X1 OAI21X1_91 ( .gnd(gnd), .vdd(vdd), .A(_506_), .B(micro_hash_ucr_Wx_153_), .C(_507_), .Y(_508_) );
AOI21X1 AOI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(_506_), .B(micro_hash_ucr_Wx_153_), .C(_508_), .Y(_509_) );
NOR2X1 NOR2X1_75 ( .gnd(gnd), .vdd(vdd), .A(_509_), .B(_400__bF_buf5), .Y(_296__225_) );
INVX4 INVX4_5 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_114_), .Y(_510_) );
INVX2 INVX2_25 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_202_), .Y(_511_) );
OAI21X1 OAI21X1_92 ( .gnd(gnd), .vdd(vdd), .A(_510_), .B(micro_hash_ucr_Wx_154_), .C(_511_), .Y(_512_) );
AOI21X1 AOI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(_510_), .B(micro_hash_ucr_Wx_154_), .C(_512_), .Y(_513_) );
NOR2X1 NOR2X1_76 ( .gnd(gnd), .vdd(vdd), .A(_513_), .B(_400__bF_buf4), .Y(_296__226_) );
INVX4 INVX4_6 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_115_), .Y(_514_) );
INVX1 INVX1_78 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_203_), .Y(_515_) );
OAI21X1 OAI21X1_93 ( .gnd(gnd), .vdd(vdd), .A(_514_), .B(micro_hash_ucr_Wx_155_), .C(_515_), .Y(_516_) );
AOI21X1 AOI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(_514_), .B(micro_hash_ucr_Wx_155_), .C(_516_), .Y(_517_) );
NOR2X1 NOR2X1_77 ( .gnd(gnd), .vdd(vdd), .A(_517_), .B(_400__bF_buf3), .Y(_296__227_) );
INVX4 INVX4_7 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_116_), .Y(_518_) );
AOI21X1 AOI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_156_), .B(_518_), .C(micro_hash_ucr_Wx_204_), .Y(_519_) );
OAI21X1 OAI21X1_94 ( .gnd(gnd), .vdd(vdd), .A(_518_), .B(micro_hash_ucr_Wx_156_), .C(_519_), .Y(_520_) );
AND2X2 AND2X2_16 ( .gnd(gnd), .vdd(vdd), .A(_520_), .B(_302__bF_buf8), .Y(_296__228_) );
INVX4 INVX4_8 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_117_), .Y(_521_) );
AOI21X1 AOI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_157_), .B(_521_), .C(micro_hash_ucr_Wx_205_), .Y(_522_) );
OAI21X1 OAI21X1_95 ( .gnd(gnd), .vdd(vdd), .A(_521_), .B(micro_hash_ucr_Wx_157_), .C(_522_), .Y(_523_) );
AND2X2 AND2X2_17 ( .gnd(gnd), .vdd(vdd), .A(_523_), .B(_302__bF_buf7), .Y(_296__229_) );
INVX4 INVX4_9 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_118_), .Y(_524_) );
INVX2 INVX2_26 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_206_), .Y(_525_) );
OAI21X1 OAI21X1_96 ( .gnd(gnd), .vdd(vdd), .A(_524_), .B(micro_hash_ucr_Wx_158_), .C(_525_), .Y(_526_) );
AOI21X1 AOI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(_524_), .B(micro_hash_ucr_Wx_158_), .C(_526_), .Y(_527_) );
NOR2X1 NOR2X1_78 ( .gnd(gnd), .vdd(vdd), .A(_527_), .B(_400__bF_buf2), .Y(_296__230_) );
INVX4 INVX4_10 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_119_), .Y(_528_) );
AOI21X1 AOI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_159_), .B(_528_), .C(micro_hash_ucr_Wx_207_), .Y(_529_) );
OAI21X1 OAI21X1_97 ( .gnd(gnd), .vdd(vdd), .A(_528_), .B(micro_hash_ucr_Wx_159_), .C(_529_), .Y(_530_) );
AND2X2 AND2X2_18 ( .gnd(gnd), .vdd(vdd), .A(_530_), .B(_302__bF_buf6), .Y(_296__231_) );
INVX4 INVX4_11 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_128_), .Y(_531_) );
AOI21X1 AOI21X1_66 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_168_), .B(_531_), .C(micro_hash_ucr_Wx_216_), .Y(_532_) );
OAI21X1 OAI21X1_98 ( .gnd(gnd), .vdd(vdd), .A(_531_), .B(micro_hash_ucr_Wx_168_), .C(_532_), .Y(_533_) );
AND2X2 AND2X2_19 ( .gnd(gnd), .vdd(vdd), .A(_533_), .B(_302__bF_buf5), .Y(_296__240_) );
INVX4 INVX4_12 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_129_), .Y(_534_) );
INVX2 INVX2_27 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_217_), .Y(_535_) );
OAI21X1 OAI21X1_99 ( .gnd(gnd), .vdd(vdd), .A(_534_), .B(micro_hash_ucr_Wx_169_), .C(_535_), .Y(_536_) );
AOI21X1 AOI21X1_67 ( .gnd(gnd), .vdd(vdd), .A(_534_), .B(micro_hash_ucr_Wx_169_), .C(_536_), .Y(_537_) );
NOR2X1 NOR2X1_79 ( .gnd(gnd), .vdd(vdd), .A(_537_), .B(_400__bF_buf1), .Y(_296__241_) );
INVX4 INVX4_13 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_130_), .Y(_538_) );
INVX2 INVX2_28 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_218_), .Y(_539_) );
OAI21X1 OAI21X1_100 ( .gnd(gnd), .vdd(vdd), .A(_538_), .B(micro_hash_ucr_Wx_170_), .C(_539_), .Y(_540_) );
AOI21X1 AOI21X1_68 ( .gnd(gnd), .vdd(vdd), .A(_538_), .B(micro_hash_ucr_Wx_170_), .C(_540_), .Y(_541_) );
NOR2X1 NOR2X1_80 ( .gnd(gnd), .vdd(vdd), .A(_541_), .B(_400__bF_buf0), .Y(_296__242_) );
INVX4 INVX4_14 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_131_), .Y(_542_) );
INVX1 INVX1_79 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_219_), .Y(_543_) );
OAI21X1 OAI21X1_101 ( .gnd(gnd), .vdd(vdd), .A(_542_), .B(micro_hash_ucr_Wx_171_), .C(_543_), .Y(_544_) );
AOI21X1 AOI21X1_69 ( .gnd(gnd), .vdd(vdd), .A(_542_), .B(micro_hash_ucr_Wx_171_), .C(_544_), .Y(_545_) );
NOR2X1 NOR2X1_81 ( .gnd(gnd), .vdd(vdd), .A(_545_), .B(_400__bF_buf12), .Y(_296__243_) );
INVX4 INVX4_15 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_132_), .Y(_546_) );
AOI21X1 AOI21X1_70 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_172_), .B(_546_), .C(micro_hash_ucr_Wx_220_), .Y(_547_) );
OAI21X1 OAI21X1_102 ( .gnd(gnd), .vdd(vdd), .A(_546_), .B(micro_hash_ucr_Wx_172_), .C(_547_), .Y(_548_) );
AND2X2 AND2X2_20 ( .gnd(gnd), .vdd(vdd), .A(_548_), .B(_302__bF_buf4), .Y(_296__244_) );
INVX4 INVX4_16 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_133_), .Y(_549_) );
INVX1 INVX1_80 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_221_), .Y(_550_) );
OAI21X1 OAI21X1_103 ( .gnd(gnd), .vdd(vdd), .A(_549_), .B(micro_hash_ucr_Wx_173_), .C(_550_), .Y(_551_) );
AOI21X1 AOI21X1_71 ( .gnd(gnd), .vdd(vdd), .A(_549_), .B(micro_hash_ucr_Wx_173_), .C(_551_), .Y(_552_) );
NOR2X1 NOR2X1_82 ( .gnd(gnd), .vdd(vdd), .A(_552_), .B(_400__bF_buf11), .Y(_296__245_) );
INVX4 INVX4_17 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_134_), .Y(_553_) );
INVX2 INVX2_29 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_222_), .Y(_554_) );
OAI21X1 OAI21X1_104 ( .gnd(gnd), .vdd(vdd), .A(_553_), .B(micro_hash_ucr_Wx_174_), .C(_554_), .Y(_555_) );
AOI21X1 AOI21X1_72 ( .gnd(gnd), .vdd(vdd), .A(_553_), .B(micro_hash_ucr_Wx_174_), .C(_555_), .Y(_556_) );
NOR2X1 NOR2X1_83 ( .gnd(gnd), .vdd(vdd), .A(_556_), .B(_400__bF_buf10), .Y(_296__246_) );
INVX4 INVX4_18 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_135_), .Y(_557_) );
AOI21X1 AOI21X1_73 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_175_), .B(_557_), .C(micro_hash_ucr_Wx_223_), .Y(_558_) );
OAI21X1 OAI21X1_105 ( .gnd(gnd), .vdd(vdd), .A(_557_), .B(micro_hash_ucr_Wx_175_), .C(_558_), .Y(_559_) );
AND2X2 AND2X2_21 ( .gnd(gnd), .vdd(vdd), .A(_559_), .B(_302__bF_buf3), .Y(_296__247_) );
INVX4 INVX4_19 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_120_), .Y(_560_) );
AOI21X1 AOI21X1_74 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_160_), .B(_560_), .C(micro_hash_ucr_Wx_208_), .Y(_561_) );
OAI21X1 OAI21X1_106 ( .gnd(gnd), .vdd(vdd), .A(_560_), .B(micro_hash_ucr_Wx_160_), .C(_561_), .Y(_562_) );
AND2X2 AND2X2_22 ( .gnd(gnd), .vdd(vdd), .A(_562_), .B(_302__bF_buf2), .Y(_296__232_) );
INVX4 INVX4_20 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_121_), .Y(_563_) );
AOI21X1 AOI21X1_75 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_161_), .B(_563_), .C(micro_hash_ucr_Wx_209_), .Y(_564_) );
OAI21X1 OAI21X1_107 ( .gnd(gnd), .vdd(vdd), .A(_563_), .B(micro_hash_ucr_Wx_161_), .C(_564_), .Y(_565_) );
AND2X2 AND2X2_23 ( .gnd(gnd), .vdd(vdd), .A(_565_), .B(_302__bF_buf1), .Y(_296__233_) );
INVX4 INVX4_21 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_122_), .Y(_566_) );
INVX2 INVX2_30 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_210_), .Y(_567_) );
OAI21X1 OAI21X1_108 ( .gnd(gnd), .vdd(vdd), .A(_566_), .B(micro_hash_ucr_Wx_162_), .C(_567_), .Y(_568_) );
AOI21X1 AOI21X1_76 ( .gnd(gnd), .vdd(vdd), .A(_566_), .B(micro_hash_ucr_Wx_162_), .C(_568_), .Y(_569_) );
NOR2X1 NOR2X1_84 ( .gnd(gnd), .vdd(vdd), .A(_569_), .B(_400__bF_buf9), .Y(_296__234_) );
INVX4 INVX4_22 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_123_), .Y(_570_) );
INVX1 INVX1_81 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_211_), .Y(_571_) );
OAI21X1 OAI21X1_109 ( .gnd(gnd), .vdd(vdd), .A(_570_), .B(micro_hash_ucr_Wx_163_), .C(_571_), .Y(_572_) );
AOI21X1 AOI21X1_77 ( .gnd(gnd), .vdd(vdd), .A(_570_), .B(micro_hash_ucr_Wx_163_), .C(_572_), .Y(_573_) );
NOR2X1 NOR2X1_85 ( .gnd(gnd), .vdd(vdd), .A(_573_), .B(_400__bF_buf8), .Y(_296__235_) );
INVX4 INVX4_23 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_124_), .Y(_574_) );
AOI21X1 AOI21X1_78 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_164_), .B(_574_), .C(micro_hash_ucr_Wx_212_), .Y(_575_) );
OAI21X1 OAI21X1_110 ( .gnd(gnd), .vdd(vdd), .A(_574_), .B(micro_hash_ucr_Wx_164_), .C(_575_), .Y(_576_) );
AND2X2 AND2X2_24 ( .gnd(gnd), .vdd(vdd), .A(_576_), .B(_302__bF_buf0), .Y(_296__236_) );
INVX4 INVX4_24 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_125_), .Y(_577_) );
AOI21X1 AOI21X1_79 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_165_), .B(_577_), .C(micro_hash_ucr_Wx_213_), .Y(_578_) );
OAI21X1 OAI21X1_111 ( .gnd(gnd), .vdd(vdd), .A(_577_), .B(micro_hash_ucr_Wx_165_), .C(_578_), .Y(_579_) );
AND2X2 AND2X2_25 ( .gnd(gnd), .vdd(vdd), .A(_579_), .B(_302__bF_buf13), .Y(_296__237_) );
INVX4 INVX4_25 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_126_), .Y(_580_) );
INVX2 INVX2_31 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_214_), .Y(_581_) );
OAI21X1 OAI21X1_112 ( .gnd(gnd), .vdd(vdd), .A(_580_), .B(micro_hash_ucr_Wx_166_), .C(_581_), .Y(_582_) );
AOI21X1 AOI21X1_80 ( .gnd(gnd), .vdd(vdd), .A(_580_), .B(micro_hash_ucr_Wx_166_), .C(_582_), .Y(_583_) );
NOR2X1 NOR2X1_86 ( .gnd(gnd), .vdd(vdd), .A(_583_), .B(_400__bF_buf7), .Y(_296__238_) );
INVX4 INVX4_26 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_127_), .Y(_584_) );
AOI21X1 AOI21X1_81 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_167_), .B(_584_), .C(micro_hash_ucr_Wx_215_), .Y(_585_) );
OAI21X1 OAI21X1_113 ( .gnd(gnd), .vdd(vdd), .A(_584_), .B(micro_hash_ucr_Wx_167_), .C(_585_), .Y(_586_) );
AND2X2 AND2X2_26 ( .gnd(gnd), .vdd(vdd), .A(_586_), .B(_302__bF_buf12), .Y(_296__239_) );
INVX2 INVX2_32 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_176_), .Y(_587_) );
OAI21X1 OAI21X1_114 ( .gnd(gnd), .vdd(vdd), .A(_531_), .B(micro_hash_ucr_Wx_88_), .C(_587_), .Y(_588_) );
AOI21X1 AOI21X1_82 ( .gnd(gnd), .vdd(vdd), .A(_531_), .B(micro_hash_ucr_Wx_88_), .C(_588_), .Y(_589_) );
NOR2X1 NOR2X1_87 ( .gnd(gnd), .vdd(vdd), .A(_589_), .B(_400__bF_buf6), .Y(_296__200_) );
INVX2 INVX2_33 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_177_), .Y(_590_) );
OAI21X1 OAI21X1_115 ( .gnd(gnd), .vdd(vdd), .A(_534_), .B(micro_hash_ucr_Wx_89_), .C(_590_), .Y(_591_) );
AOI21X1 AOI21X1_83 ( .gnd(gnd), .vdd(vdd), .A(_534_), .B(micro_hash_ucr_Wx_89_), .C(_591_), .Y(_592_) );
NOR2X1 NOR2X1_88 ( .gnd(gnd), .vdd(vdd), .A(_592_), .B(_400__bF_buf5), .Y(_296__201_) );
INVX4 INVX4_27 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_178_), .Y(_593_) );
OAI21X1 OAI21X1_116 ( .gnd(gnd), .vdd(vdd), .A(_538_), .B(micro_hash_ucr_Wx_90_), .C(_593_), .Y(_594_) );
AOI21X1 AOI21X1_84 ( .gnd(gnd), .vdd(vdd), .A(_538_), .B(micro_hash_ucr_Wx_90_), .C(_594_), .Y(_595_) );
NOR2X1 NOR2X1_89 ( .gnd(gnd), .vdd(vdd), .A(_595_), .B(_400__bF_buf4), .Y(_296__202_) );
INVX2 INVX2_34 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_179_), .Y(_596_) );
OAI21X1 OAI21X1_117 ( .gnd(gnd), .vdd(vdd), .A(_542_), .B(micro_hash_ucr_Wx_91_), .C(_596_), .Y(_597_) );
AOI21X1 AOI21X1_85 ( .gnd(gnd), .vdd(vdd), .A(_542_), .B(micro_hash_ucr_Wx_91_), .C(_597_), .Y(_598_) );
NOR2X1 NOR2X1_90 ( .gnd(gnd), .vdd(vdd), .A(_598_), .B(_400__bF_buf3), .Y(_296__203_) );
INVX4 INVX4_28 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_180_), .Y(_599_) );
OAI21X1 OAI21X1_118 ( .gnd(gnd), .vdd(vdd), .A(_546_), .B(micro_hash_ucr_Wx_92_), .C(_599_), .Y(_600_) );
AOI21X1 AOI21X1_86 ( .gnd(gnd), .vdd(vdd), .A(_546_), .B(micro_hash_ucr_Wx_92_), .C(_600_), .Y(_601_) );
NOR2X1 NOR2X1_91 ( .gnd(gnd), .vdd(vdd), .A(_601_), .B(_400__bF_buf2), .Y(_296__204_) );
INVX2 INVX2_35 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_181_), .Y(_602_) );
OAI21X1 OAI21X1_119 ( .gnd(gnd), .vdd(vdd), .A(_549_), .B(micro_hash_ucr_Wx_93_), .C(_602_), .Y(_603_) );
AOI21X1 AOI21X1_87 ( .gnd(gnd), .vdd(vdd), .A(_549_), .B(micro_hash_ucr_Wx_93_), .C(_603_), .Y(_604_) );
NOR2X1 NOR2X1_92 ( .gnd(gnd), .vdd(vdd), .A(_604_), .B(_400__bF_buf1), .Y(_296__205_) );
INVX2 INVX2_36 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_182_), .Y(_605_) );
OAI21X1 OAI21X1_120 ( .gnd(gnd), .vdd(vdd), .A(_553_), .B(micro_hash_ucr_Wx_94_), .C(_605_), .Y(_606_) );
AOI21X1 AOI21X1_88 ( .gnd(gnd), .vdd(vdd), .A(_553_), .B(micro_hash_ucr_Wx_94_), .C(_606_), .Y(_607_) );
NOR2X1 NOR2X1_93 ( .gnd(gnd), .vdd(vdd), .A(_607_), .B(_400__bF_buf0), .Y(_296__206_) );
INVX4 INVX4_29 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_183_), .Y(_608_) );
OAI21X1 OAI21X1_121 ( .gnd(gnd), .vdd(vdd), .A(_557_), .B(micro_hash_ucr_Wx_95_), .C(_608_), .Y(_609_) );
AOI21X1 AOI21X1_89 ( .gnd(gnd), .vdd(vdd), .A(_557_), .B(micro_hash_ucr_Wx_95_), .C(_609_), .Y(_610_) );
NOR2X1 NOR2X1_94 ( .gnd(gnd), .vdd(vdd), .A(_610_), .B(_400__bF_buf12), .Y(_296__207_) );
INVX2 INVX2_37 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_144_), .Y(_611_) );
INVX1 INVX1_82 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_192_), .Y(_612_) );
OAI21X1 OAI21X1_122 ( .gnd(gnd), .vdd(vdd), .A(_611_), .B(micro_hash_ucr_Wx_104_), .C(_612_), .Y(_613_) );
AOI21X1 AOI21X1_90 ( .gnd(gnd), .vdd(vdd), .A(_611_), .B(micro_hash_ucr_Wx_104_), .C(_613_), .Y(_614_) );
NOR2X1 NOR2X1_95 ( .gnd(gnd), .vdd(vdd), .A(_614_), .B(_400__bF_buf11), .Y(_296__216_) );
INVX2 INVX2_38 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_145_), .Y(_615_) );
INVX2 INVX2_39 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_193_), .Y(_616_) );
OAI21X1 OAI21X1_123 ( .gnd(gnd), .vdd(vdd), .A(_615_), .B(micro_hash_ucr_Wx_105_), .C(_616_), .Y(_617_) );
AOI21X1 AOI21X1_91 ( .gnd(gnd), .vdd(vdd), .A(_615_), .B(micro_hash_ucr_Wx_105_), .C(_617_), .Y(_618_) );
NOR2X1 NOR2X1_96 ( .gnd(gnd), .vdd(vdd), .A(_618_), .B(_400__bF_buf10), .Y(_296__217_) );
INVX4 INVX4_30 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_146_), .Y(_619_) );
INVX2 INVX2_40 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_194_), .Y(_620_) );
OAI21X1 OAI21X1_124 ( .gnd(gnd), .vdd(vdd), .A(_619_), .B(micro_hash_ucr_Wx_106_), .C(_620_), .Y(_621_) );
AOI21X1 AOI21X1_92 ( .gnd(gnd), .vdd(vdd), .A(_619_), .B(micro_hash_ucr_Wx_106_), .C(_621_), .Y(_622_) );
NOR2X1 NOR2X1_97 ( .gnd(gnd), .vdd(vdd), .A(_622_), .B(_400__bF_buf9), .Y(_296__218_) );
INVX2 INVX2_41 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_147_), .Y(_623_) );
INVX1 INVX1_83 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_195_), .Y(_624_) );
OAI21X1 OAI21X1_125 ( .gnd(gnd), .vdd(vdd), .A(_623_), .B(micro_hash_ucr_Wx_107_), .C(_624_), .Y(_625_) );
AOI21X1 AOI21X1_93 ( .gnd(gnd), .vdd(vdd), .A(_623_), .B(micro_hash_ucr_Wx_107_), .C(_625_), .Y(_626_) );
NOR2X1 NOR2X1_98 ( .gnd(gnd), .vdd(vdd), .A(_626_), .B(_400__bF_buf8), .Y(_296__219_) );
INVX2 INVX2_42 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_148_), .Y(_627_) );
AOI21X1 AOI21X1_94 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_108_), .B(_627_), .C(micro_hash_ucr_Wx_196_), .Y(_628_) );
OAI21X1 OAI21X1_126 ( .gnd(gnd), .vdd(vdd), .A(_627_), .B(micro_hash_ucr_Wx_108_), .C(_628_), .Y(_629_) );
AND2X2 AND2X2_27 ( .gnd(gnd), .vdd(vdd), .A(_629_), .B(_302__bF_buf11), .Y(_296__220_) );
INVX2 INVX2_43 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_149_), .Y(_630_) );
AOI21X1 AOI21X1_95 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_109_), .B(_630_), .C(micro_hash_ucr_Wx_197_), .Y(_631_) );
OAI21X1 OAI21X1_127 ( .gnd(gnd), .vdd(vdd), .A(_630_), .B(micro_hash_ucr_Wx_109_), .C(_631_), .Y(_632_) );
AND2X2 AND2X2_28 ( .gnd(gnd), .vdd(vdd), .A(_632_), .B(_302__bF_buf10), .Y(_296__221_) );
INVX4 INVX4_31 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_150_), .Y(_633_) );
INVX1 INVX1_84 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_198_), .Y(_634_) );
OAI21X1 OAI21X1_128 ( .gnd(gnd), .vdd(vdd), .A(_633_), .B(micro_hash_ucr_Wx_110_), .C(_634_), .Y(_635_) );
AOI21X1 AOI21X1_96 ( .gnd(gnd), .vdd(vdd), .A(_633_), .B(micro_hash_ucr_Wx_110_), .C(_635_), .Y(_636_) );
NOR2X1 NOR2X1_99 ( .gnd(gnd), .vdd(vdd), .A(_636_), .B(_400__bF_buf7), .Y(_296__222_) );
INVX4 INVX4_32 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_151_), .Y(_637_) );
AOI21X1 AOI21X1_97 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_111_), .B(_637_), .C(micro_hash_ucr_Wx_199_), .Y(_638_) );
OAI21X1 OAI21X1_129 ( .gnd(gnd), .vdd(vdd), .A(_637_), .B(micro_hash_ucr_Wx_111_), .C(_638_), .Y(_639_) );
AND2X2 AND2X2_29 ( .gnd(gnd), .vdd(vdd), .A(_639_), .B(_302__bF_buf9), .Y(_296__223_) );
INVX4 INVX4_33 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_96_), .Y(_640_) );
INVX1 INVX1_85 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_184_), .Y(_641_) );
OAI21X1 OAI21X1_130 ( .gnd(gnd), .vdd(vdd), .A(_640_), .B(micro_hash_ucr_Wx_136_), .C(_641_), .Y(_642_) );
AOI21X1 AOI21X1_98 ( .gnd(gnd), .vdd(vdd), .A(_640_), .B(micro_hash_ucr_Wx_136_), .C(_642_), .Y(_643_) );
NOR2X1 NOR2X1_100 ( .gnd(gnd), .vdd(vdd), .A(_643_), .B(_400__bF_buf6), .Y(_296__208_) );
INVX4 INVX4_34 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_97_), .Y(_644_) );
INVX1 INVX1_86 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_185_), .Y(_645_) );
OAI21X1 OAI21X1_131 ( .gnd(gnd), .vdd(vdd), .A(_644_), .B(micro_hash_ucr_Wx_137_), .C(_645_), .Y(_646_) );
AOI21X1 AOI21X1_99 ( .gnd(gnd), .vdd(vdd), .A(_644_), .B(micro_hash_ucr_Wx_137_), .C(_646_), .Y(_647_) );
NOR2X1 NOR2X1_101 ( .gnd(gnd), .vdd(vdd), .A(_647_), .B(_400__bF_buf5), .Y(_296__209_) );
INVX4 INVX4_35 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_98_), .Y(_648_) );
INVX2 INVX2_44 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_186_), .Y(_649_) );
OAI21X1 OAI21X1_132 ( .gnd(gnd), .vdd(vdd), .A(_648_), .B(micro_hash_ucr_Wx_138_), .C(_649_), .Y(_650_) );
AOI21X1 AOI21X1_100 ( .gnd(gnd), .vdd(vdd), .A(_648_), .B(micro_hash_ucr_Wx_138_), .C(_650_), .Y(_651_) );
NOR2X1 NOR2X1_102 ( .gnd(gnd), .vdd(vdd), .A(_651_), .B(_400__bF_buf4), .Y(_296__210_) );
INVX4 INVX4_36 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_99_), .Y(_652_) );
INVX1 INVX1_87 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_187_), .Y(_653_) );
OAI21X1 OAI21X1_133 ( .gnd(gnd), .vdd(vdd), .A(_652_), .B(micro_hash_ucr_Wx_139_), .C(_653_), .Y(_654_) );
AOI21X1 AOI21X1_101 ( .gnd(gnd), .vdd(vdd), .A(_652_), .B(micro_hash_ucr_Wx_139_), .C(_654_), .Y(_655_) );
NOR2X1 NOR2X1_103 ( .gnd(gnd), .vdd(vdd), .A(_655_), .B(_400__bF_buf3), .Y(_296__211_) );
INVX2 INVX2_45 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_100_), .Y(_656_) );
AOI21X1 AOI21X1_102 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_140_), .B(_656_), .C(micro_hash_ucr_Wx_188_), .Y(_657_) );
OAI21X1 OAI21X1_134 ( .gnd(gnd), .vdd(vdd), .A(_656_), .B(micro_hash_ucr_Wx_140_), .C(_657_), .Y(_658_) );
AND2X2 AND2X2_30 ( .gnd(gnd), .vdd(vdd), .A(_658_), .B(_302__bF_buf8), .Y(_296__212_) );
INVX4 INVX4_37 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_101_), .Y(_659_) );
INVX1 INVX1_88 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_189_), .Y(_660_) );
OAI21X1 OAI21X1_135 ( .gnd(gnd), .vdd(vdd), .A(_659_), .B(micro_hash_ucr_Wx_141_), .C(_660_), .Y(_661_) );
AOI21X1 AOI21X1_103 ( .gnd(gnd), .vdd(vdd), .A(_659_), .B(micro_hash_ucr_Wx_141_), .C(_661_), .Y(_662_) );
NOR2X1 NOR2X1_104 ( .gnd(gnd), .vdd(vdd), .A(_662_), .B(_400__bF_buf2), .Y(_296__213_) );
INVX4 INVX4_38 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_102_), .Y(_663_) );
INVX2 INVX2_46 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_190_), .Y(_664_) );
OAI21X1 OAI21X1_136 ( .gnd(gnd), .vdd(vdd), .A(_663_), .B(micro_hash_ucr_Wx_142_), .C(_664_), .Y(_665_) );
AOI21X1 AOI21X1_104 ( .gnd(gnd), .vdd(vdd), .A(_663_), .B(micro_hash_ucr_Wx_142_), .C(_665_), .Y(_666_) );
NOR2X1 NOR2X1_105 ( .gnd(gnd), .vdd(vdd), .A(_666_), .B(_400__bF_buf1), .Y(_296__214_) );
INVX4 INVX4_39 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_103_), .Y(_667_) );
AOI21X1 AOI21X1_105 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_143_), .B(_667_), .C(micro_hash_ucr_Wx_191_), .Y(_668_) );
OAI21X1 OAI21X1_137 ( .gnd(gnd), .vdd(vdd), .A(_667_), .B(micro_hash_ucr_Wx_143_), .C(_668_), .Y(_669_) );
AND2X2 AND2X2_31 ( .gnd(gnd), .vdd(vdd), .A(_669_), .B(_302__bF_buf7), .Y(_296__215_) );
INVX2 INVX2_47 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_104_), .Y(_670_) );
AOI21X1 AOI21X1_106 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_64_), .B(_670_), .C(micro_hash_ucr_Wx_152_), .Y(_671_) );
OAI21X1 OAI21X1_138 ( .gnd(gnd), .vdd(vdd), .A(_670_), .B(micro_hash_ucr_Wx_64_), .C(_671_), .Y(_672_) );
AND2X2 AND2X2_32 ( .gnd(gnd), .vdd(vdd), .A(_672_), .B(_302__bF_buf6), .Y(_296__176_) );
INVX2 INVX2_48 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_105_), .Y(_673_) );
AOI21X1 AOI21X1_107 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_65_), .B(_673_), .C(micro_hash_ucr_Wx_153_), .Y(_674_) );
OAI21X1 OAI21X1_139 ( .gnd(gnd), .vdd(vdd), .A(_673_), .B(micro_hash_ucr_Wx_65_), .C(_674_), .Y(_675_) );
AND2X2 AND2X2_33 ( .gnd(gnd), .vdd(vdd), .A(_675_), .B(_302__bF_buf5), .Y(_296__177_) );
INVX4 INVX4_40 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_106_), .Y(_676_) );
INVX2 INVX2_49 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_154_), .Y(_677_) );
OAI21X1 OAI21X1_140 ( .gnd(gnd), .vdd(vdd), .A(_676_), .B(micro_hash_ucr_Wx_66_), .C(_677_), .Y(_678_) );
AOI21X1 AOI21X1_108 ( .gnd(gnd), .vdd(vdd), .A(_676_), .B(micro_hash_ucr_Wx_66_), .C(_678_), .Y(_679_) );
NOR2X1 NOR2X1_106 ( .gnd(gnd), .vdd(vdd), .A(_679_), .B(_400__bF_buf0), .Y(_296__178_) );
INVX2 INVX2_50 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_107_), .Y(_680_) );
INVX1 INVX1_89 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_155_), .Y(_681_) );
OAI21X1 OAI21X1_141 ( .gnd(gnd), .vdd(vdd), .A(_680_), .B(micro_hash_ucr_Wx_67_), .C(_681_), .Y(_682_) );
AOI21X1 AOI21X1_109 ( .gnd(gnd), .vdd(vdd), .A(_680_), .B(micro_hash_ucr_Wx_67_), .C(_682_), .Y(_683_) );
NOR2X1 NOR2X1_107 ( .gnd(gnd), .vdd(vdd), .A(_683_), .B(_400__bF_buf12), .Y(_296__179_) );
INVX2 INVX2_51 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_108_), .Y(_684_) );
AOI21X1 AOI21X1_110 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_68_), .B(_684_), .C(micro_hash_ucr_Wx_156_), .Y(_685_) );
OAI21X1 OAI21X1_142 ( .gnd(gnd), .vdd(vdd), .A(_684_), .B(micro_hash_ucr_Wx_68_), .C(_685_), .Y(_686_) );
AND2X2 AND2X2_34 ( .gnd(gnd), .vdd(vdd), .A(_686_), .B(_302__bF_buf4), .Y(_296__180_) );
INVX2 INVX2_52 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_109_), .Y(_687_) );
AOI21X1 AOI21X1_111 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_69_), .B(_687_), .C(micro_hash_ucr_Wx_157_), .Y(_688_) );
OAI21X1 OAI21X1_143 ( .gnd(gnd), .vdd(vdd), .A(_687_), .B(micro_hash_ucr_Wx_69_), .C(_688_), .Y(_689_) );
AND2X2 AND2X2_35 ( .gnd(gnd), .vdd(vdd), .A(_689_), .B(_302__bF_buf3), .Y(_296__181_) );
INVX4 INVX4_41 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_70_), .Y(_690_) );
INVX2 INVX2_53 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_158_), .Y(_691_) );
OAI21X1 OAI21X1_144 ( .gnd(gnd), .vdd(vdd), .A(_690_), .B(micro_hash_ucr_Wx_110_), .C(_691_), .Y(_692_) );
AOI21X1 AOI21X1_112 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_110_), .B(_690_), .C(_692_), .Y(_693_) );
NOR2X1 NOR2X1_108 ( .gnd(gnd), .vdd(vdd), .A(_693_), .B(_400__bF_buf11), .Y(_296__182_) );
INVX4 INVX4_42 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_111_), .Y(_694_) );
AOI21X1 AOI21X1_113 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_71_), .B(_694_), .C(micro_hash_ucr_Wx_159_), .Y(_695_) );
OAI21X1 OAI21X1_145 ( .gnd(gnd), .vdd(vdd), .A(_694_), .B(micro_hash_ucr_Wx_71_), .C(_695_), .Y(_696_) );
AND2X2 AND2X2_36 ( .gnd(gnd), .vdd(vdd), .A(_696_), .B(_302__bF_buf2), .Y(_296__183_) );
AOI21X1 AOI21X1_114 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_80_), .B(_560_), .C(micro_hash_ucr_Wx_168_), .Y(_697_) );
OAI21X1 OAI21X1_146 ( .gnd(gnd), .vdd(vdd), .A(_560_), .B(micro_hash_ucr_Wx_80_), .C(_697_), .Y(_698_) );
AND2X2 AND2X2_37 ( .gnd(gnd), .vdd(vdd), .A(_698_), .B(_302__bF_buf1), .Y(_296__192_) );
INVX2 INVX2_54 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_169_), .Y(_699_) );
OAI21X1 OAI21X1_147 ( .gnd(gnd), .vdd(vdd), .A(_563_), .B(micro_hash_ucr_Wx_81_), .C(_699_), .Y(_700_) );
AOI21X1 AOI21X1_115 ( .gnd(gnd), .vdd(vdd), .A(_563_), .B(micro_hash_ucr_Wx_81_), .C(_700_), .Y(_701_) );
NOR2X1 NOR2X1_109 ( .gnd(gnd), .vdd(vdd), .A(_701_), .B(_400__bF_buf10), .Y(_296__193_) );
INVX2 INVX2_55 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_170_), .Y(_702_) );
OAI21X1 OAI21X1_148 ( .gnd(gnd), .vdd(vdd), .A(_566_), .B(micro_hash_ucr_Wx_82_), .C(_702_), .Y(_703_) );
AOI21X1 AOI21X1_116 ( .gnd(gnd), .vdd(vdd), .A(_566_), .B(micro_hash_ucr_Wx_82_), .C(_703_), .Y(_704_) );
NOR2X1 NOR2X1_110 ( .gnd(gnd), .vdd(vdd), .A(_704_), .B(_400__bF_buf9), .Y(_296__194_) );
INVX1 INVX1_90 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_171_), .Y(_705_) );
OAI21X1 OAI21X1_149 ( .gnd(gnd), .vdd(vdd), .A(_570_), .B(micro_hash_ucr_Wx_83_), .C(_705_), .Y(_706_) );
AOI21X1 AOI21X1_117 ( .gnd(gnd), .vdd(vdd), .A(_570_), .B(micro_hash_ucr_Wx_83_), .C(_706_), .Y(_707_) );
NOR2X1 NOR2X1_111 ( .gnd(gnd), .vdd(vdd), .A(_707_), .B(_400__bF_buf8), .Y(_296__195_) );
INVX1 INVX1_91 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_172_), .Y(_708_) );
OAI21X1 OAI21X1_150 ( .gnd(gnd), .vdd(vdd), .A(_574_), .B(micro_hash_ucr_Wx_84_), .C(_708_), .Y(_709_) );
AOI21X1 AOI21X1_118 ( .gnd(gnd), .vdd(vdd), .A(_574_), .B(micro_hash_ucr_Wx_84_), .C(_709_), .Y(_710_) );
NOR2X1 NOR2X1_112 ( .gnd(gnd), .vdd(vdd), .A(_710_), .B(_400__bF_buf7), .Y(_296__196_) );
INVX1 INVX1_92 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_173_), .Y(_711_) );
OAI21X1 OAI21X1_151 ( .gnd(gnd), .vdd(vdd), .A(_577_), .B(micro_hash_ucr_Wx_85_), .C(_711_), .Y(_712_) );
AOI21X1 AOI21X1_119 ( .gnd(gnd), .vdd(vdd), .A(_577_), .B(micro_hash_ucr_Wx_85_), .C(_712_), .Y(_713_) );
NOR2X1 NOR2X1_113 ( .gnd(gnd), .vdd(vdd), .A(_713_), .B(_400__bF_buf6), .Y(_296__197_) );
INVX1 INVX1_93 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_174_), .Y(_714_) );
OAI21X1 OAI21X1_152 ( .gnd(gnd), .vdd(vdd), .A(_580_), .B(micro_hash_ucr_Wx_86_), .C(_714_), .Y(_715_) );
AOI21X1 AOI21X1_120 ( .gnd(gnd), .vdd(vdd), .A(_580_), .B(micro_hash_ucr_Wx_86_), .C(_715_), .Y(_716_) );
NOR2X1 NOR2X1_114 ( .gnd(gnd), .vdd(vdd), .A(_716_), .B(_400__bF_buf5), .Y(_296__198_) );
AOI21X1 AOI21X1_121 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_87_), .B(_584_), .C(micro_hash_ucr_Wx_175_), .Y(_717_) );
OAI21X1 OAI21X1_153 ( .gnd(gnd), .vdd(vdd), .A(_584_), .B(micro_hash_ucr_Wx_87_), .C(_717_), .Y(_718_) );
AND2X2 AND2X2_38 ( .gnd(gnd), .vdd(vdd), .A(_718_), .B(_302__bF_buf0), .Y(_296__199_) );
INVX1 INVX1_94 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_160_), .Y(_719_) );
OAI21X1 OAI21X1_154 ( .gnd(gnd), .vdd(vdd), .A(_503_), .B(micro_hash_ucr_Wx_72_), .C(_719_), .Y(_720_) );
AOI21X1 AOI21X1_122 ( .gnd(gnd), .vdd(vdd), .A(_503_), .B(micro_hash_ucr_Wx_72_), .C(_720_), .Y(_721_) );
NOR2X1 NOR2X1_115 ( .gnd(gnd), .vdd(vdd), .A(_721_), .B(_400__bF_buf4), .Y(_296__184_) );
INVX2 INVX2_56 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_161_), .Y(_722_) );
OAI21X1 OAI21X1_155 ( .gnd(gnd), .vdd(vdd), .A(_506_), .B(micro_hash_ucr_Wx_73_), .C(_722_), .Y(_723_) );
AOI21X1 AOI21X1_123 ( .gnd(gnd), .vdd(vdd), .A(_506_), .B(micro_hash_ucr_Wx_73_), .C(_723_), .Y(_724_) );
NOR2X1 NOR2X1_116 ( .gnd(gnd), .vdd(vdd), .A(_724_), .B(_400__bF_buf3), .Y(_296__185_) );
INVX2 INVX2_57 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_162_), .Y(_725_) );
OAI21X1 OAI21X1_156 ( .gnd(gnd), .vdd(vdd), .A(_510_), .B(micro_hash_ucr_Wx_74_), .C(_725_), .Y(_726_) );
AOI21X1 AOI21X1_124 ( .gnd(gnd), .vdd(vdd), .A(_510_), .B(micro_hash_ucr_Wx_74_), .C(_726_), .Y(_727_) );
NOR2X1 NOR2X1_117 ( .gnd(gnd), .vdd(vdd), .A(_727_), .B(_400__bF_buf2), .Y(_296__186_) );
INVX1 INVX1_95 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_163_), .Y(_728_) );
OAI21X1 OAI21X1_157 ( .gnd(gnd), .vdd(vdd), .A(_514_), .B(micro_hash_ucr_Wx_75_), .C(_728_), .Y(_729_) );
AOI21X1 AOI21X1_125 ( .gnd(gnd), .vdd(vdd), .A(_514_), .B(micro_hash_ucr_Wx_75_), .C(_729_), .Y(_730_) );
NOR2X1 NOR2X1_118 ( .gnd(gnd), .vdd(vdd), .A(_730_), .B(_400__bF_buf1), .Y(_296__187_) );
AOI21X1 AOI21X1_126 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_76_), .B(_518_), .C(micro_hash_ucr_Wx_164_), .Y(_731_) );
OAI21X1 OAI21X1_158 ( .gnd(gnd), .vdd(vdd), .A(_518_), .B(micro_hash_ucr_Wx_76_), .C(_731_), .Y(_732_) );
AND2X2 AND2X2_39 ( .gnd(gnd), .vdd(vdd), .A(_732_), .B(_302__bF_buf13), .Y(_296__188_) );
AOI21X1 AOI21X1_127 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_77_), .B(_521_), .C(micro_hash_ucr_Wx_165_), .Y(_733_) );
OAI21X1 OAI21X1_159 ( .gnd(gnd), .vdd(vdd), .A(_521_), .B(micro_hash_ucr_Wx_77_), .C(_733_), .Y(_734_) );
AND2X2 AND2X2_40 ( .gnd(gnd), .vdd(vdd), .A(_734_), .B(_302__bF_buf12), .Y(_296__189_) );
INVX2 INVX2_58 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_166_), .Y(_735_) );
OAI21X1 OAI21X1_160 ( .gnd(gnd), .vdd(vdd), .A(_524_), .B(micro_hash_ucr_Wx_78_), .C(_735_), .Y(_736_) );
AOI21X1 AOI21X1_128 ( .gnd(gnd), .vdd(vdd), .A(_524_), .B(micro_hash_ucr_Wx_78_), .C(_736_), .Y(_737_) );
NOR2X1 NOR2X1_119 ( .gnd(gnd), .vdd(vdd), .A(_737_), .B(_400__bF_buf0), .Y(_296__190_) );
AOI21X1 AOI21X1_129 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_79_), .B(_528_), .C(micro_hash_ucr_Wx_167_), .Y(_738_) );
OAI21X1 OAI21X1_161 ( .gnd(gnd), .vdd(vdd), .A(_528_), .B(micro_hash_ucr_Wx_79_), .C(_738_), .Y(_739_) );
AND2X2 AND2X2_41 ( .gnd(gnd), .vdd(vdd), .A(_739_), .B(_302__bF_buf11), .Y(_296__191_) );
INVX2 INVX2_59 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_80_), .Y(_740_) );
OAI21X1 OAI21X1_162 ( .gnd(gnd), .vdd(vdd), .A(_740_), .B(micro_hash_ucr_Wx_40_), .C(_531_), .Y(_741_) );
AOI21X1 AOI21X1_130 ( .gnd(gnd), .vdd(vdd), .A(_740_), .B(micro_hash_ucr_Wx_40_), .C(_741_), .Y(_742_) );
NOR2X1 NOR2X1_120 ( .gnd(gnd), .vdd(vdd), .A(_742_), .B(_400__bF_buf12), .Y(_296__152_) );
INVX2 INVX2_60 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_81_), .Y(_743_) );
OAI21X1 OAI21X1_163 ( .gnd(gnd), .vdd(vdd), .A(_743_), .B(micro_hash_ucr_Wx_41_), .C(_534_), .Y(_744_) );
AOI21X1 AOI21X1_131 ( .gnd(gnd), .vdd(vdd), .A(_743_), .B(micro_hash_ucr_Wx_41_), .C(_744_), .Y(_745_) );
NOR2X1 NOR2X1_121 ( .gnd(gnd), .vdd(vdd), .A(_745_), .B(_400__bF_buf11), .Y(_296__153_) );
INVX2 INVX2_61 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_82_), .Y(_746_) );
OAI21X1 OAI21X1_164 ( .gnd(gnd), .vdd(vdd), .A(_746_), .B(micro_hash_ucr_Wx_42_), .C(_538_), .Y(_747_) );
AOI21X1 AOI21X1_132 ( .gnd(gnd), .vdd(vdd), .A(_746_), .B(micro_hash_ucr_Wx_42_), .C(_747_), .Y(_748_) );
NOR2X1 NOR2X1_122 ( .gnd(gnd), .vdd(vdd), .A(_748_), .B(_400__bF_buf10), .Y(_296__154_) );
INVX2 INVX2_62 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_83_), .Y(_749_) );
OAI21X1 OAI21X1_165 ( .gnd(gnd), .vdd(vdd), .A(_749_), .B(micro_hash_ucr_Wx_43_), .C(_542_), .Y(_750_) );
AOI21X1 AOI21X1_133 ( .gnd(gnd), .vdd(vdd), .A(_749_), .B(micro_hash_ucr_Wx_43_), .C(_750_), .Y(_751_) );
NOR2X1 NOR2X1_123 ( .gnd(gnd), .vdd(vdd), .A(_751_), .B(_400__bF_buf9), .Y(_296__155_) );
INVX2 INVX2_63 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_84_), .Y(_752_) );
OAI21X1 OAI21X1_166 ( .gnd(gnd), .vdd(vdd), .A(_752_), .B(micro_hash_ucr_Wx_44_), .C(_546_), .Y(_753_) );
AOI21X1 AOI21X1_134 ( .gnd(gnd), .vdd(vdd), .A(_752_), .B(micro_hash_ucr_Wx_44_), .C(_753_), .Y(_754_) );
NOR2X1 NOR2X1_124 ( .gnd(gnd), .vdd(vdd), .A(_754_), .B(_400__bF_buf8), .Y(_296__156_) );
INVX2 INVX2_64 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_85_), .Y(_755_) );
OAI21X1 OAI21X1_167 ( .gnd(gnd), .vdd(vdd), .A(_755_), .B(micro_hash_ucr_Wx_45_), .C(_549_), .Y(_756_) );
AOI21X1 AOI21X1_135 ( .gnd(gnd), .vdd(vdd), .A(_755_), .B(micro_hash_ucr_Wx_45_), .C(_756_), .Y(_757_) );
NOR2X1 NOR2X1_125 ( .gnd(gnd), .vdd(vdd), .A(_757_), .B(_400__bF_buf7), .Y(_296__157_) );
INVX4 INVX4_43 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_86_), .Y(_758_) );
OAI21X1 OAI21X1_168 ( .gnd(gnd), .vdd(vdd), .A(_758_), .B(micro_hash_ucr_Wx_46_), .C(_553_), .Y(_759_) );
AOI21X1 AOI21X1_136 ( .gnd(gnd), .vdd(vdd), .A(_758_), .B(micro_hash_ucr_Wx_46_), .C(_759_), .Y(_760_) );
NOR2X1 NOR2X1_126 ( .gnd(gnd), .vdd(vdd), .A(_760_), .B(_400__bF_buf6), .Y(_296__158_) );
XNOR2X1 XNOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_87_), .B(micro_hash_ucr_Wx_47_), .Y(_761_) );
AOI21X1 AOI21X1_137 ( .gnd(gnd), .vdd(vdd), .A(_557_), .B(_761_), .C(_400__bF_buf5), .Y(_296__159_) );
OAI21X1 OAI21X1_169 ( .gnd(gnd), .vdd(vdd), .A(_640_), .B(micro_hash_ucr_Wx_56_), .C(_611_), .Y(_762_) );
AOI21X1 AOI21X1_138 ( .gnd(gnd), .vdd(vdd), .A(_640_), .B(micro_hash_ucr_Wx_56_), .C(_762_), .Y(_763_) );
NOR2X1 NOR2X1_127 ( .gnd(gnd), .vdd(vdd), .A(_763_), .B(_400__bF_buf4), .Y(_296__168_) );
OAI21X1 OAI21X1_170 ( .gnd(gnd), .vdd(vdd), .A(_644_), .B(micro_hash_ucr_Wx_57_), .C(_615_), .Y(_764_) );
AOI21X1 AOI21X1_139 ( .gnd(gnd), .vdd(vdd), .A(_644_), .B(micro_hash_ucr_Wx_57_), .C(_764_), .Y(_765_) );
NOR2X1 NOR2X1_128 ( .gnd(gnd), .vdd(vdd), .A(_765_), .B(_400__bF_buf3), .Y(_296__169_) );
OAI21X1 OAI21X1_171 ( .gnd(gnd), .vdd(vdd), .A(_648_), .B(micro_hash_ucr_Wx_58_), .C(_619_), .Y(_766_) );
AOI21X1 AOI21X1_140 ( .gnd(gnd), .vdd(vdd), .A(_648_), .B(micro_hash_ucr_Wx_58_), .C(_766_), .Y(_767_) );
NOR2X1 NOR2X1_129 ( .gnd(gnd), .vdd(vdd), .A(_767_), .B(_400__bF_buf2), .Y(_296__170_) );
OAI21X1 OAI21X1_172 ( .gnd(gnd), .vdd(vdd), .A(_652_), .B(micro_hash_ucr_Wx_59_), .C(_623_), .Y(_768_) );
AOI21X1 AOI21X1_141 ( .gnd(gnd), .vdd(vdd), .A(_652_), .B(micro_hash_ucr_Wx_59_), .C(_768_), .Y(_769_) );
NOR2X1 NOR2X1_130 ( .gnd(gnd), .vdd(vdd), .A(_769_), .B(_400__bF_buf1), .Y(_296__171_) );
OAI21X1 OAI21X1_173 ( .gnd(gnd), .vdd(vdd), .A(_656_), .B(micro_hash_ucr_Wx_60_), .C(_627_), .Y(_770_) );
AOI21X1 AOI21X1_142 ( .gnd(gnd), .vdd(vdd), .A(_656_), .B(micro_hash_ucr_Wx_60_), .C(_770_), .Y(_771_) );
NOR2X1 NOR2X1_131 ( .gnd(gnd), .vdd(vdd), .A(_771_), .B(_400__bF_buf0), .Y(_296__172_) );
OAI21X1 OAI21X1_174 ( .gnd(gnd), .vdd(vdd), .A(_659_), .B(micro_hash_ucr_Wx_61_), .C(_630_), .Y(_772_) );
AOI21X1 AOI21X1_143 ( .gnd(gnd), .vdd(vdd), .A(_659_), .B(micro_hash_ucr_Wx_61_), .C(_772_), .Y(_773_) );
NOR2X1 NOR2X1_132 ( .gnd(gnd), .vdd(vdd), .A(_773_), .B(_400__bF_buf12), .Y(_296__173_) );
OAI21X1 OAI21X1_175 ( .gnd(gnd), .vdd(vdd), .A(_663_), .B(micro_hash_ucr_Wx_62_), .C(_633_), .Y(_774_) );
AOI21X1 AOI21X1_144 ( .gnd(gnd), .vdd(vdd), .A(_663_), .B(micro_hash_ucr_Wx_62_), .C(_774_), .Y(_775_) );
NOR2X1 NOR2X1_133 ( .gnd(gnd), .vdd(vdd), .A(_775_), .B(_400__bF_buf11), .Y(_296__174_) );
OAI21X1 OAI21X1_176 ( .gnd(gnd), .vdd(vdd), .A(_667_), .B(micro_hash_ucr_Wx_63_), .C(_637_), .Y(_776_) );
AOI21X1 AOI21X1_145 ( .gnd(gnd), .vdd(vdd), .A(_667_), .B(micro_hash_ucr_Wx_63_), .C(_776_), .Y(_777_) );
NOR2X1 NOR2X1_134 ( .gnd(gnd), .vdd(vdd), .A(_777_), .B(_400__bF_buf10), .Y(_296__175_) );
INVX2 INVX2_65 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_88_), .Y(_778_) );
INVX1 INVX1_96 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_136_), .Y(_779_) );
OAI21X1 OAI21X1_177 ( .gnd(gnd), .vdd(vdd), .A(_778_), .B(micro_hash_ucr_Wx_48_), .C(_779_), .Y(_780_) );
AOI21X1 AOI21X1_146 ( .gnd(gnd), .vdd(vdd), .A(_778_), .B(micro_hash_ucr_Wx_48_), .C(_780_), .Y(_781_) );
NOR2X1 NOR2X1_135 ( .gnd(gnd), .vdd(vdd), .A(_781_), .B(_400__bF_buf9), .Y(_296__160_) );
INVX2 INVX2_66 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_89_), .Y(_782_) );
INVX1 INVX1_97 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_137_), .Y(_783_) );
OAI21X1 OAI21X1_178 ( .gnd(gnd), .vdd(vdd), .A(_782_), .B(micro_hash_ucr_Wx_49_), .C(_783_), .Y(_784_) );
AOI21X1 AOI21X1_147 ( .gnd(gnd), .vdd(vdd), .A(_782_), .B(micro_hash_ucr_Wx_49_), .C(_784_), .Y(_785_) );
NOR2X1 NOR2X1_136 ( .gnd(gnd), .vdd(vdd), .A(_785_), .B(_400__bF_buf8), .Y(_296__161_) );
INVX2 INVX2_67 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_90_), .Y(_786_) );
INVX2 INVX2_68 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_138_), .Y(_787_) );
OAI21X1 OAI21X1_179 ( .gnd(gnd), .vdd(vdd), .A(_786_), .B(micro_hash_ucr_Wx_50_), .C(_787_), .Y(_788_) );
AOI21X1 AOI21X1_148 ( .gnd(gnd), .vdd(vdd), .A(_786_), .B(micro_hash_ucr_Wx_50_), .C(_788_), .Y(_789_) );
NOR2X1 NOR2X1_137 ( .gnd(gnd), .vdd(vdd), .A(_789_), .B(_400__bF_buf7), .Y(_296__162_) );
INVX2 INVX2_69 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_91_), .Y(_790_) );
INVX1 INVX1_98 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_139_), .Y(_791_) );
OAI21X1 OAI21X1_180 ( .gnd(gnd), .vdd(vdd), .A(_790_), .B(micro_hash_ucr_Wx_51_), .C(_791_), .Y(_792_) );
AOI21X1 AOI21X1_149 ( .gnd(gnd), .vdd(vdd), .A(_790_), .B(micro_hash_ucr_Wx_51_), .C(_792_), .Y(_793_) );
NOR2X1 NOR2X1_138 ( .gnd(gnd), .vdd(vdd), .A(_793_), .B(_400__bF_buf6), .Y(_296__163_) );
INVX2 INVX2_70 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_92_), .Y(_794_) );
AOI21X1 AOI21X1_150 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_52_), .B(_794_), .C(micro_hash_ucr_Wx_140_), .Y(_795_) );
OAI21X1 OAI21X1_181 ( .gnd(gnd), .vdd(vdd), .A(_794_), .B(micro_hash_ucr_Wx_52_), .C(_795_), .Y(_796_) );
AND2X2 AND2X2_42 ( .gnd(gnd), .vdd(vdd), .A(_796_), .B(_302__bF_buf10), .Y(_296__164_) );
INVX2 INVX2_71 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_93_), .Y(_797_) );
INVX1 INVX1_99 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_141_), .Y(_798_) );
OAI21X1 OAI21X1_182 ( .gnd(gnd), .vdd(vdd), .A(_797_), .B(micro_hash_ucr_Wx_53_), .C(_798_), .Y(_799_) );
AOI21X1 AOI21X1_151 ( .gnd(gnd), .vdd(vdd), .A(_797_), .B(micro_hash_ucr_Wx_53_), .C(_799_), .Y(_800_) );
NOR2X1 NOR2X1_139 ( .gnd(gnd), .vdd(vdd), .A(_800_), .B(_400__bF_buf5), .Y(_296__165_) );
INVX4 INVX4_44 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_94_), .Y(_801_) );
INVX2 INVX2_72 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_142_), .Y(_802_) );
OAI21X1 OAI21X1_183 ( .gnd(gnd), .vdd(vdd), .A(_801_), .B(micro_hash_ucr_Wx_54_), .C(_802_), .Y(_803_) );
AOI21X1 AOI21X1_152 ( .gnd(gnd), .vdd(vdd), .A(_801_), .B(micro_hash_ucr_Wx_54_), .C(_803_), .Y(_804_) );
NOR2X1 NOR2X1_140 ( .gnd(gnd), .vdd(vdd), .A(_804_), .B(_400__bF_buf4), .Y(_296__166_) );
INVX1 INVX1_100 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_143_), .Y(_805_) );
XNOR2X1 XNOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_95_), .B(micro_hash_ucr_Wx_55_), .Y(_806_) );
AOI21X1 AOI21X1_153 ( .gnd(gnd), .vdd(vdd), .A(_805_), .B(_806_), .C(_400__bF_buf3), .Y(_296__167_) );
INVX2 INVX2_73 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_56_), .Y(_807_) );
OAI21X1 OAI21X1_184 ( .gnd(gnd), .vdd(vdd), .A(_807_), .B(micro_hash_ucr_Wx_16_), .C(_670_), .Y(_808_) );
AOI21X1 AOI21X1_154 ( .gnd(gnd), .vdd(vdd), .A(_807_), .B(micro_hash_ucr_Wx_16_), .C(_808_), .Y(_809_) );
NOR2X1 NOR2X1_141 ( .gnd(gnd), .vdd(vdd), .A(_809_), .B(_400__bF_buf2), .Y(_296__128_) );
INVX2 INVX2_74 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_57_), .Y(_810_) );
OAI21X1 OAI21X1_185 ( .gnd(gnd), .vdd(vdd), .A(_810_), .B(micro_hash_ucr_Wx_17_), .C(_673_), .Y(_811_) );
AOI21X1 AOI21X1_155 ( .gnd(gnd), .vdd(vdd), .A(_810_), .B(micro_hash_ucr_Wx_17_), .C(_811_), .Y(_812_) );
NOR2X1 NOR2X1_142 ( .gnd(gnd), .vdd(vdd), .A(_812_), .B(_400__bF_buf1), .Y(_296__129_) );
INVX2 INVX2_75 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_58_), .Y(_813_) );
OAI21X1 OAI21X1_186 ( .gnd(gnd), .vdd(vdd), .A(_813_), .B(micro_hash_ucr_Wx_18_), .C(_676_), .Y(_814_) );
AOI21X1 AOI21X1_156 ( .gnd(gnd), .vdd(vdd), .A(_813_), .B(micro_hash_ucr_Wx_18_), .C(_814_), .Y(_815_) );
NOR2X1 NOR2X1_143 ( .gnd(gnd), .vdd(vdd), .A(_815_), .B(_400__bF_buf0), .Y(_296__130_) );
INVX2 INVX2_76 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_59_), .Y(_816_) );
OAI21X1 OAI21X1_187 ( .gnd(gnd), .vdd(vdd), .A(_816_), .B(micro_hash_ucr_Wx_19_), .C(_680_), .Y(_817_) );
AOI21X1 AOI21X1_157 ( .gnd(gnd), .vdd(vdd), .A(_816_), .B(micro_hash_ucr_Wx_19_), .C(_817_), .Y(_818_) );
NOR2X1 NOR2X1_144 ( .gnd(gnd), .vdd(vdd), .A(_818_), .B(_400__bF_buf12), .Y(_296__131_) );
INVX2 INVX2_77 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_60_), .Y(_819_) );
OAI21X1 OAI21X1_188 ( .gnd(gnd), .vdd(vdd), .A(_819_), .B(micro_hash_ucr_Wx_20_), .C(_684_), .Y(_820_) );
AOI21X1 AOI21X1_158 ( .gnd(gnd), .vdd(vdd), .A(_819_), .B(micro_hash_ucr_Wx_20_), .C(_820_), .Y(_821_) );
NOR2X1 NOR2X1_145 ( .gnd(gnd), .vdd(vdd), .A(_821_), .B(_400__bF_buf11), .Y(_296__132_) );
INVX2 INVX2_78 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_61_), .Y(_822_) );
OAI21X1 OAI21X1_189 ( .gnd(gnd), .vdd(vdd), .A(_822_), .B(micro_hash_ucr_Wx_21_), .C(_687_), .Y(_823_) );
AOI21X1 AOI21X1_159 ( .gnd(gnd), .vdd(vdd), .A(_822_), .B(micro_hash_ucr_Wx_21_), .C(_823_), .Y(_824_) );
NOR2X1 NOR2X1_146 ( .gnd(gnd), .vdd(vdd), .A(_824_), .B(_400__bF_buf10), .Y(_296__133_) );
INVX2 INVX2_79 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_62_), .Y(_825_) );
AOI21X1 AOI21X1_160 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_22_), .B(_825_), .C(micro_hash_ucr_Wx_110_), .Y(_826_) );
OAI21X1 OAI21X1_190 ( .gnd(gnd), .vdd(vdd), .A(_825_), .B(micro_hash_ucr_Wx_22_), .C(_826_), .Y(_827_) );
AND2X2 AND2X2_43 ( .gnd(gnd), .vdd(vdd), .A(_827_), .B(_302__bF_buf9), .Y(_296__134_) );
XNOR2X1 XNOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_63_), .B(micro_hash_ucr_Wx_23_), .Y(_828_) );
AOI21X1 AOI21X1_161 ( .gnd(gnd), .vdd(vdd), .A(_694_), .B(_828_), .C(_400__bF_buf9), .Y(_296__135_) );
INVX2 INVX2_80 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_72_), .Y(_829_) );
OAI21X1 OAI21X1_191 ( .gnd(gnd), .vdd(vdd), .A(_829_), .B(micro_hash_ucr_Wx_32_), .C(_560_), .Y(_830_) );
AOI21X1 AOI21X1_162 ( .gnd(gnd), .vdd(vdd), .A(_829_), .B(micro_hash_ucr_Wx_32_), .C(_830_), .Y(_831_) );
NOR2X1 NOR2X1_147 ( .gnd(gnd), .vdd(vdd), .A(_831_), .B(_400__bF_buf8), .Y(_296__144_) );
INVX2 INVX2_81 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_73_), .Y(_832_) );
OAI21X1 OAI21X1_192 ( .gnd(gnd), .vdd(vdd), .A(_832_), .B(micro_hash_ucr_Wx_33_), .C(_563_), .Y(_833_) );
AOI21X1 AOI21X1_163 ( .gnd(gnd), .vdd(vdd), .A(_832_), .B(micro_hash_ucr_Wx_33_), .C(_833_), .Y(_834_) );
NOR2X1 NOR2X1_148 ( .gnd(gnd), .vdd(vdd), .A(_834_), .B(_400__bF_buf7), .Y(_296__145_) );
INVX4 INVX4_45 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_74_), .Y(_835_) );
OAI21X1 OAI21X1_193 ( .gnd(gnd), .vdd(vdd), .A(_835_), .B(micro_hash_ucr_Wx_34_), .C(_566_), .Y(_836_) );
AOI21X1 AOI21X1_164 ( .gnd(gnd), .vdd(vdd), .A(_835_), .B(micro_hash_ucr_Wx_34_), .C(_836_), .Y(_837_) );
NOR2X1 NOR2X1_149 ( .gnd(gnd), .vdd(vdd), .A(_837_), .B(_400__bF_buf6), .Y(_296__146_) );
INVX2 INVX2_82 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_75_), .Y(_838_) );
OAI21X1 OAI21X1_194 ( .gnd(gnd), .vdd(vdd), .A(_838_), .B(micro_hash_ucr_Wx_35_), .C(_570_), .Y(_839_) );
AOI21X1 AOI21X1_165 ( .gnd(gnd), .vdd(vdd), .A(_838_), .B(micro_hash_ucr_Wx_35_), .C(_839_), .Y(_840_) );
NOR2X1 NOR2X1_150 ( .gnd(gnd), .vdd(vdd), .A(_840_), .B(_400__bF_buf5), .Y(_296__147_) );
INVX2 INVX2_83 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_76_), .Y(_841_) );
OAI21X1 OAI21X1_195 ( .gnd(gnd), .vdd(vdd), .A(_841_), .B(micro_hash_ucr_Wx_36_), .C(_574_), .Y(_842_) );
AOI21X1 AOI21X1_166 ( .gnd(gnd), .vdd(vdd), .A(_841_), .B(micro_hash_ucr_Wx_36_), .C(_842_), .Y(_843_) );
NOR2X1 NOR2X1_151 ( .gnd(gnd), .vdd(vdd), .A(_843_), .B(_400__bF_buf4), .Y(_296__148_) );
INVX2 INVX2_84 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_77_), .Y(_844_) );
OAI21X1 OAI21X1_196 ( .gnd(gnd), .vdd(vdd), .A(_844_), .B(micro_hash_ucr_Wx_37_), .C(_577_), .Y(_845_) );
AOI21X1 AOI21X1_167 ( .gnd(gnd), .vdd(vdd), .A(_844_), .B(micro_hash_ucr_Wx_37_), .C(_845_), .Y(_846_) );
NOR2X1 NOR2X1_152 ( .gnd(gnd), .vdd(vdd), .A(_846_), .B(_400__bF_buf3), .Y(_296__149_) );
INVX2 INVX2_85 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_78_), .Y(_847_) );
OAI21X1 OAI21X1_197 ( .gnd(gnd), .vdd(vdd), .A(_847_), .B(micro_hash_ucr_Wx_38_), .C(_580_), .Y(_848_) );
AOI21X1 AOI21X1_168 ( .gnd(gnd), .vdd(vdd), .A(_847_), .B(micro_hash_ucr_Wx_38_), .C(_848_), .Y(_849_) );
NOR2X1 NOR2X1_153 ( .gnd(gnd), .vdd(vdd), .A(_849_), .B(_400__bF_buf2), .Y(_296__150_) );
INVX2 INVX2_86 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_79_), .Y(_850_) );
OAI21X1 OAI21X1_198 ( .gnd(gnd), .vdd(vdd), .A(_850_), .B(micro_hash_ucr_Wx_39_), .C(_584_), .Y(_851_) );
AOI21X1 AOI21X1_169 ( .gnd(gnd), .vdd(vdd), .A(_850_), .B(micro_hash_ucr_Wx_39_), .C(_851_), .Y(_852_) );
NOR2X1 NOR2X1_154 ( .gnd(gnd), .vdd(vdd), .A(_852_), .B(_400__bF_buf1), .Y(_296__151_) );
INVX2 INVX2_87 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_64_), .Y(_853_) );
OAI21X1 OAI21X1_199 ( .gnd(gnd), .vdd(vdd), .A(_853_), .B(micro_hash_ucr_Wx_24_), .C(_503_), .Y(_854_) );
AOI21X1 AOI21X1_170 ( .gnd(gnd), .vdd(vdd), .A(_853_), .B(micro_hash_ucr_Wx_24_), .C(_854_), .Y(_855_) );
NOR2X1 NOR2X1_155 ( .gnd(gnd), .vdd(vdd), .A(_855_), .B(_400__bF_buf0), .Y(_296__136_) );
INVX4 INVX4_46 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_65_), .Y(_856_) );
OAI21X1 OAI21X1_200 ( .gnd(gnd), .vdd(vdd), .A(_856_), .B(micro_hash_ucr_Wx_25_), .C(_506_), .Y(_857_) );
AOI21X1 AOI21X1_171 ( .gnd(gnd), .vdd(vdd), .A(_856_), .B(micro_hash_ucr_Wx_25_), .C(_857_), .Y(_858_) );
NOR2X1 NOR2X1_156 ( .gnd(gnd), .vdd(vdd), .A(_858_), .B(_400__bF_buf12), .Y(_296__137_) );
INVX4 INVX4_47 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_66_), .Y(_859_) );
OAI21X1 OAI21X1_201 ( .gnd(gnd), .vdd(vdd), .A(_859_), .B(micro_hash_ucr_Wx_26_), .C(_510_), .Y(_860_) );
AOI21X1 AOI21X1_172 ( .gnd(gnd), .vdd(vdd), .A(_859_), .B(micro_hash_ucr_Wx_26_), .C(_860_), .Y(_861_) );
NOR2X1 NOR2X1_157 ( .gnd(gnd), .vdd(vdd), .A(_861_), .B(_400__bF_buf11), .Y(_296__138_) );
INVX2 INVX2_88 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_67_), .Y(_862_) );
OAI21X1 OAI21X1_202 ( .gnd(gnd), .vdd(vdd), .A(_862_), .B(micro_hash_ucr_Wx_27_), .C(_514_), .Y(_863_) );
AOI21X1 AOI21X1_173 ( .gnd(gnd), .vdd(vdd), .A(_862_), .B(micro_hash_ucr_Wx_27_), .C(_863_), .Y(_864_) );
NOR2X1 NOR2X1_158 ( .gnd(gnd), .vdd(vdd), .A(_864_), .B(_400__bF_buf10), .Y(_296__139_) );
INVX2 INVX2_89 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_68_), .Y(_865_) );
OAI21X1 OAI21X1_203 ( .gnd(gnd), .vdd(vdd), .A(_865_), .B(micro_hash_ucr_Wx_28_), .C(_518_), .Y(_866_) );
AOI21X1 AOI21X1_174 ( .gnd(gnd), .vdd(vdd), .A(_865_), .B(micro_hash_ucr_Wx_28_), .C(_866_), .Y(_867_) );
NOR2X1 NOR2X1_159 ( .gnd(gnd), .vdd(vdd), .A(_867_), .B(_400__bF_buf9), .Y(_296__140_) );
INVX2 INVX2_90 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_69_), .Y(_868_) );
OAI21X1 OAI21X1_204 ( .gnd(gnd), .vdd(vdd), .A(_868_), .B(micro_hash_ucr_Wx_29_), .C(_521_), .Y(_869_) );
AOI21X1 AOI21X1_175 ( .gnd(gnd), .vdd(vdd), .A(_868_), .B(micro_hash_ucr_Wx_29_), .C(_869_), .Y(_870_) );
NOR2X1 NOR2X1_160 ( .gnd(gnd), .vdd(vdd), .A(_870_), .B(_400__bF_buf8), .Y(_296__141_) );
OAI21X1 OAI21X1_205 ( .gnd(gnd), .vdd(vdd), .A(_690_), .B(micro_hash_ucr_Wx_30_), .C(_524_), .Y(_871_) );
AOI21X1 AOI21X1_176 ( .gnd(gnd), .vdd(vdd), .A(_690_), .B(micro_hash_ucr_Wx_30_), .C(_871_), .Y(_872_) );
NOR2X1 NOR2X1_161 ( .gnd(gnd), .vdd(vdd), .A(_872_), .B(_400__bF_buf7), .Y(_296__142_) );
INVX2 INVX2_91 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_71_), .Y(_873_) );
OAI21X1 OAI21X1_206 ( .gnd(gnd), .vdd(vdd), .A(_873_), .B(micro_hash_ucr_Wx_31_), .C(_528_), .Y(_874_) );
AOI21X1 AOI21X1_177 ( .gnd(gnd), .vdd(vdd), .A(_873_), .B(micro_hash_ucr_Wx_31_), .C(_874_), .Y(_875_) );
NOR2X1 NOR2X1_162 ( .gnd(gnd), .vdd(vdd), .A(_875_), .B(_400__bF_buf6), .Y(_296__143_) );
AND2X2 AND2X2_44 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf8), .B(concatenador_data_out_104_), .Y(_296__104_) );
AND2X2 AND2X2_45 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf7), .B(concatenador_data_out_105_), .Y(_296__105_) );
AND2X2 AND2X2_46 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf6), .B(concatenador_data_out_106_), .Y(_296__106_) );
AND2X2 AND2X2_47 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf5), .B(concatenador_data_out_107_), .Y(_296__107_) );
AND2X2 AND2X2_48 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf4), .B(concatenador_data_out_108_), .Y(_296__108_) );
AND2X2 AND2X2_49 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf3), .B(concatenador_data_out_109_), .Y(_296__109_) );
AND2X2 AND2X2_50 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf2), .B(concatenador_data_out_110_), .Y(_296__110_) );
AND2X2 AND2X2_51 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf1), .B(concatenador_data_out_111_), .Y(_296__111_) );
AND2X2 AND2X2_52 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf0), .B(concatenador_data_out_120_), .Y(_296__120_) );
AND2X2 AND2X2_53 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf13), .B(concatenador_data_out_121_), .Y(_296__121_) );
AND2X2 AND2X2_54 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf12), .B(concatenador_data_out_122_), .Y(_296__122_) );
AND2X2 AND2X2_55 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf11), .B(concatenador_data_out_123_), .Y(_296__123_) );
AND2X2 AND2X2_56 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf10), .B(concatenador_data_out_124_), .Y(_296__124_) );
AND2X2 AND2X2_57 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf9), .B(concatenador_data_out_125_), .Y(_296__125_) );
AND2X2 AND2X2_58 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf8), .B(concatenador_data_out_126_), .Y(_296__126_) );
AND2X2 AND2X2_59 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf7), .B(concatenador_data_out_127_), .Y(_296__127_) );
AND2X2 AND2X2_60 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf6), .B(concatenador_data_out_112_), .Y(_296__112_) );
AND2X2 AND2X2_61 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf5), .B(concatenador_data_out_113_), .Y(_296__113_) );
AND2X2 AND2X2_62 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf4), .B(concatenador_data_out_114_), .Y(_296__114_) );
AND2X2 AND2X2_63 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf3), .B(concatenador_data_out_115_), .Y(_296__115_) );
AND2X2 AND2X2_64 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf2), .B(concatenador_data_out_116_), .Y(_296__116_) );
AND2X2 AND2X2_65 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf1), .B(concatenador_data_out_117_), .Y(_296__117_) );
AND2X2 AND2X2_66 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf0), .B(concatenador_data_out_118_), .Y(_296__118_) );
AND2X2 AND2X2_67 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf13), .B(concatenador_data_out_119_), .Y(_296__119_) );
AND2X2 AND2X2_68 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf12), .B(concatenador_data_out_80_), .Y(_296__80_) );
AND2X2 AND2X2_69 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf11), .B(concatenador_data_out_81_), .Y(_296__81_) );
AND2X2 AND2X2_70 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf10), .B(concatenador_data_out_82_), .Y(_296__82_) );
AND2X2 AND2X2_71 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf9), .B(concatenador_data_out_83_), .Y(_296__83_) );
AND2X2 AND2X2_72 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf8), .B(concatenador_data_out_84_), .Y(_296__84_) );
AND2X2 AND2X2_73 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf7), .B(concatenador_data_out_85_), .Y(_296__85_) );
AND2X2 AND2X2_74 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf6), .B(concatenador_data_out_86_), .Y(_296__86_) );
AND2X2 AND2X2_75 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf5), .B(concatenador_data_out_87_), .Y(_296__87_) );
AND2X2 AND2X2_76 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf4), .B(concatenador_data_out_96_), .Y(_296__96_) );
AND2X2 AND2X2_77 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf3), .B(concatenador_data_out_97_), .Y(_296__97_) );
AND2X2 AND2X2_78 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf2), .B(concatenador_data_out_98_), .Y(_296__98_) );
AND2X2 AND2X2_79 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf1), .B(concatenador_data_out_99_), .Y(_296__99_) );
AND2X2 AND2X2_80 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf0), .B(concatenador_data_out_100_), .Y(_296__100_) );
AND2X2 AND2X2_81 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf13), .B(concatenador_data_out_101_), .Y(_296__101_) );
AND2X2 AND2X2_82 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf12), .B(concatenador_data_out_102_), .Y(_296__102_) );
AND2X2 AND2X2_83 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf11), .B(concatenador_data_out_103_), .Y(_296__103_) );
AND2X2 AND2X2_84 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf10), .B(concatenador_data_out_88_), .Y(_296__88_) );
AND2X2 AND2X2_85 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf9), .B(concatenador_data_out_89_), .Y(_296__89_) );
AND2X2 AND2X2_86 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf8), .B(concatenador_data_out_90_), .Y(_296__90_) );
AND2X2 AND2X2_87 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf7), .B(concatenador_data_out_91_), .Y(_296__91_) );
AND2X2 AND2X2_88 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf6), .B(concatenador_data_out_92_), .Y(_296__92_) );
AND2X2 AND2X2_89 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf5), .B(concatenador_data_out_93_), .Y(_296__93_) );
AND2X2 AND2X2_90 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf4), .B(concatenador_data_out_94_), .Y(_296__94_) );
AND2X2 AND2X2_91 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf3), .B(concatenador_data_out_95_), .Y(_296__95_) );
AND2X2 AND2X2_92 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf2), .B(concatenador_data_out_56_), .Y(_296__56_) );
AND2X2 AND2X2_93 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf1), .B(concatenador_data_out_57_), .Y(_296__57_) );
AND2X2 AND2X2_94 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf0), .B(concatenador_data_out_58_), .Y(_296__58_) );
AND2X2 AND2X2_95 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf13), .B(concatenador_data_out_59_), .Y(_296__59_) );
AND2X2 AND2X2_96 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf12), .B(concatenador_data_out_60_), .Y(_296__60_) );
AND2X2 AND2X2_97 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf11), .B(concatenador_data_out_61_), .Y(_296__61_) );
AND2X2 AND2X2_98 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf10), .B(concatenador_data_out_62_), .Y(_296__62_) );
AND2X2 AND2X2_99 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf9), .B(concatenador_data_out_63_), .Y(_296__63_) );
AND2X2 AND2X2_100 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf8), .B(concatenador_data_out_72_), .Y(_296__72_) );
AND2X2 AND2X2_101 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf7), .B(concatenador_data_out_73_), .Y(_296__73_) );
AND2X2 AND2X2_102 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf6), .B(concatenador_data_out_74_), .Y(_296__74_) );
AND2X2 AND2X2_103 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf5), .B(concatenador_data_out_75_), .Y(_296__75_) );
AND2X2 AND2X2_104 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf4), .B(concatenador_data_out_76_), .Y(_296__76_) );
AND2X2 AND2X2_105 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf3), .B(concatenador_data_out_77_), .Y(_296__77_) );
AND2X2 AND2X2_106 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf2), .B(concatenador_data_out_78_), .Y(_296__78_) );
AND2X2 AND2X2_107 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf1), .B(concatenador_data_out_79_), .Y(_296__79_) );
AND2X2 AND2X2_108 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf0), .B(concatenador_data_out_64_), .Y(_296__64_) );
AND2X2 AND2X2_109 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf13), .B(concatenador_data_out_65_), .Y(_296__65_) );
AND2X2 AND2X2_110 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf12), .B(concatenador_data_out_66_), .Y(_296__66_) );
AND2X2 AND2X2_111 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf11), .B(concatenador_data_out_67_), .Y(_296__67_) );
AND2X2 AND2X2_112 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf10), .B(concatenador_data_out_68_), .Y(_296__68_) );
AND2X2 AND2X2_113 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf9), .B(concatenador_data_out_69_), .Y(_296__69_) );
AND2X2 AND2X2_114 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf8), .B(concatenador_data_out_70_), .Y(_296__70_) );
AND2X2 AND2X2_115 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf7), .B(concatenador_data_out_71_), .Y(_296__71_) );
AND2X2 AND2X2_116 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf6), .B(concatenador_data_out_32_), .Y(_296__32_) );
AND2X2 AND2X2_117 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf5), .B(concatenador_data_out_33_), .Y(_296__33_) );
AND2X2 AND2X2_118 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf4), .B(concatenador_data_out_34_), .Y(_296__34_) );
AND2X2 AND2X2_119 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf3), .B(concatenador_data_out_35_), .Y(_296__35_) );
AND2X2 AND2X2_120 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf2), .B(concatenador_data_out_36_), .Y(_296__36_) );
AND2X2 AND2X2_121 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf1), .B(concatenador_data_out_37_), .Y(_296__37_) );
AND2X2 AND2X2_122 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf0), .B(concatenador_data_out_38_), .Y(_296__38_) );
AND2X2 AND2X2_123 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf13), .B(concatenador_data_out_39_), .Y(_296__39_) );
AND2X2 AND2X2_124 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf12), .B(concatenador_data_out_48_), .Y(_296__48_) );
AND2X2 AND2X2_125 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf11), .B(concatenador_data_out_49_), .Y(_296__49_) );
AND2X2 AND2X2_126 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf10), .B(concatenador_data_out_50_), .Y(_296__50_) );
AND2X2 AND2X2_127 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf9), .B(concatenador_data_out_51_), .Y(_296__51_) );
AND2X2 AND2X2_128 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf8), .B(concatenador_data_out_52_), .Y(_296__52_) );
AND2X2 AND2X2_129 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf7), .B(concatenador_data_out_53_), .Y(_296__53_) );
AND2X2 AND2X2_130 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf6), .B(concatenador_data_out_54_), .Y(_296__54_) );
AND2X2 AND2X2_131 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf5), .B(concatenador_data_out_55_), .Y(_296__55_) );
AND2X2 AND2X2_132 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf4), .B(concatenador_data_out_40_), .Y(_296__40_) );
AND2X2 AND2X2_133 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf3), .B(concatenador_data_out_41_), .Y(_296__41_) );
AND2X2 AND2X2_134 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf2), .B(concatenador_data_out_42_), .Y(_296__42_) );
AND2X2 AND2X2_135 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf1), .B(concatenador_data_out_43_), .Y(_296__43_) );
AND2X2 AND2X2_136 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf0), .B(concatenador_data_out_44_), .Y(_296__44_) );
AND2X2 AND2X2_137 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf13), .B(concatenador_data_out_45_), .Y(_296__45_) );
AND2X2 AND2X2_138 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf12), .B(concatenador_data_out_46_), .Y(_296__46_) );
AND2X2 AND2X2_139 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf11), .B(concatenador_data_out_47_), .Y(_296__47_) );
AND2X2 AND2X2_140 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf10), .B(concatenador_data_out_8_), .Y(_296__8_) );
AND2X2 AND2X2_141 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf9), .B(concatenador_data_out_9_), .Y(_296__9_) );
AND2X2 AND2X2_142 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf8), .B(concatenador_data_out_10_), .Y(_296__10_) );
AND2X2 AND2X2_143 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf7), .B(concatenador_data_out_11_), .Y(_296__11_) );
AND2X2 AND2X2_144 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf6), .B(concatenador_data_out_12_), .Y(_296__12_) );
AND2X2 AND2X2_145 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf5), .B(concatenador_data_out_13_), .Y(_296__13_) );
AND2X2 AND2X2_146 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf4), .B(concatenador_data_out_14_), .Y(_296__14_) );
AND2X2 AND2X2_147 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf3), .B(concatenador_data_out_15_), .Y(_296__15_) );
AND2X2 AND2X2_148 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf2), .B(concatenador_data_out_24_), .Y(_296__24_) );
AND2X2 AND2X2_149 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf1), .B(concatenador_data_out_25_), .Y(_296__25_) );
AND2X2 AND2X2_150 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf0), .B(concatenador_data_out_26_), .Y(_296__26_) );
AND2X2 AND2X2_151 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf13), .B(concatenador_data_out_27_), .Y(_296__27_) );
AND2X2 AND2X2_152 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf12), .B(concatenador_data_out_28_), .Y(_296__28_) );
AND2X2 AND2X2_153 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf11), .B(concatenador_data_out_29_), .Y(_296__29_) );
AND2X2 AND2X2_154 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf10), .B(concatenador_data_out_30_), .Y(_296__30_) );
AND2X2 AND2X2_155 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf9), .B(concatenador_data_out_31_), .Y(_296__31_) );
AND2X2 AND2X2_156 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf8), .B(concatenador_data_out_16_), .Y(_296__16_) );
AND2X2 AND2X2_157 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf7), .B(concatenador_data_out_17_), .Y(_296__17_) );
AND2X2 AND2X2_158 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf6), .B(concatenador_data_out_18_), .Y(_296__18_) );
AND2X2 AND2X2_159 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf5), .B(concatenador_data_out_19_), .Y(_296__19_) );
AND2X2 AND2X2_160 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf4), .B(concatenador_data_out_20_), .Y(_296__20_) );
AND2X2 AND2X2_161 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf3), .B(concatenador_data_out_21_), .Y(_296__21_) );
AND2X2 AND2X2_162 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf2), .B(concatenador_data_out_22_), .Y(_296__22_) );
AND2X2 AND2X2_163 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf1), .B(concatenador_data_out_23_), .Y(_296__23_) );
INVX8 INVX8_16 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe69), .Y(_876_) );
NOR2X1 NOR2X1_163 ( .gnd(gnd), .vdd(vdd), .A(_876__bF_buf3), .B(_400__bF_buf5), .Y(_369_) );
AND2X2 AND2X2_164 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf0), .B(concatenador_data_out_0_), .Y(_296__0_) );
AND2X2 AND2X2_165 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf13), .B(concatenador_data_out_1_), .Y(_296__1_) );
AND2X2 AND2X2_166 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf12), .B(concatenador_data_out_2_), .Y(_296__2_) );
AND2X2 AND2X2_167 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf11), .B(concatenador_data_out_3_), .Y(_296__3_) );
AND2X2 AND2X2_168 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf10), .B(concatenador_data_out_4_), .Y(_296__4_) );
AND2X2 AND2X2_169 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf9), .B(concatenador_data_out_5_), .Y(_296__5_) );
AND2X2 AND2X2_170 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf8), .B(concatenador_data_out_6_), .Y(_296__6_) );
AND2X2 AND2X2_171 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf7), .B(concatenador_data_out_7_), .Y(_296__7_) );
NOR2X1 NOR2X1_164 ( .gnd(gnd), .vdd(vdd), .A(_4479__bF_buf1), .B(_400__bF_buf4), .Y(_370_) );
INVX8 INVX8_17 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe66_bF_buf4), .Y(_877_) );
NOR2X1 NOR2X1_165 ( .gnd(gnd), .vdd(vdd), .A(_877__bF_buf3), .B(_400__bF_buf3), .Y(_365_) );
INVX8 INVX8_18 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe68), .Y(_878_) );
NOR2X1 NOR2X1_166 ( .gnd(gnd), .vdd(vdd), .A(_878__bF_buf4), .B(_400__bF_buf2), .Y(_367_) );
INVX8 INVX8_19 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe67), .Y(_879_) );
NOR2X1 NOR2X1_167 ( .gnd(gnd), .vdd(vdd), .A(_879__bF_buf3), .B(_400__bF_buf1), .Y(_366_) );
INVX8 INVX8_20 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe63), .Y(_880_) );
NOR2X1 NOR2X1_168 ( .gnd(gnd), .vdd(vdd), .A(_880__bF_buf3), .B(_400__bF_buf0), .Y(_362_) );
INVX8 INVX8_21 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe65_bF_buf3), .Y(_881_) );
NOR2X1 NOR2X1_169 ( .gnd(gnd), .vdd(vdd), .A(_881_), .B(_400__bF_buf12), .Y(_364_) );
INVX8 INVX8_22 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe64_bF_buf4), .Y(_882_) );
NOR2X1 NOR2X1_170 ( .gnd(gnd), .vdd(vdd), .A(_882__bF_buf3), .B(_400__bF_buf11), .Y(_363_) );
INVX8 INVX8_23 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe60_bF_buf4), .Y(_883_) );
NOR2X1 NOR2X1_171 ( .gnd(gnd), .vdd(vdd), .A(_883__bF_buf3), .B(_400__bF_buf10), .Y(_359_) );
INVX8 INVX8_24 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe62_bF_buf4), .Y(_884_) );
NOR2X1 NOR2X1_172 ( .gnd(gnd), .vdd(vdd), .A(_884__bF_buf4), .B(_400__bF_buf9), .Y(_361_) );
INVX8 INVX8_25 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe61_bF_buf3), .Y(_885_) );
NOR2X1 NOR2X1_173 ( .gnd(gnd), .vdd(vdd), .A(_885_), .B(_400__bF_buf8), .Y(_360_) );
INVX8 INVX8_26 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe57_bF_buf3), .Y(_886_) );
NOR2X1 NOR2X1_174 ( .gnd(gnd), .vdd(vdd), .A(_886_), .B(_400__bF_buf7), .Y(_355_) );
INVX8 INVX8_27 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe59), .Y(_887_) );
NOR2X1 NOR2X1_175 ( .gnd(gnd), .vdd(vdd), .A(_887__bF_buf3), .B(_400__bF_buf6), .Y(_358_) );
INVX8 INVX8_28 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe58_bF_buf4), .Y(_888_) );
NOR2X1 NOR2X1_176 ( .gnd(gnd), .vdd(vdd), .A(_888__bF_buf3), .B(_400__bF_buf5), .Y(_356_) );
INVX8 INVX8_29 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe54_bF_buf3), .Y(_889_) );
NOR2X1 NOR2X1_177 ( .gnd(gnd), .vdd(vdd), .A(_889__bF_buf4), .B(_400__bF_buf4), .Y(_352_) );
INVX8 INVX8_30 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe56_bF_buf3), .Y(_890_) );
NOR2X1 NOR2X1_178 ( .gnd(gnd), .vdd(vdd), .A(_890__bF_buf4), .B(_400__bF_buf3), .Y(_354_) );
INVX8 INVX8_31 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe55), .Y(_891_) );
NOR2X1 NOR2X1_179 ( .gnd(gnd), .vdd(vdd), .A(_891_), .B(_400__bF_buf2), .Y(_353_) );
INVX8 INVX8_32 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe51), .Y(_892_) );
NOR2X1 NOR2X1_180 ( .gnd(gnd), .vdd(vdd), .A(_892_), .B(_400__bF_buf1), .Y(_349_) );
INVX8 INVX8_33 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe53_bF_buf3), .Y(_893_) );
NOR2X1 NOR2X1_181 ( .gnd(gnd), .vdd(vdd), .A(_893_), .B(_400__bF_buf0), .Y(_351_) );
INVX8 INVX8_34 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe52_bF_buf4), .Y(_894_) );
NOR2X1 NOR2X1_182 ( .gnd(gnd), .vdd(vdd), .A(_894__bF_buf3), .B(_400__bF_buf12), .Y(_350_) );
INVX8 INVX8_35 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe48_bF_buf3), .Y(_895_) );
NOR2X1 NOR2X1_183 ( .gnd(gnd), .vdd(vdd), .A(_895__bF_buf4), .B(_400__bF_buf11), .Y(_345_) );
INVX8 INVX8_36 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe50_bF_buf3), .Y(_896_) );
NOR2X1 NOR2X1_184 ( .gnd(gnd), .vdd(vdd), .A(_896__bF_buf4), .B(_400__bF_buf10), .Y(_348_) );
INVX8 INVX8_37 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe49), .Y(_897_) );
NOR2X1 NOR2X1_185 ( .gnd(gnd), .vdd(vdd), .A(_897__bF_buf3), .B(_400__bF_buf9), .Y(_347_) );
INVX8 INVX8_38 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe45_bF_buf3), .Y(_898_) );
NOR2X1 NOR2X1_186 ( .gnd(gnd), .vdd(vdd), .A(_898_), .B(_400__bF_buf8), .Y(_342_) );
INVX8 INVX8_39 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe47), .Y(_899_) );
NOR2X1 NOR2X1_187 ( .gnd(gnd), .vdd(vdd), .A(_899__bF_buf3), .B(_400__bF_buf7), .Y(_344_) );
INVX8 INVX8_40 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe46_bF_buf4), .Y(_900_) );
NOR2X1 NOR2X1_188 ( .gnd(gnd), .vdd(vdd), .A(_900__bF_buf3), .B(_400__bF_buf6), .Y(_343_) );
INVX8 INVX8_41 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe42_bF_buf3), .Y(_901_) );
NOR2X1 NOR2X1_189 ( .gnd(gnd), .vdd(vdd), .A(_901__bF_buf4), .B(_400__bF_buf5), .Y(_339_) );
INVX8 INVX8_42 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe44), .Y(_902_) );
NOR2X1 NOR2X1_190 ( .gnd(gnd), .vdd(vdd), .A(_902__bF_buf4), .B(_400__bF_buf4), .Y(_341_) );
INVX8 INVX8_43 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe43), .Y(_903_) );
NOR2X1 NOR2X1_191 ( .gnd(gnd), .vdd(vdd), .A(_903__bF_buf3), .B(_400__bF_buf3), .Y(_340_) );
INVX8 INVX8_44 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe39), .Y(_904_) );
NOR2X1 NOR2X1_192 ( .gnd(gnd), .vdd(vdd), .A(_904__bF_buf3), .B(_400__bF_buf2), .Y(_336_) );
INVX8 INVX8_45 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe41), .Y(_905_) );
NOR2X1 NOR2X1_193 ( .gnd(gnd), .vdd(vdd), .A(_905__bF_buf3), .B(_400__bF_buf1), .Y(_338_) );
INVX8 INVX8_46 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe40_bF_buf4), .Y(_906_) );
NOR2X1 NOR2X1_194 ( .gnd(gnd), .vdd(vdd), .A(_906__bF_buf4), .B(_400__bF_buf0), .Y(_337_) );
INVX8 INVX8_47 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe36_bF_buf3), .Y(_907_) );
NOR2X1 NOR2X1_195 ( .gnd(gnd), .vdd(vdd), .A(_907__bF_buf4), .B(_400__bF_buf12), .Y(_332_) );
INVX8 INVX8_48 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe38_bF_buf3), .Y(_908_) );
NOR2X1 NOR2X1_196 ( .gnd(gnd), .vdd(vdd), .A(_908__bF_buf4), .B(_400__bF_buf11), .Y(_334_) );
INVX8 INVX8_49 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe37), .Y(_909_) );
NOR2X1 NOR2X1_197 ( .gnd(gnd), .vdd(vdd), .A(_909__bF_buf3), .B(_400__bF_buf10), .Y(_333_) );
INVX8 INVX8_50 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe33_bF_buf3), .Y(_910_) );
NOR2X1 NOR2X1_198 ( .gnd(gnd), .vdd(vdd), .A(_910_), .B(_400__bF_buf9), .Y(_329_) );
INVX8 INVX8_51 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe35), .Y(_911_) );
NOR2X1 NOR2X1_199 ( .gnd(gnd), .vdd(vdd), .A(_911__bF_buf4), .B(_400__bF_buf8), .Y(_331_) );
INVX8 INVX8_52 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe34_bF_buf3), .Y(_912_) );
NOR2X1 NOR2X1_200 ( .gnd(gnd), .vdd(vdd), .A(_912__bF_buf4), .B(_400__bF_buf7), .Y(_330_) );
INVX8 INVX8_53 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe30_bF_buf3), .Y(_913_) );
NOR2X1 NOR2X1_201 ( .gnd(gnd), .vdd(vdd), .A(_913__bF_buf4), .B(_400__bF_buf6), .Y(_326_) );
INVX8 INVX8_54 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe32_bF_buf3), .Y(_914_) );
NOR2X1 NOR2X1_202 ( .gnd(gnd), .vdd(vdd), .A(_914__bF_buf4), .B(_400__bF_buf5), .Y(_328_) );
INVX8 INVX8_55 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe31), .Y(_915_) );
NOR2X1 NOR2X1_203 ( .gnd(gnd), .vdd(vdd), .A(_915__bF_buf3), .B(_400__bF_buf4), .Y(_327_) );
INVX8 INVX8_56 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe27), .Y(_916_) );
NOR2X1 NOR2X1_204 ( .gnd(gnd), .vdd(vdd), .A(_916_), .B(_400__bF_buf3), .Y(_322_) );
INVX8 INVX8_57 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe29_bF_buf3), .Y(_917_) );
NOR2X1 NOR2X1_205 ( .gnd(gnd), .vdd(vdd), .A(_917_), .B(_400__bF_buf2), .Y(_325_) );
INVX8 INVX8_58 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe28_bF_buf3), .Y(_918_) );
NOR2X1 NOR2X1_206 ( .gnd(gnd), .vdd(vdd), .A(_918__bF_buf4), .B(_400__bF_buf1), .Y(_323_) );
INVX8 INVX8_59 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe24_bF_buf4), .Y(_919_) );
NOR2X1 NOR2X1_207 ( .gnd(gnd), .vdd(vdd), .A(_919__bF_buf4), .B(_400__bF_buf0), .Y(_319_) );
INVX8 INVX8_60 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe26_bF_buf3), .Y(_920_) );
NOR2X1 NOR2X1_208 ( .gnd(gnd), .vdd(vdd), .A(_920__bF_buf4), .B(_400__bF_buf12), .Y(_321_) );
INVX8 INVX8_61 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe25), .Y(_921_) );
NOR2X1 NOR2X1_209 ( .gnd(gnd), .vdd(vdd), .A(_921__bF_buf3), .B(_400__bF_buf11), .Y(_320_) );
INVX8 INVX8_62 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe21_bF_buf3), .Y(_922_) );
NOR2X1 NOR2X1_210 ( .gnd(gnd), .vdd(vdd), .A(_922_), .B(_400__bF_buf10), .Y(_316_) );
INVX8 INVX8_63 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe23_bF_buf3), .Y(_923_) );
NOR2X1 NOR2X1_211 ( .gnd(gnd), .vdd(vdd), .A(_923_), .B(_400__bF_buf9), .Y(_318_) );
INVX8 INVX8_64 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe22_bF_buf4), .Y(_924_) );
NOR2X1 NOR2X1_212 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf4), .B(_400__bF_buf8), .Y(_317_) );
INVX8 INVX8_65 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe18_bF_buf4), .Y(_925_) );
NOR2X1 NOR2X1_213 ( .gnd(gnd), .vdd(vdd), .A(_925__bF_buf4), .B(_400__bF_buf7), .Y(_312_) );
INVX8 INVX8_66 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe20_bF_buf4), .Y(_926_) );
NOR2X1 NOR2X1_214 ( .gnd(gnd), .vdd(vdd), .A(_926__bF_buf4), .B(_400__bF_buf6), .Y(_315_) );
INVX8 INVX8_67 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe19_bF_buf3), .Y(_927_) );
NOR2X1 NOR2X1_215 ( .gnd(gnd), .vdd(vdd), .A(_927__bF_buf3), .B(_400__bF_buf5), .Y(_314_) );
INVX8 INVX8_68 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe15_bF_buf3), .Y(_928_) );
NOR2X1 NOR2X1_216 ( .gnd(gnd), .vdd(vdd), .A(_928_), .B(_400__bF_buf4), .Y(_309_) );
INVX8 INVX8_69 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe17_bF_buf3), .Y(_929_) );
NOR2X1 NOR2X1_217 ( .gnd(gnd), .vdd(vdd), .A(_929_), .B(_400__bF_buf3), .Y(_311_) );
INVX8 INVX8_70 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe16_bF_buf3), .Y(_930_) );
NOR2X1 NOR2X1_218 ( .gnd(gnd), .vdd(vdd), .A(_930__bF_buf4), .B(_400__bF_buf2), .Y(_310_) );
INVX8 INVX8_71 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe12), .Y(_931_) );
NOR2X1 NOR2X1_219 ( .gnd(gnd), .vdd(vdd), .A(_931_), .B(_400__bF_buf1), .Y(_306_) );
INVX8 INVX8_72 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe14_bF_buf4), .Y(_932_) );
NOR2X1 NOR2X1_220 ( .gnd(gnd), .vdd(vdd), .A(_932_), .B(_400__bF_buf0), .Y(_308_) );
INVX4 INVX4_48 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe13), .Y(_933_) );
NOR2X1 NOR2X1_221 ( .gnd(gnd), .vdd(vdd), .A(_933_), .B(_400__bF_buf12), .Y(_307_) );
INVX2 INVX2_92 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe9), .Y(_934_) );
NOR2X1 NOR2X1_222 ( .gnd(gnd), .vdd(vdd), .A(_934_), .B(_400__bF_buf11), .Y(_303_) );
INVX2 INVX2_93 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe11), .Y(_935_) );
NOR2X1 NOR2X1_223 ( .gnd(gnd), .vdd(vdd), .A(_935_), .B(_400__bF_buf10), .Y(_305_) );
INVX8 INVX8_73 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe10), .Y(_936_) );
NOR2X1 NOR2X1_224 ( .gnd(gnd), .vdd(vdd), .A(_936_), .B(_400__bF_buf9), .Y(_304_) );
INVX4 INVX4_49 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe6), .Y(_937_) );
NOR2X1 NOR2X1_225 ( .gnd(gnd), .vdd(vdd), .A(_937_), .B(_400__bF_buf8), .Y(_371_) );
INVX4 INVX4_50 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe8), .Y(_938_) );
NOR2X1 NOR2X1_226 ( .gnd(gnd), .vdd(vdd), .A(_938_), .B(_400__bF_buf7), .Y(_373_) );
INVX4 INVX4_51 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe7), .Y(_939_) );
NOR2X1 NOR2X1_227 ( .gnd(gnd), .vdd(vdd), .A(_939_), .B(_400__bF_buf6), .Y(_372_) );
AND2X2 AND2X2_172 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf6), .B(micro_hash_ucr_pipe3), .Y(_346_) );
AND2X2 AND2X2_173 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf5), .B(micro_hash_ucr_pipe5), .Y(_368_) );
AND2X2 AND2X2_174 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf4), .B(micro_hash_ucr_pipe4), .Y(_357_) );
AND2X2 AND2X2_175 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf3), .B(micro_hash_ucr_pipe0), .Y(_313_) );
AND2X2 AND2X2_176 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf2), .B(micro_hash_ucr_pipe2), .Y(_335_) );
AND2X2 AND2X2_177 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf1), .B(micro_hash_ucr_pipe1), .Y(_324_) );
NAND2X1 NAND2X1_69 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe58_bF_buf3), .B(_436_), .Y(_940_) );
NAND2X1 NAND2X1_70 ( .gnd(gnd), .vdd(vdd), .A(_4423__bF_buf1), .B(_4481_), .Y(_941_) );
NAND2X1 NAND2X1_71 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_0_bF_buf1_), .B(micro_hash_ucr_b_0_bF_buf1_), .Y(_942_) );
NAND2X1 NAND2X1_72 ( .gnd(gnd), .vdd(vdd), .A(_942_), .B(_941_), .Y(_943_) );
INVX8 INVX8_74 ( .gnd(gnd), .vdd(vdd), .A(_943_), .Y(_944_) );
NOR2X1 NOR2X1_228 ( .gnd(gnd), .vdd(vdd), .A(_917_), .B(_944__bF_buf3), .Y(_945_) );
NAND2X1 NAND2X1_73 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe27), .B(_944__bF_buf2), .Y(_946_) );
AOI21X1 AOI21X1_178 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe12), .B(_933_), .C(micro_hash_ucr_pipe14_bF_buf3), .Y(_947_) );
OAI21X1 OAI21X1_207 ( .gnd(gnd), .vdd(vdd), .A(_947_), .B(micro_hash_ucr_pipe15_bF_buf2), .C(_930__bF_buf3), .Y(_948_) );
AOI21X1 AOI21X1_179 ( .gnd(gnd), .vdd(vdd), .A(_929_), .B(_948_), .C(micro_hash_ucr_pipe18_bF_buf3), .Y(_949_) );
OAI21X1 OAI21X1_208 ( .gnd(gnd), .vdd(vdd), .A(_949_), .B(micro_hash_ucr_pipe19_bF_buf2), .C(_926__bF_buf3), .Y(_950_) );
AOI21X1 AOI21X1_180 ( .gnd(gnd), .vdd(vdd), .A(_922_), .B(_950_), .C(micro_hash_ucr_pipe22_bF_buf3), .Y(_951_) );
OAI21X1 OAI21X1_209 ( .gnd(gnd), .vdd(vdd), .A(_951_), .B(micro_hash_ucr_pipe23_bF_buf2), .C(_919__bF_buf3), .Y(_952_) );
NAND2X1 NAND2X1_74 ( .gnd(gnd), .vdd(vdd), .A(_921__bF_buf2), .B(_952_), .Y(_953_) );
NAND2X1 NAND2X1_75 ( .gnd(gnd), .vdd(vdd), .A(_920__bF_buf3), .B(_953_), .Y(_954_) );
OAI21X1 OAI21X1_210 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe6), .B(micro_hash_ucr_pipe7), .C(_938_), .Y(_955_) );
AOI21X1 AOI21X1_181 ( .gnd(gnd), .vdd(vdd), .A(_934_), .B(_955_), .C(micro_hash_ucr_pipe10), .Y(_956_) );
OAI21X1 OAI21X1_211 ( .gnd(gnd), .vdd(vdd), .A(_956_), .B(micro_hash_ucr_pipe11), .C(_931_), .Y(_957_) );
NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_926__bF_buf2), .B(_930__bF_buf2), .C(_932_), .Y(_958_) );
NOR2X1 NOR2X1_229 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe24_bF_buf3), .B(micro_hash_ucr_pipe26_bF_buf2), .Y(_959_) );
NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf3), .B(_925__bF_buf3), .C(_959_), .Y(_960_) );
OR2X2 OR2X2_24 ( .gnd(gnd), .vdd(vdd), .A(_960_), .B(_958_), .Y(_961_) );
NOR2X1 NOR2X1_230 ( .gnd(gnd), .vdd(vdd), .A(_961_), .B(_957_), .Y(_962_) );
NOR2X1 NOR2X1_231 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_0_bF_buf1_), .B(_962_), .Y(_963_) );
NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe6), .B(_936_), .C(_938_), .Y(_964_) );
NOR2X1 NOR2X1_232 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe9), .B(micro_hash_ucr_pipe7), .Y(_965_) );
NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_434_), .B(_935_), .C(_965_), .Y(_966_) );
OAI21X1 OAI21X1_212 ( .gnd(gnd), .vdd(vdd), .A(_939_), .B(micro_hash_ucr_pipe8), .C(_934_), .Y(_967_) );
AOI21X1 AOI21X1_182 ( .gnd(gnd), .vdd(vdd), .A(_936_), .B(_967_), .C(micro_hash_ucr_pipe11), .Y(_968_) );
INVX1 INVX1_101 ( .gnd(gnd), .vdd(vdd), .A(_968_), .Y(_969_) );
NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_922_), .B(_927__bF_buf2), .C(_933_), .Y(_970_) );
NOR2X1 NOR2X1_233 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe15_bF_buf1), .B(micro_hash_ucr_pipe17_bF_buf2), .Y(_971_) );
NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_921__bF_buf1), .B(_923_), .C(_971_), .Y(_972_) );
OR2X2 OR2X2_25 ( .gnd(gnd), .vdd(vdd), .A(_972_), .B(_970_), .Y(_973_) );
OAI21X1 OAI21X1_213 ( .gnd(gnd), .vdd(vdd), .A(_969_), .B(_973_), .C(_943_), .Y(_974_) );
OAI21X1 OAI21X1_214 ( .gnd(gnd), .vdd(vdd), .A(_964_), .B(_966_), .C(_974_), .Y(_975_) );
AOI21X1 AOI21X1_183 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe13), .B(_932_), .C(micro_hash_ucr_pipe15_bF_buf0), .Y(_976_) );
OAI21X1 OAI21X1_215 ( .gnd(gnd), .vdd(vdd), .A(_976_), .B(micro_hash_ucr_pipe16_bF_buf2), .C(_929_), .Y(_977_) );
AOI21X1 AOI21X1_184 ( .gnd(gnd), .vdd(vdd), .A(_925__bF_buf2), .B(_977_), .C(micro_hash_ucr_pipe19_bF_buf1), .Y(_978_) );
OAI21X1 OAI21X1_216 ( .gnd(gnd), .vdd(vdd), .A(_978_), .B(micro_hash_ucr_pipe20_bF_buf3), .C(_922_), .Y(_979_) );
AOI21X1 AOI21X1_185 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf2), .B(_979_), .C(micro_hash_ucr_pipe23_bF_buf1), .Y(_980_) );
OAI21X1 OAI21X1_217 ( .gnd(gnd), .vdd(vdd), .A(_980_), .B(micro_hash_ucr_pipe24_bF_buf2), .C(_921__bF_buf0), .Y(_981_) );
NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_920__bF_buf2), .B(_944__bF_buf1), .C(_981_), .Y(_982_) );
OAI21X1 OAI21X1_218 ( .gnd(gnd), .vdd(vdd), .A(_963_), .B(_975_), .C(_982_), .Y(_983_) );
AOI21X1 AOI21X1_186 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_0_bF_buf0_), .B(_954_), .C(_983_), .Y(_984_) );
OAI21X1 OAI21X1_219 ( .gnd(gnd), .vdd(vdd), .A(_984_), .B(micro_hash_ucr_pipe27), .C(_946_), .Y(_985_) );
OAI21X1 OAI21X1_220 ( .gnd(gnd), .vdd(vdd), .A(_436_), .B(_918__bF_buf3), .C(_917_), .Y(_986_) );
AOI21X1 AOI21X1_187 ( .gnd(gnd), .vdd(vdd), .A(_918__bF_buf2), .B(_985_), .C(_986_), .Y(_987_) );
OAI21X1 OAI21X1_221 ( .gnd(gnd), .vdd(vdd), .A(_987_), .B(_945_), .C(_913__bF_buf3), .Y(_988_) );
AOI21X1 AOI21X1_188 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe30_bF_buf2), .B(_436_), .C(micro_hash_ucr_pipe31), .Y(_989_) );
OAI21X1 OAI21X1_222 ( .gnd(gnd), .vdd(vdd), .A(_943_), .B(_915__bF_buf2), .C(_914__bF_buf3), .Y(_990_) );
AOI21X1 AOI21X1_189 ( .gnd(gnd), .vdd(vdd), .A(_989_), .B(_988_), .C(_990_), .Y(_991_) );
NOR2X1 NOR2X1_234 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_0_bF_buf3_), .B(_914__bF_buf2), .Y(_992_) );
OAI21X1 OAI21X1_223 ( .gnd(gnd), .vdd(vdd), .A(_991_), .B(_992_), .C(_910_), .Y(_993_) );
OAI21X1 OAI21X1_224 ( .gnd(gnd), .vdd(vdd), .A(_910_), .B(_944__bF_buf0), .C(_993_), .Y(_994_) );
NAND2X1 NAND2X1_76 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_0_bF_buf2_), .B(micro_hash_ucr_pipe34_bF_buf2), .Y(_995_) );
OAI21X1 OAI21X1_225 ( .gnd(gnd), .vdd(vdd), .A(_994_), .B(micro_hash_ucr_pipe34_bF_buf1), .C(_995_), .Y(_996_) );
NAND2X1 NAND2X1_77 ( .gnd(gnd), .vdd(vdd), .A(_911__bF_buf3), .B(_996_), .Y(_997_) );
OAI21X1 OAI21X1_226 ( .gnd(gnd), .vdd(vdd), .A(_911__bF_buf2), .B(_943_), .C(_997_), .Y(_998_) );
AOI21X1 AOI21X1_190 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe36_bF_buf2), .B(_436_), .C(micro_hash_ucr_pipe37), .Y(_999_) );
OAI21X1 OAI21X1_227 ( .gnd(gnd), .vdd(vdd), .A(_998_), .B(micro_hash_ucr_pipe36_bF_buf1), .C(_999_), .Y(_1000_) );
OAI21X1 OAI21X1_228 ( .gnd(gnd), .vdd(vdd), .A(_909__bF_buf2), .B(_943_), .C(_1000_), .Y(_1001_) );
NAND2X1 NAND2X1_78 ( .gnd(gnd), .vdd(vdd), .A(_908__bF_buf3), .B(_1001_), .Y(_1002_) );
OAI21X1 OAI21X1_229 ( .gnd(gnd), .vdd(vdd), .A(_436_), .B(_908__bF_buf2), .C(_1002_), .Y(_1003_) );
OAI21X1 OAI21X1_230 ( .gnd(gnd), .vdd(vdd), .A(_943_), .B(_904__bF_buf2), .C(_906__bF_buf3), .Y(_1004_) );
AOI21X1 AOI21X1_191 ( .gnd(gnd), .vdd(vdd), .A(_904__bF_buf1), .B(_1003_), .C(_1004_), .Y(_1005_) );
OAI21X1 OAI21X1_231 ( .gnd(gnd), .vdd(vdd), .A(_906__bF_buf2), .B(micro_hash_ucr_a_0_bF_buf1_), .C(_905__bF_buf2), .Y(_1006_) );
AOI21X1 AOI21X1_192 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe41), .B(_944__bF_buf3), .C(micro_hash_ucr_pipe42_bF_buf2), .Y(_1007_) );
OAI21X1 OAI21X1_232 ( .gnd(gnd), .vdd(vdd), .A(_1005_), .B(_1006_), .C(_1007_), .Y(_1008_) );
OAI21X1 OAI21X1_233 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_0_bF_buf0_), .B(_901__bF_buf3), .C(_1008_), .Y(_1009_) );
AND2X2 AND2X2_178 ( .gnd(gnd), .vdd(vdd), .A(_1009_), .B(_903__bF_buf2), .Y(_1010_) );
NOR2X1 NOR2X1_235 ( .gnd(gnd), .vdd(vdd), .A(_903__bF_buf1), .B(_944__bF_buf2), .Y(_1011_) );
OAI21X1 OAI21X1_234 ( .gnd(gnd), .vdd(vdd), .A(_1010_), .B(_1011_), .C(_902__bF_buf3), .Y(_1012_) );
OAI21X1 OAI21X1_235 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_0_bF_buf3_), .B(_902__bF_buf2), .C(_1012_), .Y(_1013_) );
AND2X2 AND2X2_179 ( .gnd(gnd), .vdd(vdd), .A(_1013_), .B(_898_), .Y(_1014_) );
NOR2X1 NOR2X1_236 ( .gnd(gnd), .vdd(vdd), .A(_898_), .B(_944__bF_buf1), .Y(_1015_) );
OAI21X1 OAI21X1_236 ( .gnd(gnd), .vdd(vdd), .A(_1014_), .B(_1015_), .C(_900__bF_buf2), .Y(_1016_) );
OAI21X1 OAI21X1_237 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_0_bF_buf2_), .B(_900__bF_buf1), .C(_1016_), .Y(_1017_) );
AND2X2 AND2X2_180 ( .gnd(gnd), .vdd(vdd), .A(_1017_), .B(_899__bF_buf2), .Y(_1018_) );
NOR2X1 NOR2X1_237 ( .gnd(gnd), .vdd(vdd), .A(_899__bF_buf1), .B(_944__bF_buf0), .Y(_1019_) );
OAI21X1 OAI21X1_238 ( .gnd(gnd), .vdd(vdd), .A(_1018_), .B(_1019_), .C(_895__bF_buf3), .Y(_1020_) );
OAI21X1 OAI21X1_239 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_0_bF_buf1_), .B(_895__bF_buf2), .C(_1020_), .Y(_1021_) );
AND2X2 AND2X2_181 ( .gnd(gnd), .vdd(vdd), .A(_1021_), .B(_897__bF_buf2), .Y(_1022_) );
NOR2X1 NOR2X1_238 ( .gnd(gnd), .vdd(vdd), .A(_897__bF_buf1), .B(_944__bF_buf3), .Y(_1023_) );
OAI21X1 OAI21X1_240 ( .gnd(gnd), .vdd(vdd), .A(_1022_), .B(_1023_), .C(_896__bF_buf3), .Y(_1024_) );
OAI21X1 OAI21X1_241 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_0_bF_buf0_), .B(_896__bF_buf2), .C(_1024_), .Y(_1025_) );
AND2X2 AND2X2_182 ( .gnd(gnd), .vdd(vdd), .A(_1025_), .B(_892_), .Y(_1026_) );
NOR2X1 NOR2X1_239 ( .gnd(gnd), .vdd(vdd), .A(_892_), .B(_944__bF_buf2), .Y(_1027_) );
OAI21X1 OAI21X1_242 ( .gnd(gnd), .vdd(vdd), .A(_1026_), .B(_1027_), .C(_894__bF_buf2), .Y(_1028_) );
OAI21X1 OAI21X1_243 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_0_bF_buf3_), .B(_894__bF_buf1), .C(_1028_), .Y(_1029_) );
AND2X2 AND2X2_183 ( .gnd(gnd), .vdd(vdd), .A(_1029_), .B(_893_), .Y(_1030_) );
NOR2X1 NOR2X1_240 ( .gnd(gnd), .vdd(vdd), .A(_893_), .B(_944__bF_buf1), .Y(_1031_) );
OAI21X1 OAI21X1_244 ( .gnd(gnd), .vdd(vdd), .A(_1030_), .B(_1031_), .C(_889__bF_buf3), .Y(_1032_) );
OAI21X1 OAI21X1_245 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_0_bF_buf2_), .B(_889__bF_buf2), .C(_1032_), .Y(_1033_) );
AND2X2 AND2X2_184 ( .gnd(gnd), .vdd(vdd), .A(_1033_), .B(_891_), .Y(_1034_) );
NOR2X1 NOR2X1_241 ( .gnd(gnd), .vdd(vdd), .A(_891_), .B(_944__bF_buf0), .Y(_1035_) );
OAI21X1 OAI21X1_246 ( .gnd(gnd), .vdd(vdd), .A(_1034_), .B(_1035_), .C(_890__bF_buf3), .Y(_1036_) );
OAI21X1 OAI21X1_247 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_0_bF_buf1_), .B(_890__bF_buf2), .C(_1036_), .Y(_1037_) );
AND2X2 AND2X2_185 ( .gnd(gnd), .vdd(vdd), .A(_1037_), .B(_886_), .Y(_1038_) );
NOR2X1 NOR2X1_242 ( .gnd(gnd), .vdd(vdd), .A(_886_), .B(_944__bF_buf3), .Y(_1039_) );
OAI21X1 OAI21X1_248 ( .gnd(gnd), .vdd(vdd), .A(_1038_), .B(_1039_), .C(_888__bF_buf2), .Y(_1040_) );
NAND3X1 NAND3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_887__bF_buf2), .B(_940_), .C(_1040_), .Y(_1041_) );
AOI21X1 AOI21X1_193 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe59), .B(_944__bF_buf2), .C(micro_hash_ucr_pipe60_bF_buf3), .Y(_1042_) );
OAI21X1 OAI21X1_249 ( .gnd(gnd), .vdd(vdd), .A(_883__bF_buf2), .B(micro_hash_ucr_a_0_bF_buf0_), .C(_885_), .Y(_1043_) );
AOI21X1 AOI21X1_194 ( .gnd(gnd), .vdd(vdd), .A(_1042_), .B(_1041_), .C(_1043_), .Y(_1044_) );
OAI21X1 OAI21X1_250 ( .gnd(gnd), .vdd(vdd), .A(_943_), .B(_885_), .C(_884__bF_buf3), .Y(_1045_) );
OAI22X1 OAI22X1_19 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_0_bF_buf3_), .B(_884__bF_buf2), .C(_1044_), .D(_1045_), .Y(_1046_) );
OAI21X1 OAI21X1_251 ( .gnd(gnd), .vdd(vdd), .A(_944__bF_buf1), .B(_880__bF_buf2), .C(_882__bF_buf2), .Y(_1047_) );
AOI21X1 AOI21X1_195 ( .gnd(gnd), .vdd(vdd), .A(_880__bF_buf1), .B(_1046_), .C(_1047_), .Y(_1048_) );
NOR2X1 NOR2X1_243 ( .gnd(gnd), .vdd(vdd), .A(_436_), .B(_882__bF_buf1), .Y(_1049_) );
OAI21X1 OAI21X1_252 ( .gnd(gnd), .vdd(vdd), .A(_1048_), .B(_1049_), .C(_881_), .Y(_1050_) );
AOI21X1 AOI21X1_196 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe65_bF_buf2), .B(_944__bF_buf0), .C(micro_hash_ucr_pipe66_bF_buf3), .Y(_1051_) );
OAI21X1 OAI21X1_253 ( .gnd(gnd), .vdd(vdd), .A(_877__bF_buf2), .B(micro_hash_ucr_a_0_bF_buf2_), .C(_879__bF_buf2), .Y(_1052_) );
AOI21X1 AOI21X1_197 ( .gnd(gnd), .vdd(vdd), .A(_1051_), .B(_1050_), .C(_1052_), .Y(_1053_) );
OAI21X1 OAI21X1_254 ( .gnd(gnd), .vdd(vdd), .A(_943_), .B(_879__bF_buf1), .C(_878__bF_buf3), .Y(_1054_) );
OAI22X1 OAI22X1_20 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_0_bF_buf1_), .B(_878__bF_buf2), .C(_1053_), .D(_1054_), .Y(_1055_) );
OAI21X1 OAI21X1_255 ( .gnd(gnd), .vdd(vdd), .A(_944__bF_buf3), .B(_876__bF_buf2), .C(_302__bF_buf0), .Y(_1056_) );
AOI21X1 AOI21X1_198 ( .gnd(gnd), .vdd(vdd), .A(_876__bF_buf1), .B(_1055_), .C(_1056_), .Y(_297__0_) );
NOR2X1 NOR2X1_244 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_1_bF_buf1_), .B(micro_hash_ucr_b_1_bF_buf1_), .Y(_1057_) );
INVX8 INVX8_75 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_1_bF_buf0_), .Y(_1058_) );
NOR2X1 NOR2X1_245 ( .gnd(gnd), .vdd(vdd), .A(_1058__bF_buf3), .B(_4487_), .Y(_1059_) );
NOR2X1 NOR2X1_246 ( .gnd(gnd), .vdd(vdd), .A(_1057_), .B(_1059_), .Y(_1060_) );
INVX8 INVX8_76 ( .gnd(gnd), .vdd(vdd), .A(_1060_), .Y(_1061_) );
NOR2X1 NOR2X1_247 ( .gnd(gnd), .vdd(vdd), .A(_442_), .B(_884__bF_buf1), .Y(_1062_) );
NAND2X1 NAND2X1_79 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_1_), .B(micro_hash_ucr_pipe58_bF_buf2), .Y(_1063_) );
NAND2X1 NAND2X1_80 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_1_), .B(micro_hash_ucr_pipe56_bF_buf2), .Y(_1064_) );
NAND2X1 NAND2X1_81 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_1_), .B(micro_hash_ucr_pipe54_bF_buf2), .Y(_1065_) );
NAND2X1 NAND2X1_82 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_1_), .B(micro_hash_ucr_pipe52_bF_buf3), .Y(_1066_) );
NOR2X1 NOR2X1_248 ( .gnd(gnd), .vdd(vdd), .A(_442_), .B(_900__bF_buf0), .Y(_1067_) );
NAND2X1 NAND2X1_83 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe38_bF_buf2), .B(_442_), .Y(_1068_) );
NAND2X1 NAND2X1_84 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_1_), .B(micro_hash_ucr_pipe28_bF_buf2), .Y(_1069_) );
AOI21X1 AOI21X1_199 ( .gnd(gnd), .vdd(vdd), .A(_931_), .B(_969_), .C(micro_hash_ucr_pipe13), .Y(_1070_) );
OAI21X1 OAI21X1_256 ( .gnd(gnd), .vdd(vdd), .A(_1070_), .B(micro_hash_ucr_pipe14_bF_buf2), .C(_928_), .Y(_1071_) );
NAND2X1 NAND2X1_85 ( .gnd(gnd), .vdd(vdd), .A(_934_), .B(_935_), .Y(_1072_) );
NOR2X1 NOR2X1_249 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe12), .B(micro_hash_ucr_pipe14_bF_buf1), .Y(_1073_) );
NAND3X1 NAND3X1_18 ( .gnd(gnd), .vdd(vdd), .A(H_1_), .B(_928_), .C(_1073_), .Y(_1074_) );
NOR2X1 NOR2X1_250 ( .gnd(gnd), .vdd(vdd), .A(_1072_), .B(_1074_), .Y(_1075_) );
NAND3X1 NAND3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_933_), .B(_936_), .C(_939_), .Y(_1076_) );
NOR2X1 NOR2X1_251 ( .gnd(gnd), .vdd(vdd), .A(_955_), .B(_1076_), .Y(_1077_) );
AOI22X1 AOI22X1_13 ( .gnd(gnd), .vdd(vdd), .A(_1075_), .B(_1077_), .C(_1071_), .D(_1060_), .Y(_1078_) );
AOI21X1 AOI21X1_200 ( .gnd(gnd), .vdd(vdd), .A(_933_), .B(_957_), .C(micro_hash_ucr_pipe14_bF_buf0), .Y(_1079_) );
OAI21X1 OAI21X1_257 ( .gnd(gnd), .vdd(vdd), .A(_1079_), .B(micro_hash_ucr_pipe15_bF_buf3), .C(_930__bF_buf1), .Y(_1080_) );
NAND2X1 NAND2X1_86 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_1_), .B(_1080_), .Y(_1081_) );
OAI21X1 OAI21X1_258 ( .gnd(gnd), .vdd(vdd), .A(_1078_), .B(micro_hash_ucr_pipe16_bF_buf1), .C(_1081_), .Y(_1082_) );
NAND2X1 NAND2X1_87 ( .gnd(gnd), .vdd(vdd), .A(_929_), .B(_1082_), .Y(_1083_) );
OAI21X1 OAI21X1_259 ( .gnd(gnd), .vdd(vdd), .A(_929_), .B(_1061_), .C(_1083_), .Y(_1084_) );
OAI21X1 OAI21X1_260 ( .gnd(gnd), .vdd(vdd), .A(_442_), .B(_925__bF_buf1), .C(_927__bF_buf1), .Y(_1085_) );
AOI21X1 AOI21X1_201 ( .gnd(gnd), .vdd(vdd), .A(_925__bF_buf0), .B(_1084_), .C(_1085_), .Y(_1086_) );
AOI21X1 AOI21X1_202 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe19_bF_buf0), .B(_1061_), .C(_1086_), .Y(_1087_) );
NAND2X1 NAND2X1_88 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe20_bF_buf2), .B(_442_), .Y(_1088_) );
OAI21X1 OAI21X1_261 ( .gnd(gnd), .vdd(vdd), .A(_1087_), .B(micro_hash_ucr_pipe20_bF_buf1), .C(_1088_), .Y(_1089_) );
NAND2X1 NAND2X1_89 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe21_bF_buf2), .B(_1060_), .Y(_1090_) );
OAI21X1 OAI21X1_262 ( .gnd(gnd), .vdd(vdd), .A(_1089_), .B(micro_hash_ucr_pipe21_bF_buf1), .C(_1090_), .Y(_1091_) );
NAND2X1 NAND2X1_90 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe22_bF_buf2), .B(_442_), .Y(_1092_) );
OAI21X1 OAI21X1_263 ( .gnd(gnd), .vdd(vdd), .A(_1091_), .B(micro_hash_ucr_pipe22_bF_buf1), .C(_1092_), .Y(_1093_) );
AOI21X1 AOI21X1_203 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe23_bF_buf0), .B(_1060_), .C(micro_hash_ucr_pipe24_bF_buf1), .Y(_1094_) );
OAI21X1 OAI21X1_264 ( .gnd(gnd), .vdd(vdd), .A(_1093_), .B(micro_hash_ucr_pipe23_bF_buf3), .C(_1094_), .Y(_1095_) );
AOI21X1 AOI21X1_204 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe24_bF_buf0), .B(_442_), .C(micro_hash_ucr_pipe25), .Y(_1096_) );
OAI21X1 OAI21X1_265 ( .gnd(gnd), .vdd(vdd), .A(_1061_), .B(_921__bF_buf3), .C(_920__bF_buf1), .Y(_1097_) );
AOI21X1 AOI21X1_205 ( .gnd(gnd), .vdd(vdd), .A(_1096_), .B(_1095_), .C(_1097_), .Y(_1098_) );
NOR2X1 NOR2X1_252 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_1_), .B(_920__bF_buf0), .Y(_1099_) );
OAI21X1 OAI21X1_266 ( .gnd(gnd), .vdd(vdd), .A(_1098_), .B(_1099_), .C(_916_), .Y(_1100_) );
OAI21X1 OAI21X1_267 ( .gnd(gnd), .vdd(vdd), .A(_1059_), .B(_1057_), .C(micro_hash_ucr_pipe27), .Y(_1101_) );
NAND3X1 NAND3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_918__bF_buf1), .B(_1101_), .C(_1100_), .Y(_1102_) );
AOI21X1 AOI21X1_206 ( .gnd(gnd), .vdd(vdd), .A(_1069_), .B(_1102_), .C(micro_hash_ucr_pipe29_bF_buf2), .Y(_1103_) );
OAI21X1 OAI21X1_268 ( .gnd(gnd), .vdd(vdd), .A(_1061_), .B(_917_), .C(_913__bF_buf2), .Y(_1104_) );
AOI21X1 AOI21X1_207 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe30_bF_buf1), .B(_442_), .C(micro_hash_ucr_pipe31), .Y(_1105_) );
OAI21X1 OAI21X1_269 ( .gnd(gnd), .vdd(vdd), .A(_1103_), .B(_1104_), .C(_1105_), .Y(_1106_) );
OAI21X1 OAI21X1_270 ( .gnd(gnd), .vdd(vdd), .A(_915__bF_buf1), .B(_1061_), .C(_1106_), .Y(_1107_) );
NAND2X1 NAND2X1_91 ( .gnd(gnd), .vdd(vdd), .A(_914__bF_buf1), .B(_1107_), .Y(_1108_) );
OAI21X1 OAI21X1_271 ( .gnd(gnd), .vdd(vdd), .A(_442_), .B(_914__bF_buf0), .C(_1108_), .Y(_1109_) );
OAI21X1 OAI21X1_272 ( .gnd(gnd), .vdd(vdd), .A(_1061_), .B(_910_), .C(_912__bF_buf3), .Y(_1110_) );
AOI21X1 AOI21X1_208 ( .gnd(gnd), .vdd(vdd), .A(_910_), .B(_1109_), .C(_1110_), .Y(_1111_) );
OAI21X1 OAI21X1_273 ( .gnd(gnd), .vdd(vdd), .A(_912__bF_buf2), .B(micro_hash_ucr_a_1_), .C(_911__bF_buf1), .Y(_1112_) );
AOI21X1 AOI21X1_209 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe35), .B(_1060_), .C(micro_hash_ucr_pipe36_bF_buf0), .Y(_1113_) );
OAI21X1 OAI21X1_274 ( .gnd(gnd), .vdd(vdd), .A(_1111_), .B(_1112_), .C(_1113_), .Y(_1114_) );
NAND2X1 NAND2X1_92 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe36_bF_buf3), .B(_442_), .Y(_1115_) );
AOI21X1 AOI21X1_210 ( .gnd(gnd), .vdd(vdd), .A(_1115_), .B(_1114_), .C(micro_hash_ucr_pipe37), .Y(_1116_) );
NOR2X1 NOR2X1_253 ( .gnd(gnd), .vdd(vdd), .A(_909__bF_buf1), .B(_1060_), .Y(_1117_) );
OAI21X1 OAI21X1_275 ( .gnd(gnd), .vdd(vdd), .A(_1116_), .B(_1117_), .C(_908__bF_buf1), .Y(_1118_) );
NAND3X1 NAND3X1_21 ( .gnd(gnd), .vdd(vdd), .A(_904__bF_buf0), .B(_1068_), .C(_1118_), .Y(_1119_) );
AOI21X1 AOI21X1_211 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe39), .B(_1060_), .C(micro_hash_ucr_pipe40_bF_buf3), .Y(_1120_) );
OAI21X1 OAI21X1_276 ( .gnd(gnd), .vdd(vdd), .A(_906__bF_buf1), .B(micro_hash_ucr_a_1_), .C(_905__bF_buf1), .Y(_1121_) );
AOI21X1 AOI21X1_212 ( .gnd(gnd), .vdd(vdd), .A(_1120_), .B(_1119_), .C(_1121_), .Y(_1122_) );
OAI21X1 OAI21X1_277 ( .gnd(gnd), .vdd(vdd), .A(_1061_), .B(_905__bF_buf0), .C(_901__bF_buf2), .Y(_1123_) );
OAI22X1 OAI22X1_21 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_1_), .B(_901__bF_buf1), .C(_1122_), .D(_1123_), .Y(_1124_) );
OAI21X1 OAI21X1_278 ( .gnd(gnd), .vdd(vdd), .A(_1060_), .B(_903__bF_buf0), .C(_902__bF_buf1), .Y(_1125_) );
AOI21X1 AOI21X1_213 ( .gnd(gnd), .vdd(vdd), .A(_903__bF_buf3), .B(_1124_), .C(_1125_), .Y(_1126_) );
NOR2X1 NOR2X1_254 ( .gnd(gnd), .vdd(vdd), .A(_442_), .B(_902__bF_buf0), .Y(_1127_) );
OAI21X1 OAI21X1_279 ( .gnd(gnd), .vdd(vdd), .A(_1126_), .B(_1127_), .C(_898_), .Y(_1128_) );
NAND2X1 NAND2X1_93 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe45_bF_buf2), .B(_1060_), .Y(_1129_) );
AOI21X1 AOI21X1_214 ( .gnd(gnd), .vdd(vdd), .A(_1129_), .B(_1128_), .C(micro_hash_ucr_pipe46_bF_buf3), .Y(_1130_) );
OAI21X1 OAI21X1_280 ( .gnd(gnd), .vdd(vdd), .A(_1130_), .B(_1067_), .C(_899__bF_buf0), .Y(_1131_) );
NAND2X1 NAND2X1_94 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe47), .B(_1060_), .Y(_1132_) );
AOI21X1 AOI21X1_215 ( .gnd(gnd), .vdd(vdd), .A(_1132_), .B(_1131_), .C(micro_hash_ucr_pipe48_bF_buf2), .Y(_1133_) );
OAI21X1 OAI21X1_281 ( .gnd(gnd), .vdd(vdd), .A(_442_), .B(_895__bF_buf1), .C(_897__bF_buf0), .Y(_1134_) );
AOI21X1 AOI21X1_216 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe49), .B(_1061_), .C(micro_hash_ucr_pipe50_bF_buf2), .Y(_1135_) );
OAI21X1 OAI21X1_282 ( .gnd(gnd), .vdd(vdd), .A(_1133_), .B(_1134_), .C(_1135_), .Y(_1136_) );
NAND2X1 NAND2X1_95 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_1_), .B(micro_hash_ucr_pipe50_bF_buf1), .Y(_1137_) );
AOI21X1 AOI21X1_217 ( .gnd(gnd), .vdd(vdd), .A(_1137_), .B(_1136_), .C(micro_hash_ucr_pipe51), .Y(_1138_) );
NOR2X1 NOR2X1_255 ( .gnd(gnd), .vdd(vdd), .A(_892_), .B(_1061_), .Y(_1139_) );
OAI21X1 OAI21X1_283 ( .gnd(gnd), .vdd(vdd), .A(_1138_), .B(_1139_), .C(_894__bF_buf0), .Y(_1140_) );
AOI21X1 AOI21X1_218 ( .gnd(gnd), .vdd(vdd), .A(_1066_), .B(_1140_), .C(micro_hash_ucr_pipe53_bF_buf2), .Y(_1141_) );
NOR2X1 NOR2X1_256 ( .gnd(gnd), .vdd(vdd), .A(_893_), .B(_1061_), .Y(_1142_) );
OAI21X1 OAI21X1_284 ( .gnd(gnd), .vdd(vdd), .A(_1141_), .B(_1142_), .C(_889__bF_buf1), .Y(_1143_) );
AOI21X1 AOI21X1_219 ( .gnd(gnd), .vdd(vdd), .A(_1065_), .B(_1143_), .C(micro_hash_ucr_pipe55), .Y(_1144_) );
NOR2X1 NOR2X1_257 ( .gnd(gnd), .vdd(vdd), .A(_891_), .B(_1061_), .Y(_1145_) );
OAI21X1 OAI21X1_285 ( .gnd(gnd), .vdd(vdd), .A(_1144_), .B(_1145_), .C(_890__bF_buf1), .Y(_1146_) );
AOI21X1 AOI21X1_220 ( .gnd(gnd), .vdd(vdd), .A(_1064_), .B(_1146_), .C(micro_hash_ucr_pipe57_bF_buf2), .Y(_1147_) );
NOR2X1 NOR2X1_258 ( .gnd(gnd), .vdd(vdd), .A(_886_), .B(_1061_), .Y(_1148_) );
OAI21X1 OAI21X1_286 ( .gnd(gnd), .vdd(vdd), .A(_1147_), .B(_1148_), .C(_888__bF_buf1), .Y(_1149_) );
AOI21X1 AOI21X1_221 ( .gnd(gnd), .vdd(vdd), .A(_1063_), .B(_1149_), .C(micro_hash_ucr_pipe59), .Y(_1150_) );
OAI21X1 OAI21X1_287 ( .gnd(gnd), .vdd(vdd), .A(_1061_), .B(_887__bF_buf1), .C(_883__bF_buf1), .Y(_1151_) );
AOI21X1 AOI21X1_222 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe60_bF_buf2), .B(_442_), .C(micro_hash_ucr_pipe61_bF_buf2), .Y(_1152_) );
OAI21X1 OAI21X1_288 ( .gnd(gnd), .vdd(vdd), .A(_1150_), .B(_1151_), .C(_1152_), .Y(_1153_) );
NAND2X1 NAND2X1_96 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe61_bF_buf1), .B(_1060_), .Y(_1154_) );
AOI21X1 AOI21X1_223 ( .gnd(gnd), .vdd(vdd), .A(_1154_), .B(_1153_), .C(micro_hash_ucr_pipe62_bF_buf3), .Y(_1155_) );
OAI21X1 OAI21X1_289 ( .gnd(gnd), .vdd(vdd), .A(_1155_), .B(_1062_), .C(_880__bF_buf0), .Y(_1156_) );
OAI21X1 OAI21X1_290 ( .gnd(gnd), .vdd(vdd), .A(_880__bF_buf3), .B(_1061_), .C(_1156_), .Y(_1157_) );
NAND2X1 NAND2X1_97 ( .gnd(gnd), .vdd(vdd), .A(_882__bF_buf0), .B(_1157_), .Y(_1158_) );
OAI21X1 OAI21X1_291 ( .gnd(gnd), .vdd(vdd), .A(_442_), .B(_882__bF_buf3), .C(_1158_), .Y(_1159_) );
OAI21X1 OAI21X1_292 ( .gnd(gnd), .vdd(vdd), .A(_1059_), .B(_1057_), .C(micro_hash_ucr_pipe65_bF_buf1), .Y(_1160_) );
OAI21X1 OAI21X1_293 ( .gnd(gnd), .vdd(vdd), .A(_1159_), .B(micro_hash_ucr_pipe65_bF_buf0), .C(_1160_), .Y(_1161_) );
OAI21X1 OAI21X1_294 ( .gnd(gnd), .vdd(vdd), .A(_877__bF_buf1), .B(micro_hash_ucr_a_1_), .C(_879__bF_buf0), .Y(_1162_) );
AOI21X1 AOI21X1_224 ( .gnd(gnd), .vdd(vdd), .A(_877__bF_buf0), .B(_1161_), .C(_1162_), .Y(_1163_) );
OAI21X1 OAI21X1_295 ( .gnd(gnd), .vdd(vdd), .A(_1061_), .B(_879__bF_buf3), .C(_878__bF_buf1), .Y(_1164_) );
OAI22X1 OAI22X1_22 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_1_), .B(_878__bF_buf0), .C(_1163_), .D(_1164_), .Y(_1165_) );
OAI21X1 OAI21X1_296 ( .gnd(gnd), .vdd(vdd), .A(_1060_), .B(_876__bF_buf0), .C(_302__bF_buf13), .Y(_1166_) );
AOI21X1 AOI21X1_225 ( .gnd(gnd), .vdd(vdd), .A(_876__bF_buf3), .B(_1165_), .C(_1166_), .Y(_297__1_) );
INVX8 INVX8_77 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_2_), .Y(_1167_) );
NAND2X1 NAND2X1_98 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_2_), .B(micro_hash_ucr_pipe62_bF_buf2), .Y(_1168_) );
NAND2X1 NAND2X1_99 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_2_), .B(micro_hash_ucr_pipe60_bF_buf1), .Y(_1169_) );
NAND2X1 NAND2X1_100 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe54_bF_buf1), .B(_1167__bF_buf3), .Y(_1170_) );
NAND2X1 NAND2X1_101 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe52_bF_buf2), .B(_1167__bF_buf2), .Y(_1171_) );
NAND2X1 NAND2X1_102 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe50_bF_buf0), .B(_1167__bF_buf1), .Y(_1172_) );
NAND2X1 NAND2X1_103 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe48_bF_buf1), .B(_1167__bF_buf0), .Y(_1173_) );
INVX8 INVX8_78 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_2_bF_buf1_), .Y(_1174_) );
NAND2X1 NAND2X1_104 ( .gnd(gnd), .vdd(vdd), .A(_1174_), .B(_389_), .Y(_1175_) );
NAND2X1 NAND2X1_105 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_2_bF_buf0_), .B(micro_hash_ucr_b_2_bF_buf1_), .Y(_1176_) );
NAND2X1 NAND2X1_106 ( .gnd(gnd), .vdd(vdd), .A(_1176_), .B(_1175_), .Y(_1177_) );
INVX8 INVX8_79 ( .gnd(gnd), .vdd(vdd), .A(_1177_), .Y(_1178_) );
NOR2X1 NOR2X1_259 ( .gnd(gnd), .vdd(vdd), .A(_1167__bF_buf3), .B(_918__bF_buf0), .Y(_1179_) );
NOR2X1 NOR2X1_260 ( .gnd(gnd), .vdd(vdd), .A(_1167__bF_buf2), .B(_920__bF_buf4), .Y(_1180_) );
NOR2X1 NOR2X1_261 ( .gnd(gnd), .vdd(vdd), .A(_1167__bF_buf1), .B(_919__bF_buf2), .Y(_1181_) );
NOR2X1 NOR2X1_262 ( .gnd(gnd), .vdd(vdd), .A(_1167__bF_buf0), .B(_924__bF_buf1), .Y(_1182_) );
NAND2X1 NAND2X1_107 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe17_bF_buf1), .B(_1178__bF_buf3), .Y(_1183_) );
NAND2X1 NAND2X1_108 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe15_bF_buf2), .B(_1178__bF_buf2), .Y(_1184_) );
NAND2X1 NAND2X1_109 ( .gnd(gnd), .vdd(vdd), .A(_1167__bF_buf3), .B(_957_), .Y(_1185_) );
OR2X2 OR2X2_26 ( .gnd(gnd), .vdd(vdd), .A(_955_), .B(_1072_), .Y(_1186_) );
NOR2X1 NOR2X1_263 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe12), .B(micro_hash_ucr_pipe10), .Y(_1187_) );
NOR2X1 NOR2X1_264 ( .gnd(gnd), .vdd(vdd), .A(H_2_), .B(micro_hash_ucr_pipe7), .Y(_1188_) );
NAND2X1 NAND2X1_110 ( .gnd(gnd), .vdd(vdd), .A(_1187_), .B(_1188_), .Y(_1189_) );
OAI21X1 OAI21X1_297 ( .gnd(gnd), .vdd(vdd), .A(_1186_), .B(_1189_), .C(_1185_), .Y(_1190_) );
NAND2X1 NAND2X1_111 ( .gnd(gnd), .vdd(vdd), .A(_933_), .B(_1190_), .Y(_1191_) );
NOR2X1 NOR2X1_265 ( .gnd(gnd), .vdd(vdd), .A(_1178__bF_buf1), .B(_1070_), .Y(_1192_) );
NOR2X1 NOR2X1_266 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe14_bF_buf4), .B(_1192_), .Y(_1193_) );
AOI22X1 AOI22X1_14 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_2_), .B(micro_hash_ucr_pipe14_bF_buf3), .C(_1193_), .D(_1191_), .Y(_1194_) );
OAI21X1 OAI21X1_298 ( .gnd(gnd), .vdd(vdd), .A(_1194_), .B(micro_hash_ucr_pipe15_bF_buf1), .C(_1184_), .Y(_1195_) );
NAND2X1 NAND2X1_112 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe16_bF_buf0), .B(_1167__bF_buf2), .Y(_1196_) );
OAI21X1 OAI21X1_299 ( .gnd(gnd), .vdd(vdd), .A(_1195_), .B(micro_hash_ucr_pipe16_bF_buf3), .C(_1196_), .Y(_1197_) );
OAI21X1 OAI21X1_300 ( .gnd(gnd), .vdd(vdd), .A(_1197_), .B(micro_hash_ucr_pipe17_bF_buf0), .C(_1183_), .Y(_1198_) );
OAI21X1 OAI21X1_301 ( .gnd(gnd), .vdd(vdd), .A(_1167__bF_buf1), .B(_925__bF_buf4), .C(_927__bF_buf0), .Y(_1199_) );
AOI21X1 AOI21X1_226 ( .gnd(gnd), .vdd(vdd), .A(_925__bF_buf3), .B(_1198_), .C(_1199_), .Y(_1200_) );
OAI21X1 OAI21X1_302 ( .gnd(gnd), .vdd(vdd), .A(_1178__bF_buf0), .B(_927__bF_buf3), .C(_926__bF_buf1), .Y(_1201_) );
OAI22X1 OAI22X1_23 ( .gnd(gnd), .vdd(vdd), .A(_1167__bF_buf0), .B(_926__bF_buf0), .C(_1200_), .D(_1201_), .Y(_1202_) );
NAND2X1 NAND2X1_113 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe21_bF_buf0), .B(_1177_), .Y(_1203_) );
OAI21X1 OAI21X1_303 ( .gnd(gnd), .vdd(vdd), .A(_1202_), .B(micro_hash_ucr_pipe21_bF_buf3), .C(_1203_), .Y(_1204_) );
NOR2X1 NOR2X1_267 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe22_bF_buf0), .B(_1204_), .Y(_1205_) );
OAI21X1 OAI21X1_304 ( .gnd(gnd), .vdd(vdd), .A(_1205_), .B(_1182_), .C(_923_), .Y(_1206_) );
NAND2X1 NAND2X1_114 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe23_bF_buf2), .B(_1178__bF_buf3), .Y(_1207_) );
AOI21X1 AOI21X1_227 ( .gnd(gnd), .vdd(vdd), .A(_1207_), .B(_1206_), .C(micro_hash_ucr_pipe24_bF_buf4), .Y(_1208_) );
OAI21X1 OAI21X1_305 ( .gnd(gnd), .vdd(vdd), .A(_1208_), .B(_1181_), .C(_921__bF_buf2), .Y(_1209_) );
NAND2X1 NAND2X1_115 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe25), .B(_1178__bF_buf2), .Y(_1210_) );
AOI21X1 AOI21X1_228 ( .gnd(gnd), .vdd(vdd), .A(_1210_), .B(_1209_), .C(micro_hash_ucr_pipe26_bF_buf1), .Y(_1211_) );
OAI21X1 OAI21X1_306 ( .gnd(gnd), .vdd(vdd), .A(_1211_), .B(_1180_), .C(_916_), .Y(_1212_) );
NAND2X1 NAND2X1_116 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe27), .B(_1178__bF_buf1), .Y(_1213_) );
AOI21X1 AOI21X1_229 ( .gnd(gnd), .vdd(vdd), .A(_1213_), .B(_1212_), .C(micro_hash_ucr_pipe28_bF_buf1), .Y(_1214_) );
OAI21X1 OAI21X1_307 ( .gnd(gnd), .vdd(vdd), .A(_1214_), .B(_1179_), .C(_917_), .Y(_1215_) );
AOI21X1 AOI21X1_230 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe29_bF_buf1), .B(_1178__bF_buf0), .C(micro_hash_ucr_pipe30_bF_buf0), .Y(_1216_) );
OAI21X1 OAI21X1_308 ( .gnd(gnd), .vdd(vdd), .A(_913__bF_buf1), .B(micro_hash_ucr_a_2_), .C(_915__bF_buf0), .Y(_1217_) );
AOI21X1 AOI21X1_231 ( .gnd(gnd), .vdd(vdd), .A(_1216_), .B(_1215_), .C(_1217_), .Y(_1218_) );
OAI21X1 OAI21X1_309 ( .gnd(gnd), .vdd(vdd), .A(_1177_), .B(_915__bF_buf3), .C(_914__bF_buf4), .Y(_1219_) );
OAI22X1 OAI22X1_24 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_2_), .B(_914__bF_buf3), .C(_1218_), .D(_1219_), .Y(_1220_) );
AOI21X1 AOI21X1_232 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe33_bF_buf2), .B(_1178__bF_buf3), .C(micro_hash_ucr_pipe34_bF_buf0), .Y(_1221_) );
OAI21X1 OAI21X1_310 ( .gnd(gnd), .vdd(vdd), .A(_1220_), .B(micro_hash_ucr_pipe33_bF_buf1), .C(_1221_), .Y(_1222_) );
AOI21X1 AOI21X1_233 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe34_bF_buf3), .B(_1167__bF_buf3), .C(micro_hash_ucr_pipe35), .Y(_1223_) );
OAI21X1 OAI21X1_311 ( .gnd(gnd), .vdd(vdd), .A(_1177_), .B(_911__bF_buf0), .C(_907__bF_buf3), .Y(_1224_) );
AOI21X1 AOI21X1_234 ( .gnd(gnd), .vdd(vdd), .A(_1223_), .B(_1222_), .C(_1224_), .Y(_1225_) );
NOR2X1 NOR2X1_268 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_2_), .B(_907__bF_buf2), .Y(_1226_) );
OAI21X1 OAI21X1_312 ( .gnd(gnd), .vdd(vdd), .A(_1225_), .B(_1226_), .C(_909__bF_buf0), .Y(_1227_) );
OAI21X1 OAI21X1_313 ( .gnd(gnd), .vdd(vdd), .A(_909__bF_buf3), .B(_1178__bF_buf2), .C(_1227_), .Y(_1228_) );
NAND2X1 NAND2X1_117 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_2_), .B(micro_hash_ucr_pipe38_bF_buf1), .Y(_1229_) );
OAI21X1 OAI21X1_314 ( .gnd(gnd), .vdd(vdd), .A(_1228_), .B(micro_hash_ucr_pipe38_bF_buf0), .C(_1229_), .Y(_1230_) );
NAND2X1 NAND2X1_118 ( .gnd(gnd), .vdd(vdd), .A(_904__bF_buf3), .B(_1230_), .Y(_1231_) );
OAI21X1 OAI21X1_315 ( .gnd(gnd), .vdd(vdd), .A(_904__bF_buf2), .B(_1177_), .C(_1231_), .Y(_1232_) );
AOI21X1 AOI21X1_235 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe40_bF_buf2), .B(_1167__bF_buf2), .C(micro_hash_ucr_pipe41), .Y(_1233_) );
OAI21X1 OAI21X1_316 ( .gnd(gnd), .vdd(vdd), .A(_1232_), .B(micro_hash_ucr_pipe40_bF_buf1), .C(_1233_), .Y(_1234_) );
OAI21X1 OAI21X1_317 ( .gnd(gnd), .vdd(vdd), .A(_905__bF_buf3), .B(_1177_), .C(_1234_), .Y(_1235_) );
NAND2X1 NAND2X1_119 ( .gnd(gnd), .vdd(vdd), .A(_901__bF_buf0), .B(_1235_), .Y(_1236_) );
OAI21X1 OAI21X1_318 ( .gnd(gnd), .vdd(vdd), .A(_1167__bF_buf1), .B(_901__bF_buf4), .C(_1236_), .Y(_1237_) );
OAI21X1 OAI21X1_319 ( .gnd(gnd), .vdd(vdd), .A(_1177_), .B(_903__bF_buf2), .C(_902__bF_buf4), .Y(_1238_) );
AOI21X1 AOI21X1_236 ( .gnd(gnd), .vdd(vdd), .A(_903__bF_buf1), .B(_1237_), .C(_1238_), .Y(_1239_) );
OAI21X1 OAI21X1_320 ( .gnd(gnd), .vdd(vdd), .A(_902__bF_buf3), .B(micro_hash_ucr_a_2_), .C(_898_), .Y(_1240_) );
AOI21X1 AOI21X1_237 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe45_bF_buf1), .B(_1178__bF_buf1), .C(micro_hash_ucr_pipe46_bF_buf2), .Y(_1241_) );
OAI21X1 OAI21X1_321 ( .gnd(gnd), .vdd(vdd), .A(_1239_), .B(_1240_), .C(_1241_), .Y(_1242_) );
NAND2X1 NAND2X1_120 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe46_bF_buf1), .B(_1167__bF_buf0), .Y(_1243_) );
AOI21X1 AOI21X1_238 ( .gnd(gnd), .vdd(vdd), .A(_1243_), .B(_1242_), .C(micro_hash_ucr_pipe47), .Y(_1244_) );
NOR2X1 NOR2X1_269 ( .gnd(gnd), .vdd(vdd), .A(_899__bF_buf3), .B(_1178__bF_buf0), .Y(_1245_) );
OAI21X1 OAI21X1_322 ( .gnd(gnd), .vdd(vdd), .A(_1244_), .B(_1245_), .C(_895__bF_buf0), .Y(_1246_) );
NAND3X1 NAND3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_897__bF_buf3), .B(_1173_), .C(_1246_), .Y(_1247_) );
NAND2X1 NAND2X1_121 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe49), .B(_1178__bF_buf3), .Y(_1248_) );
NAND3X1 NAND3X1_23 ( .gnd(gnd), .vdd(vdd), .A(_896__bF_buf1), .B(_1248_), .C(_1247_), .Y(_1249_) );
NAND3X1 NAND3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_892_), .B(_1172_), .C(_1249_), .Y(_1250_) );
NAND2X1 NAND2X1_122 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe51), .B(_1178__bF_buf2), .Y(_1251_) );
NAND3X1 NAND3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_894__bF_buf3), .B(_1251_), .C(_1250_), .Y(_1252_) );
NAND3X1 NAND3X1_26 ( .gnd(gnd), .vdd(vdd), .A(_893_), .B(_1171_), .C(_1252_), .Y(_1253_) );
NAND2X1 NAND2X1_123 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe53_bF_buf1), .B(_1178__bF_buf1), .Y(_1254_) );
NAND3X1 NAND3X1_27 ( .gnd(gnd), .vdd(vdd), .A(_889__bF_buf0), .B(_1254_), .C(_1253_), .Y(_1255_) );
NAND3X1 NAND3X1_28 ( .gnd(gnd), .vdd(vdd), .A(_891_), .B(_1170_), .C(_1255_), .Y(_1256_) );
NAND2X1 NAND2X1_124 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe55), .B(_1178__bF_buf0), .Y(_1257_) );
AOI21X1 AOI21X1_239 ( .gnd(gnd), .vdd(vdd), .A(_1257_), .B(_1256_), .C(micro_hash_ucr_pipe56_bF_buf1), .Y(_1258_) );
OAI21X1 OAI21X1_323 ( .gnd(gnd), .vdd(vdd), .A(_1167__bF_buf3), .B(_890__bF_buf0), .C(_886_), .Y(_1259_) );
AOI21X1 AOI21X1_240 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe57_bF_buf1), .B(_1177_), .C(micro_hash_ucr_pipe58_bF_buf1), .Y(_1260_) );
OAI21X1 OAI21X1_324 ( .gnd(gnd), .vdd(vdd), .A(_1258_), .B(_1259_), .C(_1260_), .Y(_1261_) );
NAND2X1 NAND2X1_125 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_2_), .B(micro_hash_ucr_pipe58_bF_buf0), .Y(_1262_) );
NAND3X1 NAND3X1_29 ( .gnd(gnd), .vdd(vdd), .A(_887__bF_buf0), .B(_1262_), .C(_1261_), .Y(_1263_) );
NAND2X1 NAND2X1_126 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe59), .B(_1177_), .Y(_1264_) );
NAND3X1 NAND3X1_30 ( .gnd(gnd), .vdd(vdd), .A(_883__bF_buf0), .B(_1264_), .C(_1263_), .Y(_1265_) );
NAND3X1 NAND3X1_31 ( .gnd(gnd), .vdd(vdd), .A(_885_), .B(_1169_), .C(_1265_), .Y(_1266_) );
NAND2X1 NAND2X1_127 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe61_bF_buf0), .B(_1177_), .Y(_1267_) );
NAND3X1 NAND3X1_32 ( .gnd(gnd), .vdd(vdd), .A(_884__bF_buf0), .B(_1267_), .C(_1266_), .Y(_1268_) );
AOI21X1 AOI21X1_241 ( .gnd(gnd), .vdd(vdd), .A(_1168_), .B(_1268_), .C(micro_hash_ucr_pipe63), .Y(_1269_) );
OAI21X1 OAI21X1_325 ( .gnd(gnd), .vdd(vdd), .A(_1177_), .B(_880__bF_buf2), .C(_882__bF_buf2), .Y(_1270_) );
AOI21X1 AOI21X1_242 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe64_bF_buf3), .B(_1167__bF_buf2), .C(micro_hash_ucr_pipe65_bF_buf3), .Y(_1271_) );
OAI21X1 OAI21X1_326 ( .gnd(gnd), .vdd(vdd), .A(_1269_), .B(_1270_), .C(_1271_), .Y(_1272_) );
AOI21X1 AOI21X1_243 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe65_bF_buf2), .B(_1178__bF_buf3), .C(micro_hash_ucr_pipe66_bF_buf2), .Y(_1273_) );
AOI22X1 AOI22X1_15 ( .gnd(gnd), .vdd(vdd), .A(_1167__bF_buf1), .B(micro_hash_ucr_pipe66_bF_buf1), .C(_1272_), .D(_1273_), .Y(_1274_) );
AOI21X1 AOI21X1_244 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe67), .B(_1177_), .C(micro_hash_ucr_pipe68), .Y(_1275_) );
OAI21X1 OAI21X1_327 ( .gnd(gnd), .vdd(vdd), .A(_1274_), .B(micro_hash_ucr_pipe67), .C(_1275_), .Y(_1276_) );
AOI21X1 AOI21X1_245 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_2_), .B(micro_hash_ucr_pipe68), .C(micro_hash_ucr_pipe69), .Y(_1277_) );
OAI21X1 OAI21X1_328 ( .gnd(gnd), .vdd(vdd), .A(_1178__bF_buf2), .B(_876__bF_buf2), .C(_302__bF_buf12), .Y(_1278_) );
AOI21X1 AOI21X1_246 ( .gnd(gnd), .vdd(vdd), .A(_1277_), .B(_1276_), .C(_1278_), .Y(_297__2_) );
NOR2X1 NOR2X1_270 ( .gnd(gnd), .vdd(vdd), .A(_460__bF_buf2), .B(_882__bF_buf1), .Y(_1279_) );
NOR2X1 NOR2X1_271 ( .gnd(gnd), .vdd(vdd), .A(_460__bF_buf1), .B(_884__bF_buf4), .Y(_1280_) );
NAND2X1 NAND2X1_128 ( .gnd(gnd), .vdd(vdd), .A(_4445_), .B(_394_), .Y(_1281_) );
NAND2X1 NAND2X1_129 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_3_bF_buf2_), .B(micro_hash_ucr_b_3_bF_buf1_), .Y(_1282_) );
NAND2X1 NAND2X1_130 ( .gnd(gnd), .vdd(vdd), .A(_1282_), .B(_1281_), .Y(_1283_) );
NOR2X1 NOR2X1_272 ( .gnd(gnd), .vdd(vdd), .A(_460__bF_buf0), .B(_889__bF_buf4), .Y(_1284_) );
NOR2X1 NOR2X1_273 ( .gnd(gnd), .vdd(vdd), .A(_460__bF_buf3), .B(_894__bF_buf2), .Y(_1285_) );
NOR2X1 NOR2X1_274 ( .gnd(gnd), .vdd(vdd), .A(_460__bF_buf2), .B(_896__bF_buf0), .Y(_1286_) );
NOR2X1 NOR2X1_275 ( .gnd(gnd), .vdd(vdd), .A(_460__bF_buf1), .B(_895__bF_buf4), .Y(_1287_) );
NOR2X1 NOR2X1_276 ( .gnd(gnd), .vdd(vdd), .A(_460__bF_buf0), .B(_900__bF_buf3), .Y(_1288_) );
NOR2X1 NOR2X1_277 ( .gnd(gnd), .vdd(vdd), .A(_460__bF_buf3), .B(_902__bF_buf2), .Y(_1289_) );
INVX8 INVX8_80 ( .gnd(gnd), .vdd(vdd), .A(_1283_), .Y(_1290_) );
NOR2X1 NOR2X1_278 ( .gnd(gnd), .vdd(vdd), .A(_460__bF_buf2), .B(_920__bF_buf3), .Y(_1291_) );
NAND2X1 NAND2X1_131 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_3_), .B(micro_hash_ucr_pipe16_bF_buf2), .Y(_1292_) );
OR2X2 OR2X2_27 ( .gnd(gnd), .vdd(vdd), .A(_1079_), .B(micro_hash_ucr_a_3_), .Y(_1293_) );
NOR2X1 NOR2X1_279 ( .gnd(gnd), .vdd(vdd), .A(H_3_), .B(micro_hash_ucr_pipe9), .Y(_1294_) );
NAND2X1 NAND2X1_132 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe6), .B(_938_), .Y(_1295_) );
NOR2X1 NOR2X1_280 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe13), .B(micro_hash_ucr_pipe11), .Y(_1296_) );
NAND2X1 NAND2X1_133 ( .gnd(gnd), .vdd(vdd), .A(_1187_), .B(_1296_), .Y(_1297_) );
NOR2X1 NOR2X1_281 ( .gnd(gnd), .vdd(vdd), .A(_1295_), .B(_1297_), .Y(_1298_) );
NAND3X1 NAND3X1_33 ( .gnd(gnd), .vdd(vdd), .A(_939_), .B(_1294_), .C(_1298_), .Y(_1299_) );
OAI21X1 OAI21X1_329 ( .gnd(gnd), .vdd(vdd), .A(_1070_), .B(_1290__bF_buf3), .C(_1299_), .Y(_1300_) );
AOI21X1 AOI21X1_247 ( .gnd(gnd), .vdd(vdd), .A(_932_), .B(_1300_), .C(micro_hash_ucr_pipe15_bF_buf0), .Y(_1301_) );
AOI22X1 AOI22X1_16 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe15_bF_buf3), .B(_1290__bF_buf2), .C(_1301_), .D(_1293_), .Y(_1302_) );
OAI21X1 OAI21X1_330 ( .gnd(gnd), .vdd(vdd), .A(_1302_), .B(micro_hash_ucr_pipe16_bF_buf1), .C(_1292_), .Y(_1303_) );
NAND2X1 NAND2X1_134 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe17_bF_buf3), .B(_1283_), .Y(_1304_) );
OAI21X1 OAI21X1_331 ( .gnd(gnd), .vdd(vdd), .A(_1303_), .B(micro_hash_ucr_pipe17_bF_buf2), .C(_1304_), .Y(_1305_) );
NOR2X1 NOR2X1_282 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe18_bF_buf2), .B(_1305_), .Y(_1306_) );
OAI21X1 OAI21X1_332 ( .gnd(gnd), .vdd(vdd), .A(_460__bF_buf1), .B(_925__bF_buf2), .C(_927__bF_buf2), .Y(_1307_) );
AOI21X1 AOI21X1_248 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe19_bF_buf3), .B(_1283_), .C(micro_hash_ucr_pipe20_bF_buf0), .Y(_1308_) );
OAI21X1 OAI21X1_333 ( .gnd(gnd), .vdd(vdd), .A(_1306_), .B(_1307_), .C(_1308_), .Y(_1309_) );
OAI21X1 OAI21X1_334 ( .gnd(gnd), .vdd(vdd), .A(_460__bF_buf0), .B(_926__bF_buf4), .C(_1309_), .Y(_1310_) );
AND2X2 AND2X2_186 ( .gnd(gnd), .vdd(vdd), .A(_1310_), .B(_922_), .Y(_1311_) );
NOR2X1 NOR2X1_283 ( .gnd(gnd), .vdd(vdd), .A(_922_), .B(_1283_), .Y(_1312_) );
OAI21X1 OAI21X1_335 ( .gnd(gnd), .vdd(vdd), .A(_1311_), .B(_1312_), .C(_924__bF_buf0), .Y(_1313_) );
AOI21X1 AOI21X1_249 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_3_), .B(micro_hash_ucr_pipe22_bF_buf4), .C(micro_hash_ucr_pipe23_bF_buf1), .Y(_1314_) );
OAI21X1 OAI21X1_336 ( .gnd(gnd), .vdd(vdd), .A(_1290__bF_buf1), .B(_923_), .C(_919__bF_buf1), .Y(_1315_) );
AOI21X1 AOI21X1_250 ( .gnd(gnd), .vdd(vdd), .A(_1314_), .B(_1313_), .C(_1315_), .Y(_1316_) );
NOR2X1 NOR2X1_284 ( .gnd(gnd), .vdd(vdd), .A(_460__bF_buf3), .B(_919__bF_buf0), .Y(_1317_) );
OAI21X1 OAI21X1_337 ( .gnd(gnd), .vdd(vdd), .A(_1316_), .B(_1317_), .C(_921__bF_buf1), .Y(_1318_) );
NAND2X1 NAND2X1_135 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe25), .B(_1290__bF_buf0), .Y(_1319_) );
AOI21X1 AOI21X1_251 ( .gnd(gnd), .vdd(vdd), .A(_1319_), .B(_1318_), .C(micro_hash_ucr_pipe26_bF_buf0), .Y(_1320_) );
OAI21X1 OAI21X1_338 ( .gnd(gnd), .vdd(vdd), .A(_1320_), .B(_1291_), .C(_916_), .Y(_1321_) );
NAND2X1 NAND2X1_136 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe27), .B(_1290__bF_buf3), .Y(_1322_) );
AOI21X1 AOI21X1_252 ( .gnd(gnd), .vdd(vdd), .A(_1322_), .B(_1321_), .C(micro_hash_ucr_pipe28_bF_buf0), .Y(_1323_) );
OAI21X1 OAI21X1_339 ( .gnd(gnd), .vdd(vdd), .A(_460__bF_buf2), .B(_918__bF_buf4), .C(_917_), .Y(_1324_) );
OAI22X1 OAI22X1_25 ( .gnd(gnd), .vdd(vdd), .A(_917_), .B(_1290__bF_buf2), .C(_1323_), .D(_1324_), .Y(_1325_) );
OAI21X1 OAI21X1_340 ( .gnd(gnd), .vdd(vdd), .A(_913__bF_buf0), .B(micro_hash_ucr_a_3_), .C(_915__bF_buf2), .Y(_1326_) );
AOI21X1 AOI21X1_253 ( .gnd(gnd), .vdd(vdd), .A(_913__bF_buf4), .B(_1325_), .C(_1326_), .Y(_1327_) );
OAI21X1 OAI21X1_341 ( .gnd(gnd), .vdd(vdd), .A(_1283_), .B(_915__bF_buf1), .C(_914__bF_buf2), .Y(_1328_) );
OAI22X1 OAI22X1_26 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_3_), .B(_914__bF_buf1), .C(_1327_), .D(_1328_), .Y(_1329_) );
NAND2X1 NAND2X1_137 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe33_bF_buf0), .B(_1290__bF_buf1), .Y(_1330_) );
OAI21X1 OAI21X1_342 ( .gnd(gnd), .vdd(vdd), .A(_1329_), .B(micro_hash_ucr_pipe33_bF_buf3), .C(_1330_), .Y(_1331_) );
OAI21X1 OAI21X1_343 ( .gnd(gnd), .vdd(vdd), .A(_460__bF_buf1), .B(_912__bF_buf1), .C(_911__bF_buf4), .Y(_1332_) );
AOI21X1 AOI21X1_254 ( .gnd(gnd), .vdd(vdd), .A(_912__bF_buf0), .B(_1331_), .C(_1332_), .Y(_1333_) );
NOR2X1 NOR2X1_285 ( .gnd(gnd), .vdd(vdd), .A(_911__bF_buf3), .B(_1290__bF_buf0), .Y(_1334_) );
OAI21X1 OAI21X1_344 ( .gnd(gnd), .vdd(vdd), .A(_1333_), .B(_1334_), .C(_907__bF_buf1), .Y(_1335_) );
AOI21X1 AOI21X1_255 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe36_bF_buf2), .B(_460__bF_buf0), .C(micro_hash_ucr_pipe37), .Y(_1336_) );
OAI21X1 OAI21X1_345 ( .gnd(gnd), .vdd(vdd), .A(_1283_), .B(_909__bF_buf2), .C(_908__bF_buf0), .Y(_1337_) );
AOI21X1 AOI21X1_256 ( .gnd(gnd), .vdd(vdd), .A(_1336_), .B(_1335_), .C(_1337_), .Y(_1338_) );
NOR2X1 NOR2X1_286 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_3_), .B(_908__bF_buf4), .Y(_1339_) );
OAI21X1 OAI21X1_346 ( .gnd(gnd), .vdd(vdd), .A(_1338_), .B(_1339_), .C(_904__bF_buf1), .Y(_1340_) );
NAND2X1 NAND2X1_138 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe39), .B(_1283_), .Y(_1341_) );
NAND3X1 NAND3X1_34 ( .gnd(gnd), .vdd(vdd), .A(_906__bF_buf0), .B(_1341_), .C(_1340_), .Y(_1342_) );
AOI21X1 AOI21X1_257 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_3_), .B(micro_hash_ucr_pipe40_bF_buf0), .C(micro_hash_ucr_pipe41), .Y(_1343_) );
OAI21X1 OAI21X1_347 ( .gnd(gnd), .vdd(vdd), .A(_1290__bF_buf3), .B(_905__bF_buf2), .C(_901__bF_buf3), .Y(_1344_) );
AOI21X1 AOI21X1_258 ( .gnd(gnd), .vdd(vdd), .A(_1343_), .B(_1342_), .C(_1344_), .Y(_1345_) );
NOR2X1 NOR2X1_287 ( .gnd(gnd), .vdd(vdd), .A(_460__bF_buf3), .B(_901__bF_buf2), .Y(_1346_) );
OAI21X1 OAI21X1_348 ( .gnd(gnd), .vdd(vdd), .A(_1345_), .B(_1346_), .C(_903__bF_buf0), .Y(_1347_) );
NAND2X1 NAND2X1_139 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe43), .B(_1290__bF_buf2), .Y(_1348_) );
AOI21X1 AOI21X1_259 ( .gnd(gnd), .vdd(vdd), .A(_1348_), .B(_1347_), .C(micro_hash_ucr_pipe44), .Y(_1349_) );
OAI21X1 OAI21X1_349 ( .gnd(gnd), .vdd(vdd), .A(_1349_), .B(_1289_), .C(_898_), .Y(_1350_) );
NAND2X1 NAND2X1_140 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe45_bF_buf0), .B(_1290__bF_buf1), .Y(_1351_) );
AOI21X1 AOI21X1_260 ( .gnd(gnd), .vdd(vdd), .A(_1351_), .B(_1350_), .C(micro_hash_ucr_pipe46_bF_buf0), .Y(_1352_) );
OAI21X1 OAI21X1_350 ( .gnd(gnd), .vdd(vdd), .A(_1352_), .B(_1288_), .C(_899__bF_buf2), .Y(_1353_) );
NAND2X1 NAND2X1_141 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe47), .B(_1290__bF_buf0), .Y(_1354_) );
AOI21X1 AOI21X1_261 ( .gnd(gnd), .vdd(vdd), .A(_1354_), .B(_1353_), .C(micro_hash_ucr_pipe48_bF_buf0), .Y(_1355_) );
OAI21X1 OAI21X1_351 ( .gnd(gnd), .vdd(vdd), .A(_1355_), .B(_1287_), .C(_897__bF_buf2), .Y(_1356_) );
NAND2X1 NAND2X1_142 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe49), .B(_1290__bF_buf3), .Y(_1357_) );
AOI21X1 AOI21X1_262 ( .gnd(gnd), .vdd(vdd), .A(_1357_), .B(_1356_), .C(micro_hash_ucr_pipe50_bF_buf3), .Y(_1358_) );
OAI21X1 OAI21X1_352 ( .gnd(gnd), .vdd(vdd), .A(_1358_), .B(_1286_), .C(_892_), .Y(_1359_) );
NAND2X1 NAND2X1_143 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe51), .B(_1290__bF_buf2), .Y(_1360_) );
AOI21X1 AOI21X1_263 ( .gnd(gnd), .vdd(vdd), .A(_1360_), .B(_1359_), .C(micro_hash_ucr_pipe52_bF_buf1), .Y(_1361_) );
OAI21X1 OAI21X1_353 ( .gnd(gnd), .vdd(vdd), .A(_1361_), .B(_1285_), .C(_893_), .Y(_1362_) );
NAND2X1 NAND2X1_144 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe53_bF_buf0), .B(_1290__bF_buf1), .Y(_1363_) );
AOI21X1 AOI21X1_264 ( .gnd(gnd), .vdd(vdd), .A(_1363_), .B(_1362_), .C(micro_hash_ucr_pipe54_bF_buf0), .Y(_1364_) );
OAI21X1 OAI21X1_354 ( .gnd(gnd), .vdd(vdd), .A(_1364_), .B(_1284_), .C(_891_), .Y(_1365_) );
NAND2X1 NAND2X1_145 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe55), .B(_1290__bF_buf0), .Y(_1366_) );
AOI21X1 AOI21X1_265 ( .gnd(gnd), .vdd(vdd), .A(_1366_), .B(_1365_), .C(micro_hash_ucr_pipe56_bF_buf0), .Y(_1367_) );
OAI21X1 OAI21X1_355 ( .gnd(gnd), .vdd(vdd), .A(_460__bF_buf2), .B(_890__bF_buf4), .C(_886_), .Y(_1368_) );
AOI21X1 AOI21X1_266 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe57_bF_buf0), .B(_1283_), .C(micro_hash_ucr_pipe58_bF_buf4), .Y(_1369_) );
OAI21X1 OAI21X1_356 ( .gnd(gnd), .vdd(vdd), .A(_1367_), .B(_1368_), .C(_1369_), .Y(_1370_) );
NAND2X1 NAND2X1_146 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_3_), .B(micro_hash_ucr_pipe58_bF_buf3), .Y(_1371_) );
AOI21X1 AOI21X1_267 ( .gnd(gnd), .vdd(vdd), .A(_1371_), .B(_1370_), .C(micro_hash_ucr_pipe59), .Y(_1372_) );
OAI21X1 OAI21X1_357 ( .gnd(gnd), .vdd(vdd), .A(_1283_), .B(_887__bF_buf3), .C(_883__bF_buf3), .Y(_1373_) );
AOI21X1 AOI21X1_268 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe60_bF_buf0), .B(_460__bF_buf1), .C(micro_hash_ucr_pipe61_bF_buf3), .Y(_1374_) );
OAI21X1 OAI21X1_358 ( .gnd(gnd), .vdd(vdd), .A(_1372_), .B(_1373_), .C(_1374_), .Y(_1375_) );
OAI21X1 OAI21X1_359 ( .gnd(gnd), .vdd(vdd), .A(_885_), .B(_1283_), .C(_1375_), .Y(_1376_) );
AND2X2 AND2X2_187 ( .gnd(gnd), .vdd(vdd), .A(_1376_), .B(_884__bF_buf3), .Y(_1377_) );
OAI21X1 OAI21X1_360 ( .gnd(gnd), .vdd(vdd), .A(_1377_), .B(_1280_), .C(_880__bF_buf1), .Y(_1378_) );
NAND2X1 NAND2X1_147 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe63), .B(_1290__bF_buf3), .Y(_1379_) );
AOI21X1 AOI21X1_269 ( .gnd(gnd), .vdd(vdd), .A(_1379_), .B(_1378_), .C(micro_hash_ucr_pipe64_bF_buf2), .Y(_1380_) );
OAI21X1 OAI21X1_361 ( .gnd(gnd), .vdd(vdd), .A(_1380_), .B(_1279_), .C(_881_), .Y(_1381_) );
AOI21X1 AOI21X1_270 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe65_bF_buf1), .B(_1290__bF_buf2), .C(micro_hash_ucr_pipe66_bF_buf0), .Y(_1382_) );
OAI21X1 OAI21X1_362 ( .gnd(gnd), .vdd(vdd), .A(_877__bF_buf3), .B(micro_hash_ucr_a_3_), .C(_879__bF_buf2), .Y(_1383_) );
AOI21X1 AOI21X1_271 ( .gnd(gnd), .vdd(vdd), .A(_1382_), .B(_1381_), .C(_1383_), .Y(_1384_) );
OAI21X1 OAI21X1_363 ( .gnd(gnd), .vdd(vdd), .A(_1283_), .B(_879__bF_buf1), .C(_878__bF_buf4), .Y(_1385_) );
OAI22X1 OAI22X1_27 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_3_), .B(_878__bF_buf3), .C(_1384_), .D(_1385_), .Y(_1386_) );
OAI21X1 OAI21X1_364 ( .gnd(gnd), .vdd(vdd), .A(_1290__bF_buf1), .B(_876__bF_buf1), .C(_302__bF_buf11), .Y(_1387_) );
AOI21X1 AOI21X1_272 ( .gnd(gnd), .vdd(vdd), .A(_876__bF_buf0), .B(_1386_), .C(_1387_), .Y(_297__3_) );
NAND2X1 NAND2X1_148 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe64_bF_buf1), .B(_474__bF_buf2), .Y(_1388_) );
NOR2X1 NOR2X1_288 ( .gnd(gnd), .vdd(vdd), .A(_474__bF_buf1), .B(_895__bF_buf3), .Y(_1389_) );
NOR2X1 NOR2X1_289 ( .gnd(gnd), .vdd(vdd), .A(_474__bF_buf0), .B(_900__bF_buf2), .Y(_1390_) );
NAND2X1 NAND2X1_149 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe36_bF_buf1), .B(_474__bF_buf3), .Y(_1391_) );
NAND2X1 NAND2X1_150 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe34_bF_buf2), .B(_474__bF_buf2), .Y(_1392_) );
NAND2X1 NAND2X1_151 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe32_bF_buf2), .B(_474__bF_buf1), .Y(_1393_) );
INVX1 INVX1_102 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_4_), .Y(_1394_) );
INVX8 INVX8_81 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_4_bF_buf1_), .Y(_1395_) );
NAND2X1 NAND2X1_152 ( .gnd(gnd), .vdd(vdd), .A(_1394_), .B(_1395_), .Y(_1396_) );
NAND2X1 NAND2X1_153 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_4_), .B(micro_hash_ucr_b_4_bF_buf0_), .Y(_1397_) );
NAND2X1 NAND2X1_154 ( .gnd(gnd), .vdd(vdd), .A(_1397_), .B(_1396_), .Y(_1398_) );
NAND2X1 NAND2X1_155 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_4_), .B(micro_hash_ucr_pipe22_bF_buf3), .Y(_1399_) );
NAND2X1 NAND2X1_156 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_4_), .B(micro_hash_ucr_pipe20_bF_buf4), .Y(_1400_) );
NAND2X1 NAND2X1_157 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_4_), .B(micro_hash_ucr_pipe18_bF_buf1), .Y(_1401_) );
INVX8 INVX8_82 ( .gnd(gnd), .vdd(vdd), .A(_1398_), .Y(_1402_) );
INVX1 INVX1_103 ( .gnd(gnd), .vdd(vdd), .A(_1296_), .Y(_1403_) );
NOR2X1 NOR2X1_290 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe9), .B(_1403_), .Y(_1404_) );
NAND3X1 NAND3X1_35 ( .gnd(gnd), .vdd(vdd), .A(_471_), .B(_939_), .C(_1187_), .Y(_1405_) );
NOR2X1 NOR2X1_291 ( .gnd(gnd), .vdd(vdd), .A(_1295_), .B(_1405_), .Y(_1406_) );
NAND2X1 NAND2X1_158 ( .gnd(gnd), .vdd(vdd), .A(_1404_), .B(_1406_), .Y(_1407_) );
OAI21X1 OAI21X1_365 ( .gnd(gnd), .vdd(vdd), .A(_1070_), .B(_1402__bF_buf3), .C(_1407_), .Y(_1408_) );
AND2X2 AND2X2_188 ( .gnd(gnd), .vdd(vdd), .A(_1408_), .B(_932_), .Y(_1409_) );
OAI21X1 OAI21X1_366 ( .gnd(gnd), .vdd(vdd), .A(_1079_), .B(micro_hash_ucr_a_4_), .C(_928_), .Y(_1410_) );
OAI22X1 OAI22X1_28 ( .gnd(gnd), .vdd(vdd), .A(_928_), .B(_1398_), .C(_1409_), .D(_1410_), .Y(_1411_) );
NAND2X1 NAND2X1_159 ( .gnd(gnd), .vdd(vdd), .A(_930__bF_buf0), .B(_1411_), .Y(_1412_) );
OAI21X1 OAI21X1_367 ( .gnd(gnd), .vdd(vdd), .A(_474__bF_buf0), .B(_930__bF_buf4), .C(_1412_), .Y(_1413_) );
NAND2X1 NAND2X1_160 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe17_bF_buf1), .B(_1398_), .Y(_1414_) );
OAI21X1 OAI21X1_368 ( .gnd(gnd), .vdd(vdd), .A(_1413_), .B(micro_hash_ucr_pipe17_bF_buf0), .C(_1414_), .Y(_1415_) );
OAI21X1 OAI21X1_369 ( .gnd(gnd), .vdd(vdd), .A(_1415_), .B(micro_hash_ucr_pipe18_bF_buf0), .C(_1401_), .Y(_1416_) );
NAND2X1 NAND2X1_161 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe19_bF_buf2), .B(_1398_), .Y(_1417_) );
OAI21X1 OAI21X1_370 ( .gnd(gnd), .vdd(vdd), .A(_1416_), .B(micro_hash_ucr_pipe19_bF_buf1), .C(_1417_), .Y(_1418_) );
OAI21X1 OAI21X1_371 ( .gnd(gnd), .vdd(vdd), .A(_1418_), .B(micro_hash_ucr_pipe20_bF_buf3), .C(_1400_), .Y(_1419_) );
NAND2X1 NAND2X1_162 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe21_bF_buf2), .B(_1398_), .Y(_1420_) );
OAI21X1 OAI21X1_372 ( .gnd(gnd), .vdd(vdd), .A(_1419_), .B(micro_hash_ucr_pipe21_bF_buf1), .C(_1420_), .Y(_1421_) );
OAI21X1 OAI21X1_373 ( .gnd(gnd), .vdd(vdd), .A(_1421_), .B(micro_hash_ucr_pipe22_bF_buf2), .C(_1399_), .Y(_1422_) );
NAND2X1 NAND2X1_163 ( .gnd(gnd), .vdd(vdd), .A(_923_), .B(_1422_), .Y(_1423_) );
OAI21X1 OAI21X1_374 ( .gnd(gnd), .vdd(vdd), .A(_923_), .B(_1398_), .C(_1423_), .Y(_1424_) );
AOI21X1 AOI21X1_273 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe24_bF_buf3), .B(_474__bF_buf3), .C(micro_hash_ucr_pipe25), .Y(_1425_) );
OAI21X1 OAI21X1_375 ( .gnd(gnd), .vdd(vdd), .A(_1424_), .B(micro_hash_ucr_pipe24_bF_buf2), .C(_1425_), .Y(_1426_) );
OAI21X1 OAI21X1_376 ( .gnd(gnd), .vdd(vdd), .A(_921__bF_buf0), .B(_1398_), .C(_1426_), .Y(_1427_) );
NAND2X1 NAND2X1_164 ( .gnd(gnd), .vdd(vdd), .A(_920__bF_buf2), .B(_1427_), .Y(_1428_) );
OAI21X1 OAI21X1_377 ( .gnd(gnd), .vdd(vdd), .A(_474__bF_buf2), .B(_920__bF_buf1), .C(_1428_), .Y(_1429_) );
OAI21X1 OAI21X1_378 ( .gnd(gnd), .vdd(vdd), .A(_1398_), .B(_916_), .C(_918__bF_buf3), .Y(_1430_) );
AOI21X1 AOI21X1_274 ( .gnd(gnd), .vdd(vdd), .A(_916_), .B(_1429_), .C(_1430_), .Y(_1431_) );
OAI21X1 OAI21X1_379 ( .gnd(gnd), .vdd(vdd), .A(_918__bF_buf2), .B(micro_hash_ucr_a_4_), .C(_917_), .Y(_1432_) );
AOI21X1 AOI21X1_275 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe29_bF_buf0), .B(_1402__bF_buf2), .C(micro_hash_ucr_pipe30_bF_buf3), .Y(_1433_) );
OAI21X1 OAI21X1_380 ( .gnd(gnd), .vdd(vdd), .A(_1431_), .B(_1432_), .C(_1433_), .Y(_1434_) );
NAND2X1 NAND2X1_165 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe30_bF_buf2), .B(_474__bF_buf1), .Y(_1435_) );
AOI21X1 AOI21X1_276 ( .gnd(gnd), .vdd(vdd), .A(_1435_), .B(_1434_), .C(micro_hash_ucr_pipe31), .Y(_1436_) );
NOR2X1 NOR2X1_292 ( .gnd(gnd), .vdd(vdd), .A(_915__bF_buf0), .B(_1402__bF_buf1), .Y(_1437_) );
OAI21X1 OAI21X1_381 ( .gnd(gnd), .vdd(vdd), .A(_1436_), .B(_1437_), .C(_914__bF_buf0), .Y(_1438_) );
AOI21X1 AOI21X1_277 ( .gnd(gnd), .vdd(vdd), .A(_1393_), .B(_1438_), .C(micro_hash_ucr_pipe33_bF_buf2), .Y(_1439_) );
NOR2X1 NOR2X1_293 ( .gnd(gnd), .vdd(vdd), .A(_910_), .B(_1402__bF_buf0), .Y(_1440_) );
OAI21X1 OAI21X1_382 ( .gnd(gnd), .vdd(vdd), .A(_1439_), .B(_1440_), .C(_912__bF_buf4), .Y(_1441_) );
AOI21X1 AOI21X1_278 ( .gnd(gnd), .vdd(vdd), .A(_1392_), .B(_1441_), .C(micro_hash_ucr_pipe35), .Y(_1442_) );
NOR2X1 NOR2X1_294 ( .gnd(gnd), .vdd(vdd), .A(_911__bF_buf2), .B(_1402__bF_buf3), .Y(_1443_) );
OAI21X1 OAI21X1_383 ( .gnd(gnd), .vdd(vdd), .A(_1442_), .B(_1443_), .C(_907__bF_buf0), .Y(_1444_) );
NAND3X1 NAND3X1_36 ( .gnd(gnd), .vdd(vdd), .A(_909__bF_buf1), .B(_1391_), .C(_1444_), .Y(_1445_) );
AOI21X1 AOI21X1_279 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe37), .B(_1402__bF_buf2), .C(micro_hash_ucr_pipe38_bF_buf3), .Y(_1446_) );
OAI21X1 OAI21X1_384 ( .gnd(gnd), .vdd(vdd), .A(_908__bF_buf3), .B(micro_hash_ucr_a_4_), .C(_904__bF_buf0), .Y(_1447_) );
AOI21X1 AOI21X1_280 ( .gnd(gnd), .vdd(vdd), .A(_1446_), .B(_1445_), .C(_1447_), .Y(_1448_) );
OAI21X1 OAI21X1_385 ( .gnd(gnd), .vdd(vdd), .A(_1398_), .B(_904__bF_buf3), .C(_906__bF_buf4), .Y(_1449_) );
OAI22X1 OAI22X1_29 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_4_), .B(_906__bF_buf3), .C(_1448_), .D(_1449_), .Y(_1450_) );
NOR2X1 NOR2X1_295 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe41), .B(_1450_), .Y(_1451_) );
NOR2X1 NOR2X1_296 ( .gnd(gnd), .vdd(vdd), .A(_905__bF_buf1), .B(_1398_), .Y(_1452_) );
OAI21X1 OAI21X1_386 ( .gnd(gnd), .vdd(vdd), .A(_1451_), .B(_1452_), .C(_901__bF_buf1), .Y(_1453_) );
AOI21X1 AOI21X1_281 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_4_), .B(micro_hash_ucr_pipe42_bF_buf1), .C(micro_hash_ucr_pipe43), .Y(_1454_) );
OAI21X1 OAI21X1_387 ( .gnd(gnd), .vdd(vdd), .A(_1402__bF_buf1), .B(_903__bF_buf3), .C(_902__bF_buf1), .Y(_1455_) );
AOI21X1 AOI21X1_282 ( .gnd(gnd), .vdd(vdd), .A(_1454_), .B(_1453_), .C(_1455_), .Y(_1456_) );
NOR2X1 NOR2X1_297 ( .gnd(gnd), .vdd(vdd), .A(_474__bF_buf0), .B(_902__bF_buf0), .Y(_1457_) );
OAI21X1 OAI21X1_388 ( .gnd(gnd), .vdd(vdd), .A(_1456_), .B(_1457_), .C(_898_), .Y(_1458_) );
NAND2X1 NAND2X1_166 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe45_bF_buf3), .B(_1402__bF_buf0), .Y(_1459_) );
AOI21X1 AOI21X1_283 ( .gnd(gnd), .vdd(vdd), .A(_1459_), .B(_1458_), .C(micro_hash_ucr_pipe46_bF_buf4), .Y(_1460_) );
OAI21X1 OAI21X1_389 ( .gnd(gnd), .vdd(vdd), .A(_1460_), .B(_1390_), .C(_899__bF_buf1), .Y(_1461_) );
NAND2X1 NAND2X1_167 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe47), .B(_1402__bF_buf3), .Y(_1462_) );
AOI21X1 AOI21X1_284 ( .gnd(gnd), .vdd(vdd), .A(_1462_), .B(_1461_), .C(micro_hash_ucr_pipe48_bF_buf3), .Y(_1463_) );
OAI21X1 OAI21X1_390 ( .gnd(gnd), .vdd(vdd), .A(_1463_), .B(_1389_), .C(_897__bF_buf1), .Y(_1464_) );
AOI21X1 AOI21X1_285 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe49), .B(_1402__bF_buf2), .C(micro_hash_ucr_pipe50_bF_buf2), .Y(_1465_) );
OAI21X1 OAI21X1_391 ( .gnd(gnd), .vdd(vdd), .A(_896__bF_buf4), .B(micro_hash_ucr_a_4_), .C(_892_), .Y(_1466_) );
AOI21X1 AOI21X1_286 ( .gnd(gnd), .vdd(vdd), .A(_1465_), .B(_1464_), .C(_1466_), .Y(_1467_) );
OAI21X1 OAI21X1_392 ( .gnd(gnd), .vdd(vdd), .A(_1398_), .B(_892_), .C(_894__bF_buf1), .Y(_1468_) );
OAI22X1 OAI22X1_30 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_4_), .B(_894__bF_buf0), .C(_1467_), .D(_1468_), .Y(_1469_) );
NAND2X1 NAND2X1_168 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe53_bF_buf3), .B(_1402__bF_buf1), .Y(_1470_) );
OAI21X1 OAI21X1_393 ( .gnd(gnd), .vdd(vdd), .A(_1469_), .B(micro_hash_ucr_pipe53_bF_buf2), .C(_1470_), .Y(_1471_) );
NAND2X1 NAND2X1_169 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe54_bF_buf3), .B(_474__bF_buf3), .Y(_1472_) );
OAI21X1 OAI21X1_394 ( .gnd(gnd), .vdd(vdd), .A(_1471_), .B(micro_hash_ucr_pipe54_bF_buf2), .C(_1472_), .Y(_1473_) );
NAND2X1 NAND2X1_170 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe55), .B(_1402__bF_buf0), .Y(_1474_) );
OAI21X1 OAI21X1_395 ( .gnd(gnd), .vdd(vdd), .A(_1473_), .B(micro_hash_ucr_pipe55), .C(_1474_), .Y(_1475_) );
OAI21X1 OAI21X1_396 ( .gnd(gnd), .vdd(vdd), .A(_474__bF_buf2), .B(_890__bF_buf3), .C(_886_), .Y(_1476_) );
AOI21X1 AOI21X1_287 ( .gnd(gnd), .vdd(vdd), .A(_890__bF_buf2), .B(_1475_), .C(_1476_), .Y(_1477_) );
OAI21X1 OAI21X1_397 ( .gnd(gnd), .vdd(vdd), .A(_1402__bF_buf3), .B(_886_), .C(_888__bF_buf0), .Y(_1478_) );
OAI22X1 OAI22X1_31 ( .gnd(gnd), .vdd(vdd), .A(_474__bF_buf1), .B(_888__bF_buf3), .C(_1477_), .D(_1478_), .Y(_1479_) );
OAI21X1 OAI21X1_398 ( .gnd(gnd), .vdd(vdd), .A(_1398_), .B(_887__bF_buf2), .C(_883__bF_buf2), .Y(_1480_) );
AOI21X1 AOI21X1_288 ( .gnd(gnd), .vdd(vdd), .A(_887__bF_buf1), .B(_1479_), .C(_1480_), .Y(_1481_) );
OAI21X1 OAI21X1_399 ( .gnd(gnd), .vdd(vdd), .A(_883__bF_buf1), .B(micro_hash_ucr_a_4_), .C(_885_), .Y(_1482_) );
AOI21X1 AOI21X1_289 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe61_bF_buf2), .B(_1402__bF_buf2), .C(micro_hash_ucr_pipe62_bF_buf1), .Y(_1483_) );
OAI21X1 OAI21X1_400 ( .gnd(gnd), .vdd(vdd), .A(_1481_), .B(_1482_), .C(_1483_), .Y(_1484_) );
NAND2X1 NAND2X1_171 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe62_bF_buf0), .B(_474__bF_buf0), .Y(_1485_) );
AOI21X1 AOI21X1_290 ( .gnd(gnd), .vdd(vdd), .A(_1485_), .B(_1484_), .C(micro_hash_ucr_pipe63), .Y(_1486_) );
NOR2X1 NOR2X1_298 ( .gnd(gnd), .vdd(vdd), .A(_880__bF_buf0), .B(_1402__bF_buf1), .Y(_1487_) );
OAI21X1 OAI21X1_401 ( .gnd(gnd), .vdd(vdd), .A(_1486_), .B(_1487_), .C(_882__bF_buf0), .Y(_1488_) );
NAND3X1 NAND3X1_37 ( .gnd(gnd), .vdd(vdd), .A(_881_), .B(_1388_), .C(_1488_), .Y(_1489_) );
NAND2X1 NAND2X1_172 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe65_bF_buf0), .B(_1402__bF_buf0), .Y(_1490_) );
AOI21X1 AOI21X1_291 ( .gnd(gnd), .vdd(vdd), .A(_1490_), .B(_1489_), .C(micro_hash_ucr_pipe66_bF_buf4), .Y(_1491_) );
OAI21X1 OAI21X1_402 ( .gnd(gnd), .vdd(vdd), .A(_474__bF_buf3), .B(_877__bF_buf2), .C(_879__bF_buf0), .Y(_1492_) );
AOI21X1 AOI21X1_292 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe67), .B(_1398_), .C(micro_hash_ucr_pipe68), .Y(_1493_) );
OAI21X1 OAI21X1_403 ( .gnd(gnd), .vdd(vdd), .A(_1491_), .B(_1492_), .C(_1493_), .Y(_1494_) );
AOI21X1 AOI21X1_293 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_4_), .B(micro_hash_ucr_pipe68), .C(micro_hash_ucr_pipe69), .Y(_1495_) );
OAI21X1 OAI21X1_404 ( .gnd(gnd), .vdd(vdd), .A(_1402__bF_buf3), .B(_876__bF_buf3), .C(_302__bF_buf10), .Y(_1496_) );
AOI21X1 AOI21X1_294 ( .gnd(gnd), .vdd(vdd), .A(_1495_), .B(_1494_), .C(_1496_), .Y(_297__4_) );
NAND2X1 NAND2X1_173 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_5_bF_buf1_), .B(micro_hash_ucr_pipe66_bF_buf3), .Y(_1497_) );
NAND2X1 NAND2X1_174 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_5_bF_buf0_), .B(micro_hash_ucr_pipe64_bF_buf0), .Y(_1498_) );
NAND2X1 NAND2X1_175 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_5_bF_buf3_), .B(micro_hash_ucr_pipe62_bF_buf4), .Y(_1499_) );
NAND2X1 NAND2X1_176 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_5_bF_buf2_), .B(micro_hash_ucr_pipe54_bF_buf1), .Y(_1500_) );
NOR2X1 NOR2X1_299 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_5_), .B(micro_hash_ucr_b_5_bF_buf1_), .Y(_1501_) );
NOR2X1 NOR2X1_300 ( .gnd(gnd), .vdd(vdd), .A(_4460_), .B(_414__bF_buf2), .Y(_1502_) );
NOR2X1 NOR2X1_301 ( .gnd(gnd), .vdd(vdd), .A(_1501_), .B(_1502_), .Y(_1503_) );
INVX8 INVX8_83 ( .gnd(gnd), .vdd(vdd), .A(_1503_), .Y(_1504_) );
NAND2X1 NAND2X1_177 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_5_bF_buf1_), .B(micro_hash_ucr_pipe42_bF_buf0), .Y(_1505_) );
NAND2X1 NAND2X1_178 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_5_bF_buf0_), .B(micro_hash_ucr_pipe40_bF_buf4), .Y(_1506_) );
NOR2X1 NOR2X1_302 ( .gnd(gnd), .vdd(vdd), .A(_480_), .B(_912__bF_buf3), .Y(_1507_) );
NOR2X1 NOR2X1_303 ( .gnd(gnd), .vdd(vdd), .A(_480_), .B(_914__bF_buf4), .Y(_1508_) );
NOR2X1 NOR2X1_304 ( .gnd(gnd), .vdd(vdd), .A(_480_), .B(_913__bF_buf3), .Y(_1509_) );
NOR2X1 NOR2X1_305 ( .gnd(gnd), .vdd(vdd), .A(_480_), .B(_924__bF_buf4), .Y(_1510_) );
NOR2X1 NOR2X1_306 ( .gnd(gnd), .vdd(vdd), .A(_480_), .B(_926__bF_buf3), .Y(_1511_) );
NOR2X1 NOR2X1_307 ( .gnd(gnd), .vdd(vdd), .A(_480_), .B(_925__bF_buf1), .Y(_1512_) );
NOR2X1 NOR2X1_308 ( .gnd(gnd), .vdd(vdd), .A(_480_), .B(_930__bF_buf3), .Y(_1513_) );
NAND2X1 NAND2X1_179 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe15_bF_buf2), .B(_1503_), .Y(_1514_) );
NAND2X1 NAND2X1_180 ( .gnd(gnd), .vdd(vdd), .A(_928_), .B(_1070_), .Y(_1515_) );
NAND3X1 NAND3X1_38 ( .gnd(gnd), .vdd(vdd), .A(_479_), .B(_939_), .C(_1187_), .Y(_1516_) );
NOR2X1 NOR2X1_309 ( .gnd(gnd), .vdd(vdd), .A(_1295_), .B(_1516_), .Y(_1517_) );
AOI22X1 AOI22X1_17 ( .gnd(gnd), .vdd(vdd), .A(_1404_), .B(_1517_), .C(_1515_), .D(_1504_), .Y(_1518_) );
NOR2X1 NOR2X1_310 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe15_bF_buf1), .B(_932_), .Y(_1519_) );
OAI22X1 OAI22X1_32 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_5_bF_buf3_), .B(_1079_), .C(_1518_), .D(_1519_), .Y(_1520_) );
AOI21X1 AOI21X1_295 ( .gnd(gnd), .vdd(vdd), .A(_1514_), .B(_1520_), .C(micro_hash_ucr_pipe16_bF_buf0), .Y(_1521_) );
OAI21X1 OAI21X1_405 ( .gnd(gnd), .vdd(vdd), .A(_1521_), .B(_1513_), .C(_929_), .Y(_1522_) );
NAND2X1 NAND2X1_181 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe17_bF_buf3), .B(_1503_), .Y(_1523_) );
AOI21X1 AOI21X1_296 ( .gnd(gnd), .vdd(vdd), .A(_1523_), .B(_1522_), .C(micro_hash_ucr_pipe18_bF_buf4), .Y(_1524_) );
OAI21X1 OAI21X1_406 ( .gnd(gnd), .vdd(vdd), .A(_1524_), .B(_1512_), .C(_927__bF_buf1), .Y(_1525_) );
NAND2X1 NAND2X1_182 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe19_bF_buf0), .B(_1503_), .Y(_1526_) );
AOI21X1 AOI21X1_297 ( .gnd(gnd), .vdd(vdd), .A(_1526_), .B(_1525_), .C(micro_hash_ucr_pipe20_bF_buf2), .Y(_1527_) );
OAI21X1 OAI21X1_407 ( .gnd(gnd), .vdd(vdd), .A(_1527_), .B(_1511_), .C(_922_), .Y(_1528_) );
NAND2X1 NAND2X1_183 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe21_bF_buf0), .B(_1503_), .Y(_1529_) );
AOI21X1 AOI21X1_298 ( .gnd(gnd), .vdd(vdd), .A(_1529_), .B(_1528_), .C(micro_hash_ucr_pipe22_bF_buf1), .Y(_1530_) );
OAI21X1 OAI21X1_408 ( .gnd(gnd), .vdd(vdd), .A(_1530_), .B(_1510_), .C(_923_), .Y(_1531_) );
AOI21X1 AOI21X1_299 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe23_bF_buf0), .B(_1503_), .C(micro_hash_ucr_pipe24_bF_buf1), .Y(_1532_) );
OAI21X1 OAI21X1_409 ( .gnd(gnd), .vdd(vdd), .A(_919__bF_buf4), .B(micro_hash_ucr_a_5_bF_buf2_), .C(_921__bF_buf3), .Y(_1533_) );
AOI21X1 AOI21X1_300 ( .gnd(gnd), .vdd(vdd), .A(_1532_), .B(_1531_), .C(_1533_), .Y(_1534_) );
OAI21X1 OAI21X1_410 ( .gnd(gnd), .vdd(vdd), .A(_1504_), .B(_921__bF_buf2), .C(_920__bF_buf0), .Y(_1535_) );
OAI22X1 OAI22X1_33 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_5_bF_buf1_), .B(_920__bF_buf4), .C(_1534_), .D(_1535_), .Y(_1536_) );
OAI21X1 OAI21X1_411 ( .gnd(gnd), .vdd(vdd), .A(_1503_), .B(_916_), .C(_918__bF_buf1), .Y(_1537_) );
AOI21X1 AOI21X1_301 ( .gnd(gnd), .vdd(vdd), .A(_916_), .B(_1536_), .C(_1537_), .Y(_1538_) );
NOR2X1 NOR2X1_311 ( .gnd(gnd), .vdd(vdd), .A(_480_), .B(_918__bF_buf0), .Y(_1539_) );
OAI21X1 OAI21X1_412 ( .gnd(gnd), .vdd(vdd), .A(_1538_), .B(_1539_), .C(_917_), .Y(_1540_) );
NAND2X1 NAND2X1_184 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe29_bF_buf3), .B(_1503_), .Y(_1541_) );
AOI21X1 AOI21X1_302 ( .gnd(gnd), .vdd(vdd), .A(_1541_), .B(_1540_), .C(micro_hash_ucr_pipe30_bF_buf1), .Y(_1542_) );
OAI21X1 OAI21X1_413 ( .gnd(gnd), .vdd(vdd), .A(_1542_), .B(_1509_), .C(_915__bF_buf3), .Y(_1543_) );
NAND2X1 NAND2X1_185 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe31), .B(_1503_), .Y(_1544_) );
AOI21X1 AOI21X1_303 ( .gnd(gnd), .vdd(vdd), .A(_1544_), .B(_1543_), .C(micro_hash_ucr_pipe32_bF_buf1), .Y(_1545_) );
OAI21X1 OAI21X1_414 ( .gnd(gnd), .vdd(vdd), .A(_1545_), .B(_1508_), .C(_910_), .Y(_1546_) );
NAND2X1 NAND2X1_186 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe33_bF_buf1), .B(_1503_), .Y(_1547_) );
AOI21X1 AOI21X1_304 ( .gnd(gnd), .vdd(vdd), .A(_1547_), .B(_1546_), .C(micro_hash_ucr_pipe34_bF_buf1), .Y(_1548_) );
OAI21X1 OAI21X1_415 ( .gnd(gnd), .vdd(vdd), .A(_1548_), .B(_1507_), .C(_911__bF_buf1), .Y(_1549_) );
OAI21X1 OAI21X1_416 ( .gnd(gnd), .vdd(vdd), .A(_911__bF_buf0), .B(_1504_), .C(_1549_), .Y(_1550_) );
AND2X2 AND2X2_189 ( .gnd(gnd), .vdd(vdd), .A(_1550_), .B(_907__bF_buf4), .Y(_1551_) );
OAI21X1 OAI21X1_417 ( .gnd(gnd), .vdd(vdd), .A(_480_), .B(_907__bF_buf3), .C(_909__bF_buf0), .Y(_1552_) );
AOI21X1 AOI21X1_305 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe37), .B(_1504_), .C(micro_hash_ucr_pipe38_bF_buf2), .Y(_1553_) );
OAI21X1 OAI21X1_418 ( .gnd(gnd), .vdd(vdd), .A(_1551_), .B(_1552_), .C(_1553_), .Y(_1554_) );
NAND2X1 NAND2X1_187 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_5_bF_buf0_), .B(micro_hash_ucr_pipe38_bF_buf1), .Y(_1555_) );
AOI21X1 AOI21X1_306 ( .gnd(gnd), .vdd(vdd), .A(_1555_), .B(_1554_), .C(micro_hash_ucr_pipe39), .Y(_1556_) );
NOR2X1 NOR2X1_312 ( .gnd(gnd), .vdd(vdd), .A(_904__bF_buf2), .B(_1504_), .Y(_1557_) );
OAI21X1 OAI21X1_419 ( .gnd(gnd), .vdd(vdd), .A(_1556_), .B(_1557_), .C(_906__bF_buf2), .Y(_1558_) );
AOI21X1 AOI21X1_307 ( .gnd(gnd), .vdd(vdd), .A(_1506_), .B(_1558_), .C(micro_hash_ucr_pipe41), .Y(_1559_) );
NOR2X1 NOR2X1_313 ( .gnd(gnd), .vdd(vdd), .A(_905__bF_buf0), .B(_1504_), .Y(_1560_) );
OAI21X1 OAI21X1_420 ( .gnd(gnd), .vdd(vdd), .A(_1559_), .B(_1560_), .C(_901__bF_buf0), .Y(_1561_) );
AOI21X1 AOI21X1_308 ( .gnd(gnd), .vdd(vdd), .A(_1505_), .B(_1561_), .C(micro_hash_ucr_pipe43), .Y(_1562_) );
NOR2X1 NOR2X1_314 ( .gnd(gnd), .vdd(vdd), .A(_903__bF_buf2), .B(_1504_), .Y(_1563_) );
OAI21X1 OAI21X1_421 ( .gnd(gnd), .vdd(vdd), .A(_1562_), .B(_1563_), .C(_902__bF_buf4), .Y(_1564_) );
AOI21X1 AOI21X1_309 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_5_bF_buf3_), .B(micro_hash_ucr_pipe44), .C(micro_hash_ucr_pipe45_bF_buf2), .Y(_1565_) );
AOI22X1 AOI22X1_18 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe45_bF_buf1), .B(_1504_), .C(_1564_), .D(_1565_), .Y(_1566_) );
AOI21X1 AOI21X1_310 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe46_bF_buf3), .B(_480_), .C(micro_hash_ucr_pipe47), .Y(_1567_) );
OAI21X1 OAI21X1_422 ( .gnd(gnd), .vdd(vdd), .A(_1566_), .B(micro_hash_ucr_pipe46_bF_buf2), .C(_1567_), .Y(_1568_) );
AOI21X1 AOI21X1_311 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe47), .B(_1503_), .C(micro_hash_ucr_pipe48_bF_buf2), .Y(_1569_) );
NAND2X1 NAND2X1_188 ( .gnd(gnd), .vdd(vdd), .A(_1569_), .B(_1568_), .Y(_1570_) );
NAND2X1 NAND2X1_189 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe48_bF_buf1), .B(_480_), .Y(_1571_) );
NAND3X1 NAND3X1_39 ( .gnd(gnd), .vdd(vdd), .A(_897__bF_buf0), .B(_1571_), .C(_1570_), .Y(_1572_) );
NAND2X1 NAND2X1_190 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe49), .B(_1503_), .Y(_1573_) );
AOI21X1 AOI21X1_312 ( .gnd(gnd), .vdd(vdd), .A(_1573_), .B(_1572_), .C(micro_hash_ucr_pipe50_bF_buf1), .Y(_1574_) );
OAI21X1 OAI21X1_423 ( .gnd(gnd), .vdd(vdd), .A(_480_), .B(_896__bF_buf3), .C(_892_), .Y(_1575_) );
AOI21X1 AOI21X1_313 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe51), .B(_1504_), .C(micro_hash_ucr_pipe52_bF_buf0), .Y(_1576_) );
OAI21X1 OAI21X1_424 ( .gnd(gnd), .vdd(vdd), .A(_1574_), .B(_1575_), .C(_1576_), .Y(_1577_) );
NAND2X1 NAND2X1_191 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_5_bF_buf2_), .B(micro_hash_ucr_pipe52_bF_buf4), .Y(_1578_) );
NAND3X1 NAND3X1_40 ( .gnd(gnd), .vdd(vdd), .A(_893_), .B(_1578_), .C(_1577_), .Y(_1579_) );
OAI21X1 OAI21X1_425 ( .gnd(gnd), .vdd(vdd), .A(_1502_), .B(_1501_), .C(micro_hash_ucr_pipe53_bF_buf1), .Y(_1580_) );
NAND3X1 NAND3X1_41 ( .gnd(gnd), .vdd(vdd), .A(_889__bF_buf3), .B(_1580_), .C(_1579_), .Y(_1581_) );
AOI21X1 AOI21X1_314 ( .gnd(gnd), .vdd(vdd), .A(_1500_), .B(_1581_), .C(micro_hash_ucr_pipe55), .Y(_1582_) );
OAI21X1 OAI21X1_426 ( .gnd(gnd), .vdd(vdd), .A(_1504_), .B(_891_), .C(_890__bF_buf1), .Y(_1583_) );
AOI21X1 AOI21X1_315 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe56_bF_buf3), .B(_480_), .C(micro_hash_ucr_pipe57_bF_buf3), .Y(_1584_) );
OAI21X1 OAI21X1_427 ( .gnd(gnd), .vdd(vdd), .A(_1582_), .B(_1583_), .C(_1584_), .Y(_1585_) );
AOI21X1 AOI21X1_316 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe57_bF_buf2), .B(_1503_), .C(micro_hash_ucr_pipe58_bF_buf2), .Y(_1586_) );
AOI22X1 AOI22X1_19 ( .gnd(gnd), .vdd(vdd), .A(_480_), .B(micro_hash_ucr_pipe58_bF_buf1), .C(_1585_), .D(_1586_), .Y(_1587_) );
AOI21X1 AOI21X1_317 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe59), .B(_1504_), .C(micro_hash_ucr_pipe60_bF_buf4), .Y(_1588_) );
OAI21X1 OAI21X1_428 ( .gnd(gnd), .vdd(vdd), .A(_1587_), .B(micro_hash_ucr_pipe59), .C(_1588_), .Y(_1589_) );
NAND2X1 NAND2X1_192 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_5_bF_buf1_), .B(micro_hash_ucr_pipe60_bF_buf3), .Y(_1590_) );
NAND3X1 NAND3X1_42 ( .gnd(gnd), .vdd(vdd), .A(_885_), .B(_1590_), .C(_1589_), .Y(_1591_) );
OAI21X1 OAI21X1_429 ( .gnd(gnd), .vdd(vdd), .A(_1502_), .B(_1501_), .C(micro_hash_ucr_pipe61_bF_buf1), .Y(_1592_) );
NAND3X1 NAND3X1_43 ( .gnd(gnd), .vdd(vdd), .A(_884__bF_buf2), .B(_1592_), .C(_1591_), .Y(_1593_) );
NAND3X1 NAND3X1_44 ( .gnd(gnd), .vdd(vdd), .A(_880__bF_buf3), .B(_1499_), .C(_1593_), .Y(_1594_) );
OAI21X1 OAI21X1_430 ( .gnd(gnd), .vdd(vdd), .A(_1502_), .B(_1501_), .C(micro_hash_ucr_pipe63), .Y(_1595_) );
NAND3X1 NAND3X1_45 ( .gnd(gnd), .vdd(vdd), .A(_882__bF_buf3), .B(_1595_), .C(_1594_), .Y(_1596_) );
NAND3X1 NAND3X1_46 ( .gnd(gnd), .vdd(vdd), .A(_881_), .B(_1498_), .C(_1596_), .Y(_1597_) );
OAI21X1 OAI21X1_431 ( .gnd(gnd), .vdd(vdd), .A(_1502_), .B(_1501_), .C(micro_hash_ucr_pipe65_bF_buf3), .Y(_1598_) );
NAND3X1 NAND3X1_47 ( .gnd(gnd), .vdd(vdd), .A(_877__bF_buf1), .B(_1598_), .C(_1597_), .Y(_1599_) );
NAND3X1 NAND3X1_48 ( .gnd(gnd), .vdd(vdd), .A(_879__bF_buf3), .B(_1497_), .C(_1599_), .Y(_1600_) );
OAI21X1 OAI21X1_432 ( .gnd(gnd), .vdd(vdd), .A(_1502_), .B(_1501_), .C(micro_hash_ucr_pipe67), .Y(_1601_) );
NAND3X1 NAND3X1_49 ( .gnd(gnd), .vdd(vdd), .A(_878__bF_buf2), .B(_1601_), .C(_1600_), .Y(_1602_) );
AOI21X1 AOI21X1_318 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_5_bF_buf0_), .B(micro_hash_ucr_pipe68), .C(micro_hash_ucr_pipe69), .Y(_1603_) );
OAI21X1 OAI21X1_433 ( .gnd(gnd), .vdd(vdd), .A(_1503_), .B(_876__bF_buf2), .C(_302__bF_buf9), .Y(_1604_) );
AOI21X1 AOI21X1_319 ( .gnd(gnd), .vdd(vdd), .A(_1603_), .B(_1602_), .C(_1604_), .Y(_297__5_) );
NAND2X1 NAND2X1_193 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_6_bF_buf1_), .B(micro_hash_ucr_pipe66_bF_buf2), .Y(_1605_) );
NAND2X1 NAND2X1_194 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_6_bF_buf0_), .B(micro_hash_ucr_pipe64_bF_buf4), .Y(_1606_) );
NAND2X1 NAND2X1_195 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_6_bF_buf3_), .B(micro_hash_ucr_pipe62_bF_buf3), .Y(_1607_) );
NAND2X1 NAND2X1_196 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_6_bF_buf2_), .B(micro_hash_ucr_pipe52_bF_buf3), .Y(_1608_) );
NAND2X1 NAND2X1_197 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_6_bF_buf1_), .B(micro_hash_ucr_pipe50_bF_buf0), .Y(_1609_) );
NAND2X1 NAND2X1_198 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_6_bF_buf0_), .B(micro_hash_ucr_pipe48_bF_buf0), .Y(_1610_) );
NAND2X1 NAND2X1_199 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_6_bF_buf3_), .B(micro_hash_ucr_pipe46_bF_buf1), .Y(_1611_) );
NAND2X1 NAND2X1_200 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_6_bF_buf2_), .B(micro_hash_ucr_pipe44), .Y(_1612_) );
NAND2X1 NAND2X1_201 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe32_bF_buf0), .B(_494_), .Y(_1613_) );
NOR2X1 NOR2X1_315 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_6_), .B(micro_hash_ucr_b_6_bF_buf1_), .Y(_1614_) );
NOR2X1 NOR2X1_316 ( .gnd(gnd), .vdd(vdd), .A(_4472_), .B(_428__bF_buf2), .Y(_1615_) );
NOR2X1 NOR2X1_317 ( .gnd(gnd), .vdd(vdd), .A(_1614_), .B(_1615_), .Y(_1616_) );
INVX4 INVX4_52 ( .gnd(gnd), .vdd(vdd), .A(_1616_), .Y(_1617_) );
NOR2X1 NOR2X1_318 ( .gnd(gnd), .vdd(vdd), .A(_494_), .B(_926__bF_buf2), .Y(_1618_) );
NOR2X1 NOR2X1_319 ( .gnd(gnd), .vdd(vdd), .A(_494_), .B(_925__bF_buf0), .Y(_1619_) );
NAND2X1 NAND2X1_202 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe15_bF_buf0), .B(_1616_), .Y(_1620_) );
NOR2X1 NOR2X1_320 ( .gnd(gnd), .vdd(vdd), .A(H_6_), .B(micro_hash_ucr_pipe12), .Y(_1621_) );
NAND3X1 NAND3X1_50 ( .gnd(gnd), .vdd(vdd), .A(_936_), .B(_965_), .C(_1621_), .Y(_1622_) );
OAI22X1 OAI22X1_34 ( .gnd(gnd), .vdd(vdd), .A(_955_), .B(_1622_), .C(_956_), .D(micro_hash_ucr_a_6_bF_buf1_), .Y(_1623_) );
NAND2X1 NAND2X1_203 ( .gnd(gnd), .vdd(vdd), .A(_935_), .B(_1623_), .Y(_1624_) );
OAI21X1 OAI21X1_434 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_6_bF_buf0_), .B(_931_), .C(_1624_), .Y(_1625_) );
NAND2X1 NAND2X1_204 ( .gnd(gnd), .vdd(vdd), .A(_933_), .B(_1625_), .Y(_1626_) );
NOR2X1 NOR2X1_321 ( .gnd(gnd), .vdd(vdd), .A(_1616_), .B(_1070_), .Y(_1627_) );
NOR2X1 NOR2X1_322 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe14_bF_buf2), .B(_1627_), .Y(_1628_) );
AOI22X1 AOI22X1_20 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_6_bF_buf3_), .B(micro_hash_ucr_pipe14_bF_buf1), .C(_1628_), .D(_1626_), .Y(_1629_) );
OAI21X1 OAI21X1_435 ( .gnd(gnd), .vdd(vdd), .A(_1629_), .B(micro_hash_ucr_pipe15_bF_buf3), .C(_1620_), .Y(_1630_) );
NAND2X1 NAND2X1_205 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe16_bF_buf3), .B(_494_), .Y(_1631_) );
OAI21X1 OAI21X1_436 ( .gnd(gnd), .vdd(vdd), .A(_1630_), .B(micro_hash_ucr_pipe16_bF_buf2), .C(_1631_), .Y(_1632_) );
OAI21X1 OAI21X1_437 ( .gnd(gnd), .vdd(vdd), .A(_1616_), .B(_929_), .C(_925__bF_buf4), .Y(_1633_) );
AOI21X1 AOI21X1_320 ( .gnd(gnd), .vdd(vdd), .A(_929_), .B(_1632_), .C(_1633_), .Y(_1634_) );
OAI21X1 OAI21X1_438 ( .gnd(gnd), .vdd(vdd), .A(_1634_), .B(_1619_), .C(_927__bF_buf0), .Y(_1635_) );
NAND2X1 NAND2X1_206 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe19_bF_buf3), .B(_1616_), .Y(_1636_) );
AOI21X1 AOI21X1_321 ( .gnd(gnd), .vdd(vdd), .A(_1636_), .B(_1635_), .C(micro_hash_ucr_pipe20_bF_buf1), .Y(_1637_) );
OAI21X1 OAI21X1_439 ( .gnd(gnd), .vdd(vdd), .A(_1637_), .B(_1618_), .C(_922_), .Y(_1638_) );
OAI21X1 OAI21X1_440 ( .gnd(gnd), .vdd(vdd), .A(_922_), .B(_1617_), .C(_1638_), .Y(_1639_) );
NAND2X1 NAND2X1_207 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf3), .B(_1639_), .Y(_1640_) );
OAI21X1 OAI21X1_441 ( .gnd(gnd), .vdd(vdd), .A(_494_), .B(_924__bF_buf2), .C(_1640_), .Y(_1641_) );
OAI21X1 OAI21X1_442 ( .gnd(gnd), .vdd(vdd), .A(_1615_), .B(_1614_), .C(micro_hash_ucr_pipe23_bF_buf3), .Y(_1642_) );
OAI21X1 OAI21X1_443 ( .gnd(gnd), .vdd(vdd), .A(_1641_), .B(micro_hash_ucr_pipe23_bF_buf2), .C(_1642_), .Y(_1643_) );
OAI21X1 OAI21X1_444 ( .gnd(gnd), .vdd(vdd), .A(_919__bF_buf3), .B(micro_hash_ucr_a_6_bF_buf2_), .C(_921__bF_buf1), .Y(_1644_) );
AOI21X1 AOI21X1_322 ( .gnd(gnd), .vdd(vdd), .A(_919__bF_buf2), .B(_1643_), .C(_1644_), .Y(_1645_) );
OAI21X1 OAI21X1_445 ( .gnd(gnd), .vdd(vdd), .A(_1617_), .B(_921__bF_buf0), .C(_920__bF_buf3), .Y(_1646_) );
OAI22X1 OAI22X1_35 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_6_bF_buf1_), .B(_920__bF_buf2), .C(_1645_), .D(_1646_), .Y(_1647_) );
NAND2X1 NAND2X1_208 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe27), .B(_1616_), .Y(_1648_) );
OAI21X1 OAI21X1_446 ( .gnd(gnd), .vdd(vdd), .A(_1647_), .B(micro_hash_ucr_pipe27), .C(_1648_), .Y(_1649_) );
NOR2X1 NOR2X1_323 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe28_bF_buf3), .B(_1649_), .Y(_1650_) );
OAI21X1 OAI21X1_447 ( .gnd(gnd), .vdd(vdd), .A(_918__bF_buf4), .B(micro_hash_ucr_a_6_bF_buf0_), .C(_917_), .Y(_1651_) );
AOI21X1 AOI21X1_323 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe29_bF_buf2), .B(_1616_), .C(micro_hash_ucr_pipe30_bF_buf0), .Y(_1652_) );
OAI21X1 OAI21X1_448 ( .gnd(gnd), .vdd(vdd), .A(_1650_), .B(_1651_), .C(_1652_), .Y(_1653_) );
NAND2X1 NAND2X1_209 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe30_bF_buf3), .B(_494_), .Y(_1654_) );
AOI21X1 AOI21X1_324 ( .gnd(gnd), .vdd(vdd), .A(_1654_), .B(_1653_), .C(micro_hash_ucr_pipe31), .Y(_1655_) );
NOR2X1 NOR2X1_324 ( .gnd(gnd), .vdd(vdd), .A(_915__bF_buf2), .B(_1616_), .Y(_1656_) );
OAI21X1 OAI21X1_449 ( .gnd(gnd), .vdd(vdd), .A(_1655_), .B(_1656_), .C(_914__bF_buf3), .Y(_1657_) );
NAND3X1 NAND3X1_51 ( .gnd(gnd), .vdd(vdd), .A(_910_), .B(_1613_), .C(_1657_), .Y(_1658_) );
AOI21X1 AOI21X1_325 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe33_bF_buf0), .B(_1616_), .C(micro_hash_ucr_pipe34_bF_buf0), .Y(_1659_) );
OAI21X1 OAI21X1_450 ( .gnd(gnd), .vdd(vdd), .A(_912__bF_buf2), .B(micro_hash_ucr_a_6_bF_buf3_), .C(_911__bF_buf4), .Y(_1660_) );
AOI21X1 AOI21X1_326 ( .gnd(gnd), .vdd(vdd), .A(_1659_), .B(_1658_), .C(_1660_), .Y(_1661_) );
OAI21X1 OAI21X1_451 ( .gnd(gnd), .vdd(vdd), .A(_1617_), .B(_911__bF_buf3), .C(_907__bF_buf2), .Y(_1662_) );
OAI22X1 OAI22X1_36 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_6_bF_buf2_), .B(_907__bF_buf1), .C(_1661_), .D(_1662_), .Y(_1663_) );
OAI21X1 OAI21X1_452 ( .gnd(gnd), .vdd(vdd), .A(_1616_), .B(_909__bF_buf3), .C(_908__bF_buf2), .Y(_1664_) );
AOI21X1 AOI21X1_327 ( .gnd(gnd), .vdd(vdd), .A(_909__bF_buf2), .B(_1663_), .C(_1664_), .Y(_1665_) );
NOR2X1 NOR2X1_325 ( .gnd(gnd), .vdd(vdd), .A(_494_), .B(_908__bF_buf1), .Y(_1666_) );
OAI21X1 OAI21X1_453 ( .gnd(gnd), .vdd(vdd), .A(_1665_), .B(_1666_), .C(_904__bF_buf1), .Y(_1667_) );
NAND2X1 NAND2X1_210 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe39), .B(_1616_), .Y(_1668_) );
AOI21X1 AOI21X1_328 ( .gnd(gnd), .vdd(vdd), .A(_1668_), .B(_1667_), .C(micro_hash_ucr_pipe40_bF_buf3), .Y(_1669_) );
OAI21X1 OAI21X1_454 ( .gnd(gnd), .vdd(vdd), .A(_494_), .B(_906__bF_buf1), .C(_905__bF_buf3), .Y(_1670_) );
AOI21X1 AOI21X1_329 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe41), .B(_1617_), .C(micro_hash_ucr_pipe42_bF_buf3), .Y(_1671_) );
OAI21X1 OAI21X1_455 ( .gnd(gnd), .vdd(vdd), .A(_1669_), .B(_1670_), .C(_1671_), .Y(_1672_) );
NAND2X1 NAND2X1_211 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_6_bF_buf1_), .B(micro_hash_ucr_pipe42_bF_buf2), .Y(_1673_) );
AOI21X1 AOI21X1_330 ( .gnd(gnd), .vdd(vdd), .A(_1673_), .B(_1672_), .C(micro_hash_ucr_pipe43), .Y(_1674_) );
NOR2X1 NOR2X1_326 ( .gnd(gnd), .vdd(vdd), .A(_903__bF_buf1), .B(_1617_), .Y(_1675_) );
OAI21X1 OAI21X1_456 ( .gnd(gnd), .vdd(vdd), .A(_1674_), .B(_1675_), .C(_902__bF_buf3), .Y(_1676_) );
AOI21X1 AOI21X1_331 ( .gnd(gnd), .vdd(vdd), .A(_1612_), .B(_1676_), .C(micro_hash_ucr_pipe45_bF_buf0), .Y(_1677_) );
NOR2X1 NOR2X1_327 ( .gnd(gnd), .vdd(vdd), .A(_898_), .B(_1617_), .Y(_1678_) );
OAI21X1 OAI21X1_457 ( .gnd(gnd), .vdd(vdd), .A(_1677_), .B(_1678_), .C(_900__bF_buf1), .Y(_1679_) );
NAND3X1 NAND3X1_52 ( .gnd(gnd), .vdd(vdd), .A(_899__bF_buf0), .B(_1611_), .C(_1679_), .Y(_1680_) );
OAI21X1 OAI21X1_458 ( .gnd(gnd), .vdd(vdd), .A(_1615_), .B(_1614_), .C(micro_hash_ucr_pipe47), .Y(_1681_) );
NAND3X1 NAND3X1_53 ( .gnd(gnd), .vdd(vdd), .A(_895__bF_buf2), .B(_1681_), .C(_1680_), .Y(_1682_) );
NAND3X1 NAND3X1_54 ( .gnd(gnd), .vdd(vdd), .A(_897__bF_buf3), .B(_1610_), .C(_1682_), .Y(_1683_) );
OAI21X1 OAI21X1_459 ( .gnd(gnd), .vdd(vdd), .A(_1615_), .B(_1614_), .C(micro_hash_ucr_pipe49), .Y(_1684_) );
NAND3X1 NAND3X1_55 ( .gnd(gnd), .vdd(vdd), .A(_896__bF_buf2), .B(_1684_), .C(_1683_), .Y(_1685_) );
NAND3X1 NAND3X1_56 ( .gnd(gnd), .vdd(vdd), .A(_892_), .B(_1609_), .C(_1685_), .Y(_1686_) );
OAI21X1 OAI21X1_460 ( .gnd(gnd), .vdd(vdd), .A(_1615_), .B(_1614_), .C(micro_hash_ucr_pipe51), .Y(_1687_) );
NAND3X1 NAND3X1_57 ( .gnd(gnd), .vdd(vdd), .A(_894__bF_buf3), .B(_1687_), .C(_1686_), .Y(_1688_) );
AOI21X1 AOI21X1_332 ( .gnd(gnd), .vdd(vdd), .A(_1608_), .B(_1688_), .C(micro_hash_ucr_pipe53_bF_buf0), .Y(_1689_) );
OAI21X1 OAI21X1_461 ( .gnd(gnd), .vdd(vdd), .A(_1617_), .B(_893_), .C(_889__bF_buf2), .Y(_1690_) );
AOI21X1 AOI21X1_333 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe54_bF_buf0), .B(_494_), .C(micro_hash_ucr_pipe55), .Y(_1691_) );
OAI21X1 OAI21X1_462 ( .gnd(gnd), .vdd(vdd), .A(_1689_), .B(_1690_), .C(_1691_), .Y(_1692_) );
AOI21X1 AOI21X1_334 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe55), .B(_1616_), .C(micro_hash_ucr_pipe56_bF_buf2), .Y(_1693_) );
NAND2X1 NAND2X1_212 ( .gnd(gnd), .vdd(vdd), .A(_1693_), .B(_1692_), .Y(_1694_) );
NAND2X1 NAND2X1_213 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe56_bF_buf1), .B(_494_), .Y(_1695_) );
NAND3X1 NAND3X1_58 ( .gnd(gnd), .vdd(vdd), .A(_886_), .B(_1695_), .C(_1694_), .Y(_1696_) );
NAND2X1 NAND2X1_214 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe57_bF_buf1), .B(_1616_), .Y(_1697_) );
AOI21X1 AOI21X1_335 ( .gnd(gnd), .vdd(vdd), .A(_1697_), .B(_1696_), .C(micro_hash_ucr_pipe58_bF_buf0), .Y(_1698_) );
OAI21X1 OAI21X1_463 ( .gnd(gnd), .vdd(vdd), .A(_494_), .B(_888__bF_buf2), .C(_887__bF_buf0), .Y(_1699_) );
AOI21X1 AOI21X1_336 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe59), .B(_1617_), .C(micro_hash_ucr_pipe60_bF_buf2), .Y(_1700_) );
OAI21X1 OAI21X1_464 ( .gnd(gnd), .vdd(vdd), .A(_1698_), .B(_1699_), .C(_1700_), .Y(_1701_) );
NAND2X1 NAND2X1_215 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_6_bF_buf0_), .B(micro_hash_ucr_pipe60_bF_buf1), .Y(_1702_) );
NAND3X1 NAND3X1_59 ( .gnd(gnd), .vdd(vdd), .A(_885_), .B(_1702_), .C(_1701_), .Y(_1703_) );
OAI21X1 OAI21X1_465 ( .gnd(gnd), .vdd(vdd), .A(_1615_), .B(_1614_), .C(micro_hash_ucr_pipe61_bF_buf0), .Y(_1704_) );
NAND3X1 NAND3X1_60 ( .gnd(gnd), .vdd(vdd), .A(_884__bF_buf1), .B(_1704_), .C(_1703_), .Y(_1705_) );
NAND3X1 NAND3X1_61 ( .gnd(gnd), .vdd(vdd), .A(_880__bF_buf2), .B(_1607_), .C(_1705_), .Y(_1706_) );
OAI21X1 OAI21X1_466 ( .gnd(gnd), .vdd(vdd), .A(_1615_), .B(_1614_), .C(micro_hash_ucr_pipe63), .Y(_1707_) );
NAND3X1 NAND3X1_62 ( .gnd(gnd), .vdd(vdd), .A(_882__bF_buf2), .B(_1707_), .C(_1706_), .Y(_1708_) );
NAND3X1 NAND3X1_63 ( .gnd(gnd), .vdd(vdd), .A(_881_), .B(_1606_), .C(_1708_), .Y(_1709_) );
OAI21X1 OAI21X1_467 ( .gnd(gnd), .vdd(vdd), .A(_1615_), .B(_1614_), .C(micro_hash_ucr_pipe65_bF_buf2), .Y(_1710_) );
NAND3X1 NAND3X1_64 ( .gnd(gnd), .vdd(vdd), .A(_877__bF_buf0), .B(_1710_), .C(_1709_), .Y(_1711_) );
NAND3X1 NAND3X1_65 ( .gnd(gnd), .vdd(vdd), .A(_879__bF_buf2), .B(_1605_), .C(_1711_), .Y(_1712_) );
OAI21X1 OAI21X1_468 ( .gnd(gnd), .vdd(vdd), .A(_1615_), .B(_1614_), .C(micro_hash_ucr_pipe67), .Y(_1713_) );
NAND3X1 NAND3X1_66 ( .gnd(gnd), .vdd(vdd), .A(_878__bF_buf1), .B(_1713_), .C(_1712_), .Y(_1714_) );
AOI21X1 AOI21X1_337 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_6_bF_buf3_), .B(micro_hash_ucr_pipe68), .C(micro_hash_ucr_pipe69), .Y(_1715_) );
OAI21X1 OAI21X1_469 ( .gnd(gnd), .vdd(vdd), .A(_1616_), .B(_876__bF_buf1), .C(_302__bF_buf8), .Y(_1716_) );
AOI21X1 AOI21X1_338 ( .gnd(gnd), .vdd(vdd), .A(_1715_), .B(_1714_), .C(_1716_), .Y(_297__6_) );
INVX8 INVX8_84 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_7_), .Y(_1717_) );
NAND2X1 NAND2X1_216 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe62_bF_buf2), .B(_1717__bF_buf3), .Y(_1718_) );
NAND2X1 NAND2X1_217 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe60_bF_buf0), .B(_1717__bF_buf2), .Y(_1719_) );
INVX1 INVX1_104 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_7_), .Y(_1720_) );
INVX8 INVX8_85 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_7_), .Y(_1721_) );
NAND2X1 NAND2X1_218 ( .gnd(gnd), .vdd(vdd), .A(_1720_), .B(_1721__bF_buf4), .Y(_1722_) );
NAND2X1 NAND2X1_219 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_7_), .B(micro_hash_ucr_b_7_), .Y(_1723_) );
NAND2X1 NAND2X1_220 ( .gnd(gnd), .vdd(vdd), .A(_1723_), .B(_1722_), .Y(_1724_) );
INVX8 INVX8_86 ( .gnd(gnd), .vdd(vdd), .A(_1724_), .Y(_1725_) );
NAND2X1 NAND2X1_221 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe44), .B(_1717__bF_buf1), .Y(_1726_) );
NOR2X1 NOR2X1_328 ( .gnd(gnd), .vdd(vdd), .A(_1717__bF_buf0), .B(_901__bF_buf4), .Y(_1727_) );
NOR2X1 NOR2X1_329 ( .gnd(gnd), .vdd(vdd), .A(_1717__bF_buf3), .B(_906__bF_buf0), .Y(_1728_) );
NOR2X1 NOR2X1_330 ( .gnd(gnd), .vdd(vdd), .A(_1717__bF_buf2), .B(_908__bF_buf0), .Y(_1729_) );
NOR2X1 NOR2X1_331 ( .gnd(gnd), .vdd(vdd), .A(_1717__bF_buf1), .B(_907__bF_buf0), .Y(_1730_) );
NOR2X1 NOR2X1_332 ( .gnd(gnd), .vdd(vdd), .A(_1717__bF_buf0), .B(_912__bF_buf1), .Y(_1731_) );
NOR2X1 NOR2X1_333 ( .gnd(gnd), .vdd(vdd), .A(_1717__bF_buf3), .B(_918__bF_buf3), .Y(_1732_) );
NAND2X1 NAND2X1_222 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe17_bF_buf2), .B(_1725__bF_buf3), .Y(_1733_) );
NAND2X1 NAND2X1_223 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe15_bF_buf2), .B(_1725__bF_buf2), .Y(_1734_) );
NAND2X1 NAND2X1_224 ( .gnd(gnd), .vdd(vdd), .A(_1717__bF_buf2), .B(_957_), .Y(_1735_) );
NAND3X1 NAND3X1_67 ( .gnd(gnd), .vdd(vdd), .A(_500_), .B(_939_), .C(_1187_), .Y(_1736_) );
OAI21X1 OAI21X1_470 ( .gnd(gnd), .vdd(vdd), .A(_1186_), .B(_1736_), .C(_1735_), .Y(_1737_) );
NAND2X1 NAND2X1_225 ( .gnd(gnd), .vdd(vdd), .A(_933_), .B(_1737_), .Y(_1738_) );
NOR2X1 NOR2X1_334 ( .gnd(gnd), .vdd(vdd), .A(_1725__bF_buf1), .B(_1070_), .Y(_1739_) );
NOR2X1 NOR2X1_335 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe14_bF_buf0), .B(_1739_), .Y(_1740_) );
AOI22X1 AOI22X1_21 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_7_), .B(micro_hash_ucr_pipe14_bF_buf4), .C(_1740_), .D(_1738_), .Y(_1741_) );
OAI21X1 OAI21X1_471 ( .gnd(gnd), .vdd(vdd), .A(_1741_), .B(micro_hash_ucr_pipe15_bF_buf1), .C(_1734_), .Y(_1742_) );
NAND2X1 NAND2X1_226 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe16_bF_buf1), .B(_1717__bF_buf1), .Y(_1743_) );
OAI21X1 OAI21X1_472 ( .gnd(gnd), .vdd(vdd), .A(_1742_), .B(micro_hash_ucr_pipe16_bF_buf0), .C(_1743_), .Y(_1744_) );
OAI21X1 OAI21X1_473 ( .gnd(gnd), .vdd(vdd), .A(_1744_), .B(micro_hash_ucr_pipe17_bF_buf1), .C(_1733_), .Y(_1745_) );
OAI21X1 OAI21X1_474 ( .gnd(gnd), .vdd(vdd), .A(_1717__bF_buf0), .B(_925__bF_buf3), .C(_927__bF_buf3), .Y(_1746_) );
AOI21X1 AOI21X1_339 ( .gnd(gnd), .vdd(vdd), .A(_925__bF_buf2), .B(_1745_), .C(_1746_), .Y(_1747_) );
OAI21X1 OAI21X1_475 ( .gnd(gnd), .vdd(vdd), .A(_1725__bF_buf0), .B(_927__bF_buf2), .C(_926__bF_buf1), .Y(_1748_) );
NOR2X1 NOR2X1_336 ( .gnd(gnd), .vdd(vdd), .A(_1748_), .B(_1747_), .Y(_1749_) );
NOR2X1 NOR2X1_337 ( .gnd(gnd), .vdd(vdd), .A(_1717__bF_buf3), .B(_926__bF_buf0), .Y(_1750_) );
OAI21X1 OAI21X1_476 ( .gnd(gnd), .vdd(vdd), .A(_1749_), .B(_1750_), .C(_922_), .Y(_1751_) );
AOI21X1 AOI21X1_340 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe21_bF_buf3), .B(_1725__bF_buf3), .C(micro_hash_ucr_pipe22_bF_buf0), .Y(_1752_) );
OAI21X1 OAI21X1_477 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf1), .B(micro_hash_ucr_a_7_), .C(_923_), .Y(_1753_) );
AOI21X1 AOI21X1_341 ( .gnd(gnd), .vdd(vdd), .A(_1752_), .B(_1751_), .C(_1753_), .Y(_1754_) );
OAI21X1 OAI21X1_478 ( .gnd(gnd), .vdd(vdd), .A(_1724_), .B(_923_), .C(_919__bF_buf1), .Y(_1755_) );
OAI22X1 OAI22X1_37 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_7_), .B(_919__bF_buf0), .C(_1754_), .D(_1755_), .Y(_1756_) );
OAI21X1 OAI21X1_479 ( .gnd(gnd), .vdd(vdd), .A(_1725__bF_buf2), .B(_921__bF_buf3), .C(_920__bF_buf1), .Y(_1757_) );
AOI21X1 AOI21X1_342 ( .gnd(gnd), .vdd(vdd), .A(_921__bF_buf2), .B(_1756_), .C(_1757_), .Y(_1758_) );
NOR2X1 NOR2X1_338 ( .gnd(gnd), .vdd(vdd), .A(_1717__bF_buf2), .B(_920__bF_buf0), .Y(_1759_) );
OAI21X1 OAI21X1_480 ( .gnd(gnd), .vdd(vdd), .A(_1758_), .B(_1759_), .C(_916_), .Y(_1760_) );
NAND2X1 NAND2X1_227 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe27), .B(_1725__bF_buf1), .Y(_1761_) );
AOI21X1 AOI21X1_343 ( .gnd(gnd), .vdd(vdd), .A(_1761_), .B(_1760_), .C(micro_hash_ucr_pipe28_bF_buf2), .Y(_1762_) );
OAI21X1 OAI21X1_481 ( .gnd(gnd), .vdd(vdd), .A(_1762_), .B(_1732_), .C(_917_), .Y(_1763_) );
OAI21X1 OAI21X1_482 ( .gnd(gnd), .vdd(vdd), .A(_917_), .B(_1724_), .C(_1763_), .Y(_1764_) );
NOR2X1 NOR2X1_339 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe30_bF_buf2), .B(_1764_), .Y(_1765_) );
OAI21X1 OAI21X1_483 ( .gnd(gnd), .vdd(vdd), .A(_913__bF_buf2), .B(micro_hash_ucr_a_7_), .C(_915__bF_buf1), .Y(_1766_) );
AOI21X1 AOI21X1_344 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe31), .B(_1725__bF_buf0), .C(micro_hash_ucr_pipe32_bF_buf3), .Y(_1767_) );
OAI21X1 OAI21X1_484 ( .gnd(gnd), .vdd(vdd), .A(_1765_), .B(_1766_), .C(_1767_), .Y(_1768_) );
OAI21X1 OAI21X1_485 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_7_), .B(_914__bF_buf2), .C(_1768_), .Y(_1769_) );
NAND2X1 NAND2X1_228 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe33_bF_buf3), .B(_1725__bF_buf3), .Y(_1770_) );
OAI21X1 OAI21X1_486 ( .gnd(gnd), .vdd(vdd), .A(_1769_), .B(micro_hash_ucr_pipe33_bF_buf2), .C(_1770_), .Y(_1771_) );
AND2X2 AND2X2_190 ( .gnd(gnd), .vdd(vdd), .A(_1771_), .B(_912__bF_buf0), .Y(_1772_) );
OAI21X1 OAI21X1_487 ( .gnd(gnd), .vdd(vdd), .A(_1772_), .B(_1731_), .C(_911__bF_buf2), .Y(_1773_) );
NAND2X1 NAND2X1_229 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe35), .B(_1725__bF_buf2), .Y(_1774_) );
AOI21X1 AOI21X1_345 ( .gnd(gnd), .vdd(vdd), .A(_1774_), .B(_1773_), .C(micro_hash_ucr_pipe36_bF_buf0), .Y(_1775_) );
OAI21X1 OAI21X1_488 ( .gnd(gnd), .vdd(vdd), .A(_1775_), .B(_1730_), .C(_909__bF_buf1), .Y(_1776_) );
NAND2X1 NAND2X1_230 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe37), .B(_1725__bF_buf1), .Y(_1777_) );
AOI21X1 AOI21X1_346 ( .gnd(gnd), .vdd(vdd), .A(_1777_), .B(_1776_), .C(micro_hash_ucr_pipe38_bF_buf0), .Y(_1778_) );
OAI21X1 OAI21X1_489 ( .gnd(gnd), .vdd(vdd), .A(_1778_), .B(_1729_), .C(_904__bF_buf0), .Y(_1779_) );
NAND2X1 NAND2X1_231 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe39), .B(_1725__bF_buf0), .Y(_1780_) );
AOI21X1 AOI21X1_347 ( .gnd(gnd), .vdd(vdd), .A(_1780_), .B(_1779_), .C(micro_hash_ucr_pipe40_bF_buf2), .Y(_1781_) );
OAI21X1 OAI21X1_490 ( .gnd(gnd), .vdd(vdd), .A(_1781_), .B(_1728_), .C(_905__bF_buf2), .Y(_1782_) );
NAND2X1 NAND2X1_232 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe41), .B(_1725__bF_buf3), .Y(_1783_) );
AOI21X1 AOI21X1_348 ( .gnd(gnd), .vdd(vdd), .A(_1783_), .B(_1782_), .C(micro_hash_ucr_pipe42_bF_buf1), .Y(_1784_) );
OAI21X1 OAI21X1_491 ( .gnd(gnd), .vdd(vdd), .A(_1784_), .B(_1727_), .C(_903__bF_buf0), .Y(_1785_) );
NAND2X1 NAND2X1_233 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe43), .B(_1725__bF_buf2), .Y(_1786_) );
NAND3X1 NAND3X1_68 ( .gnd(gnd), .vdd(vdd), .A(_902__bF_buf2), .B(_1786_), .C(_1785_), .Y(_1787_) );
NAND3X1 NAND3X1_69 ( .gnd(gnd), .vdd(vdd), .A(_898_), .B(_1726_), .C(_1787_), .Y(_1788_) );
AOI21X1 AOI21X1_349 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe45_bF_buf3), .B(_1725__bF_buf1), .C(micro_hash_ucr_pipe46_bF_buf0), .Y(_1789_) );
OAI21X1 OAI21X1_492 ( .gnd(gnd), .vdd(vdd), .A(_900__bF_buf0), .B(micro_hash_ucr_a_7_), .C(_899__bF_buf3), .Y(_1790_) );
AOI21X1 AOI21X1_350 ( .gnd(gnd), .vdd(vdd), .A(_1789_), .B(_1788_), .C(_1790_), .Y(_1791_) );
OAI21X1 OAI21X1_493 ( .gnd(gnd), .vdd(vdd), .A(_1724_), .B(_899__bF_buf2), .C(_895__bF_buf1), .Y(_1792_) );
OAI22X1 OAI22X1_38 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_7_), .B(_895__bF_buf0), .C(_1791_), .D(_1792_), .Y(_1793_) );
NAND2X1 NAND2X1_234 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe49), .B(_1725__bF_buf0), .Y(_1794_) );
OAI21X1 OAI21X1_494 ( .gnd(gnd), .vdd(vdd), .A(_1793_), .B(micro_hash_ucr_pipe49), .C(_1794_), .Y(_1795_) );
NAND2X1 NAND2X1_235 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe50_bF_buf3), .B(_1717__bF_buf1), .Y(_1796_) );
OAI21X1 OAI21X1_495 ( .gnd(gnd), .vdd(vdd), .A(_1795_), .B(micro_hash_ucr_pipe50_bF_buf2), .C(_1796_), .Y(_1797_) );
AOI21X1 AOI21X1_351 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe51), .B(_1725__bF_buf3), .C(micro_hash_ucr_pipe52_bF_buf2), .Y(_1798_) );
OAI21X1 OAI21X1_496 ( .gnd(gnd), .vdd(vdd), .A(_1797_), .B(micro_hash_ucr_pipe51), .C(_1798_), .Y(_1799_) );
AOI21X1 AOI21X1_352 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe52_bF_buf1), .B(_1717__bF_buf0), .C(micro_hash_ucr_pipe53_bF_buf3), .Y(_1800_) );
AOI22X1 AOI22X1_22 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe53_bF_buf2), .B(_1725__bF_buf2), .C(_1799_), .D(_1800_), .Y(_1801_) );
AOI21X1 AOI21X1_353 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_7_), .B(micro_hash_ucr_pipe54_bF_buf3), .C(micro_hash_ucr_pipe55), .Y(_1802_) );
OAI21X1 OAI21X1_497 ( .gnd(gnd), .vdd(vdd), .A(_1801_), .B(micro_hash_ucr_pipe54_bF_buf2), .C(_1802_), .Y(_1803_) );
NAND2X1 NAND2X1_236 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe55), .B(_1724_), .Y(_1804_) );
AOI21X1 AOI21X1_354 ( .gnd(gnd), .vdd(vdd), .A(_1804_), .B(_1803_), .C(micro_hash_ucr_pipe56_bF_buf0), .Y(_1805_) );
OAI21X1 OAI21X1_498 ( .gnd(gnd), .vdd(vdd), .A(_890__bF_buf0), .B(micro_hash_ucr_a_7_), .C(_886_), .Y(_1806_) );
AOI21X1 AOI21X1_355 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe57_bF_buf0), .B(_1725__bF_buf1), .C(micro_hash_ucr_pipe58_bF_buf4), .Y(_1807_) );
OAI21X1 OAI21X1_499 ( .gnd(gnd), .vdd(vdd), .A(_1805_), .B(_1806_), .C(_1807_), .Y(_1808_) );
NAND2X1 NAND2X1_237 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe58_bF_buf3), .B(_1717__bF_buf3), .Y(_1809_) );
NAND3X1 NAND3X1_70 ( .gnd(gnd), .vdd(vdd), .A(_887__bF_buf3), .B(_1809_), .C(_1808_), .Y(_1810_) );
NAND2X1 NAND2X1_238 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe59), .B(_1725__bF_buf0), .Y(_1811_) );
NAND3X1 NAND3X1_71 ( .gnd(gnd), .vdd(vdd), .A(_883__bF_buf0), .B(_1811_), .C(_1810_), .Y(_1812_) );
NAND3X1 NAND3X1_72 ( .gnd(gnd), .vdd(vdd), .A(_885_), .B(_1719_), .C(_1812_), .Y(_1813_) );
NAND2X1 NAND2X1_239 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe61_bF_buf3), .B(_1725__bF_buf3), .Y(_1814_) );
NAND3X1 NAND3X1_73 ( .gnd(gnd), .vdd(vdd), .A(_884__bF_buf0), .B(_1814_), .C(_1813_), .Y(_1815_) );
NAND3X1 NAND3X1_74 ( .gnd(gnd), .vdd(vdd), .A(_880__bF_buf1), .B(_1718_), .C(_1815_), .Y(_1816_) );
NAND2X1 NAND2X1_240 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe63), .B(_1725__bF_buf2), .Y(_1817_) );
AOI21X1 AOI21X1_356 ( .gnd(gnd), .vdd(vdd), .A(_1817_), .B(_1816_), .C(micro_hash_ucr_pipe64_bF_buf3), .Y(_1818_) );
OAI21X1 OAI21X1_500 ( .gnd(gnd), .vdd(vdd), .A(_1717__bF_buf2), .B(_882__bF_buf1), .C(_881_), .Y(_1819_) );
AOI21X1 AOI21X1_357 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe65_bF_buf1), .B(_1724_), .C(micro_hash_ucr_pipe66_bF_buf1), .Y(_1820_) );
OAI21X1 OAI21X1_501 ( .gnd(gnd), .vdd(vdd), .A(_1818_), .B(_1819_), .C(_1820_), .Y(_1821_) );
NAND2X1 NAND2X1_241 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_7_), .B(micro_hash_ucr_pipe66_bF_buf0), .Y(_1822_) );
NAND3X1 NAND3X1_75 ( .gnd(gnd), .vdd(vdd), .A(_879__bF_buf1), .B(_1822_), .C(_1821_), .Y(_1823_) );
NAND2X1 NAND2X1_242 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe67), .B(_1724_), .Y(_1824_) );
NAND3X1 NAND3X1_76 ( .gnd(gnd), .vdd(vdd), .A(_878__bF_buf0), .B(_1824_), .C(_1823_), .Y(_1825_) );
AOI21X1 AOI21X1_358 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_a_7_), .B(micro_hash_ucr_pipe68), .C(micro_hash_ucr_pipe69), .Y(_1826_) );
OAI21X1 OAI21X1_502 ( .gnd(gnd), .vdd(vdd), .A(_1725__bF_buf1), .B(_876__bF_buf0), .C(_302__bF_buf7), .Y(_1827_) );
AOI21X1 AOI21X1_359 ( .gnd(gnd), .vdd(vdd), .A(_1826_), .B(_1825_), .C(_1827_), .Y(_297__7_) );
INVX1 INVX1_105 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_k_0_), .Y(_1828_) );
NOR2X1 NOR2X1_340 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe40_bF_buf1), .B(micro_hash_ucr_pipe7), .Y(_1829_) );
AOI21X1 AOI21X1_360 ( .gnd(gnd), .vdd(vdd), .A(_1828_), .B(_1829_), .C(_400__bF_buf5), .Y(_301__0_) );
NAND2X1 NAND2X1_243 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_k_1_), .B(_1829_), .Y(_1830_) );
NOR2X1 NOR2X1_341 ( .gnd(gnd), .vdd(vdd), .A(_1830_), .B(_400__bF_buf4), .Y(_301__1_) );
NAND2X1 NAND2X1_244 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_k_2_), .B(_1829_), .Y(_1831_) );
NOR2X1 NOR2X1_342 ( .gnd(gnd), .vdd(vdd), .A(_1831_), .B(_400__bF_buf3), .Y(_301__2_) );
OAI21X1 OAI21X1_503 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe7), .B(micro_hash_ucr_k_3_), .C(_906__bF_buf4), .Y(_1832_) );
NOR2X1 NOR2X1_343 ( .gnd(gnd), .vdd(vdd), .A(_1832_), .B(_400__bF_buf2), .Y(_301__3_) );
OAI21X1 OAI21X1_504 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe7), .B(micro_hash_ucr_k_4_), .C(_906__bF_buf3), .Y(_1833_) );
NOR2X1 NOR2X1_344 ( .gnd(gnd), .vdd(vdd), .A(_1833_), .B(_400__bF_buf1), .Y(_301__4_) );
INVX2 INVX2_94 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_k_5_), .Y(_1834_) );
OAI21X1 OAI21X1_505 ( .gnd(gnd), .vdd(vdd), .A(_1834_), .B(micro_hash_ucr_pipe7), .C(_906__bF_buf2), .Y(_1835_) );
AND2X2 AND2X2_191 ( .gnd(gnd), .vdd(vdd), .A(_302__bF_buf6), .B(_1835_), .Y(_301__5_) );
NAND2X1 NAND2X1_245 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_k_6_), .B(_1829_), .Y(_1836_) );
NOR2X1 NOR2X1_345 ( .gnd(gnd), .vdd(vdd), .A(_1836_), .B(_400__bF_buf0), .Y(_301__6_) );
INVX1 INVX1_106 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_k_7_), .Y(_1837_) );
AOI21X1 AOI21X1_361 ( .gnd(gnd), .vdd(vdd), .A(_1837_), .B(_1829_), .C(_400__bF_buf12), .Y(_301__7_) );
NAND2X1 NAND2X1_246 ( .gnd(gnd), .vdd(vdd), .A(_4481_), .B(_436_), .Y(_1838_) );
NOR2X1 NOR2X1_346 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe21_bF_buf2), .B(micro_hash_ucr_pipe23_bF_buf1), .Y(_1839_) );
INVX1 INVX1_107 ( .gnd(gnd), .vdd(vdd), .A(_1839_), .Y(_1840_) );
NOR2X1 NOR2X1_347 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe39), .B(micro_hash_ucr_pipe37), .Y(_1841_) );
INVX1 INVX1_108 ( .gnd(gnd), .vdd(vdd), .A(_1841_), .Y(_1842_) );
NOR2X1 NOR2X1_348 ( .gnd(gnd), .vdd(vdd), .A(_1840_), .B(_1842_), .Y(_1843_) );
NOR2X1 NOR2X1_349 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe27), .B(micro_hash_ucr_pipe29_bF_buf1), .Y(_1844_) );
AND2X2 AND2X2_192 ( .gnd(gnd), .vdd(vdd), .A(_1844_), .B(_911__bF_buf1), .Y(_1845_) );
AND2X2 AND2X2_193 ( .gnd(gnd), .vdd(vdd), .A(_1843_), .B(_1845_), .Y(_1846_) );
NAND3X1 NAND3X1_77 ( .gnd(gnd), .vdd(vdd), .A(_910_), .B(_915__bF_buf0), .C(_971_), .Y(_1847_) );
NOR2X1 NOR2X1_350 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe25), .B(micro_hash_ucr_pipe19_bF_buf2), .Y(_1848_) );
NAND2X1 NAND2X1_247 ( .gnd(gnd), .vdd(vdd), .A(_965_), .B(_1296_), .Y(_1849_) );
INVX1 INVX1_109 ( .gnd(gnd), .vdd(vdd), .A(_1849_), .Y(_1850_) );
NAND2X1 NAND2X1_248 ( .gnd(gnd), .vdd(vdd), .A(_1848_), .B(_1850_), .Y(_1851_) );
NOR2X1 NOR2X1_351 ( .gnd(gnd), .vdd(vdd), .A(_1847_), .B(_1851_), .Y(_1852_) );
NAND2X1 NAND2X1_249 ( .gnd(gnd), .vdd(vdd), .A(_1846_), .B(_1852_), .Y(_1853_) );
INVX4 INVX4_53 ( .gnd(gnd), .vdd(vdd), .A(_1853_), .Y(_1854_) );
AOI21X1 AOI21X1_362 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_0_bF_buf0_), .B(micro_hash_ucr_a_0_bF_buf0_), .C(_1854_), .Y(_1855_) );
NOR2X1 NOR2X1_352 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe45_bF_buf2), .B(micro_hash_ucr_pipe47), .Y(_1856_) );
NAND3X1 NAND3X1_78 ( .gnd(gnd), .vdd(vdd), .A(_903__bF_buf3), .B(_905__bF_buf1), .C(_1856_), .Y(_1857_) );
NOR2X1 NOR2X1_353 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe55), .B(micro_hash_ucr_pipe51), .Y(_1858_) );
NAND3X1 NAND3X1_79 ( .gnd(gnd), .vdd(vdd), .A(_893_), .B(_897__bF_buf2), .C(_1858_), .Y(_1859_) );
NOR2X1 NOR2X1_354 ( .gnd(gnd), .vdd(vdd), .A(_1857_), .B(_1859_), .Y(_1860_) );
NOR2X1 NOR2X1_355 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe67), .B(micro_hash_ucr_pipe65_bF_buf0), .Y(_1861_) );
INVX2 INVX2_95 ( .gnd(gnd), .vdd(vdd), .A(_1861_), .Y(_1862_) );
NOR2X1 NOR2X1_356 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe63), .B(micro_hash_ucr_pipe61_bF_buf2), .Y(_1863_) );
NAND3X1 NAND3X1_80 ( .gnd(gnd), .vdd(vdd), .A(_886_), .B(_887__bF_buf2), .C(_1863_), .Y(_1864_) );
NOR2X1 NOR2X1_357 ( .gnd(gnd), .vdd(vdd), .A(_1862_), .B(_1864_), .Y(_1865_) );
NAND2X1 NAND2X1_250 ( .gnd(gnd), .vdd(vdd), .A(_1865_), .B(_1860_), .Y(_1866_) );
OAI21X1 OAI21X1_506 ( .gnd(gnd), .vdd(vdd), .A(_1855_), .B(_1866_), .C(_1838_), .Y(_1867_) );
INVX2 INVX2_96 ( .gnd(gnd), .vdd(vdd), .A(_1860_), .Y(_1868_) );
NOR2X1 NOR2X1_358 ( .gnd(gnd), .vdd(vdd), .A(_1864_), .B(_1868_), .Y(_1869_) );
NOR2X1 NOR2X1_359 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe19_bF_buf1), .B(_1840_), .Y(_1870_) );
NAND3X1 NAND3X1_81 ( .gnd(gnd), .vdd(vdd), .A(_910_), .B(micro_hash_ucr_x_0_), .C(_965_), .Y(_1871_) );
NOR2X1 NOR2X1_360 ( .gnd(gnd), .vdd(vdd), .A(_1862_), .B(_1871_), .Y(_1872_) );
NAND2X1 NAND2X1_251 ( .gnd(gnd), .vdd(vdd), .A(_1870_), .B(_1872_), .Y(_1873_) );
NOR2X1 NOR2X1_361 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe31), .B(micro_hash_ucr_pipe29_bF_buf0), .Y(_1874_) );
NAND3X1 NAND3X1_82 ( .gnd(gnd), .vdd(vdd), .A(_971_), .B(_1296_), .C(_1874_), .Y(_1875_) );
NOR2X1 NOR2X1_362 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe27), .B(micro_hash_ucr_pipe25), .Y(_1876_) );
NAND3X1 NAND3X1_83 ( .gnd(gnd), .vdd(vdd), .A(_911__bF_buf0), .B(_1841_), .C(_1876_), .Y(_1877_) );
OR2X2 OR2X2_28 ( .gnd(gnd), .vdd(vdd), .A(_1875_), .B(_1877_), .Y(_1878_) );
NOR2X1 NOR2X1_363 ( .gnd(gnd), .vdd(vdd), .A(_1878_), .B(_1873_), .Y(_1879_) );
AOI21X1 AOI21X1_363 ( .gnd(gnd), .vdd(vdd), .A(_1869_), .B(_1879_), .C(micro_hash_ucr_pipe69), .Y(_1880_) );
OAI21X1 OAI21X1_507 ( .gnd(gnd), .vdd(vdd), .A(_876__bF_buf3), .B(_1838_), .C(_302__bF_buf5), .Y(_1881_) );
AOI21X1 AOI21X1_364 ( .gnd(gnd), .vdd(vdd), .A(_1880_), .B(_1867_), .C(_1881_), .Y(_375__0_) );
NAND2X1 NAND2X1_252 ( .gnd(gnd), .vdd(vdd), .A(_4487_), .B(_442_), .Y(_1882_) );
AOI21X1 AOI21X1_365 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_1_bF_buf0_), .B(micro_hash_ucr_a_1_), .C(_1854_), .Y(_1883_) );
OAI21X1 OAI21X1_508 ( .gnd(gnd), .vdd(vdd), .A(_1883_), .B(_1866_), .C(_1882_), .Y(_1884_) );
INVX1 INVX1_110 ( .gnd(gnd), .vdd(vdd), .A(_1869_), .Y(_1885_) );
NAND2X1 NAND2X1_253 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_x_1_), .B(_1861_), .Y(_1886_) );
NOR2X1 NOR2X1_364 ( .gnd(gnd), .vdd(vdd), .A(_1886_), .B(_1885_), .Y(_1887_) );
AOI21X1 AOI21X1_366 ( .gnd(gnd), .vdd(vdd), .A(_1854_), .B(_1887_), .C(micro_hash_ucr_pipe69), .Y(_1888_) );
OAI21X1 OAI21X1_509 ( .gnd(gnd), .vdd(vdd), .A(_876__bF_buf2), .B(_1882_), .C(_302__bF_buf4), .Y(_1889_) );
AOI21X1 AOI21X1_367 ( .gnd(gnd), .vdd(vdd), .A(_1888_), .B(_1884_), .C(_1889_), .Y(_375__1_) );
AOI21X1 AOI21X1_368 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_2_bF_buf0_), .B(micro_hash_ucr_a_2_), .C(_1854_), .Y(_1890_) );
NOR2X1 NOR2X1_365 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe69), .B(_1862_), .Y(_1891_) );
NAND2X1 NAND2X1_254 ( .gnd(gnd), .vdd(vdd), .A(_1891_), .B(_1869_), .Y(_1892_) );
OAI22X1 OAI22X1_39 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_2_bF_buf3_), .B(micro_hash_ucr_a_2_), .C(_1890_), .D(_1892_), .Y(_1893_) );
NAND3X1 NAND3X1_84 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_x_2_), .B(_1839_), .C(_1844_), .Y(_1894_) );
NOR2X1 NOR2X1_366 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe35), .B(_1842_), .Y(_1895_) );
NAND2X1 NAND2X1_255 ( .gnd(gnd), .vdd(vdd), .A(_1895_), .B(_1891_), .Y(_1896_) );
NOR2X1 NOR2X1_367 ( .gnd(gnd), .vdd(vdd), .A(_1894_), .B(_1896_), .Y(_1897_) );
NAND3X1 NAND3X1_85 ( .gnd(gnd), .vdd(vdd), .A(_1852_), .B(_1897_), .C(_1869_), .Y(_1898_) );
AOI21X1 AOI21X1_369 ( .gnd(gnd), .vdd(vdd), .A(_1898_), .B(_1893_), .C(_400__bF_buf11), .Y(_375__2_) );
AOI21X1 AOI21X1_370 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_3_bF_buf0_), .B(micro_hash_ucr_a_3_), .C(_1854_), .Y(_1899_) );
OAI22X1 OAI22X1_40 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_3_bF_buf3_), .B(micro_hash_ucr_a_3_), .C(_1899_), .D(_1892_), .Y(_1900_) );
NOR2X1 NOR2X1_368 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe33_bF_buf1), .B(_1877_), .Y(_1901_) );
NAND2X1 NAND2X1_256 ( .gnd(gnd), .vdd(vdd), .A(_928_), .B(_1296_), .Y(_1902_) );
NAND3X1 NAND3X1_86 ( .gnd(gnd), .vdd(vdd), .A(_876__bF_buf1), .B(micro_hash_ucr_x_3_), .C(_1874_), .Y(_1903_) );
NOR2X1 NOR2X1_369 ( .gnd(gnd), .vdd(vdd), .A(_1902_), .B(_1903_), .Y(_1904_) );
AND2X2 AND2X2_194 ( .gnd(gnd), .vdd(vdd), .A(_1860_), .B(_1904_), .Y(_1905_) );
NOR2X1 NOR2X1_370 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe19_bF_buf0), .B(micro_hash_ucr_pipe17_bF_buf0), .Y(_1906_) );
NAND3X1 NAND3X1_87 ( .gnd(gnd), .vdd(vdd), .A(_965_), .B(_1839_), .C(_1906_), .Y(_1907_) );
INVX2 INVX2_97 ( .gnd(gnd), .vdd(vdd), .A(_1865_), .Y(_1908_) );
NOR2X1 NOR2X1_371 ( .gnd(gnd), .vdd(vdd), .A(_1907_), .B(_1908_), .Y(_1909_) );
NAND3X1 NAND3X1_88 ( .gnd(gnd), .vdd(vdd), .A(_1901_), .B(_1909_), .C(_1905_), .Y(_1910_) );
AOI21X1 AOI21X1_371 ( .gnd(gnd), .vdd(vdd), .A(_1910_), .B(_1900_), .C(_400__bF_buf10), .Y(_375__3_) );
NOR2X1 NOR2X1_372 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_4_bF_buf3_), .B(micro_hash_ucr_a_4_), .Y(_1911_) );
OAI21X1 OAI21X1_510 ( .gnd(gnd), .vdd(vdd), .A(_1862_), .B(_1911_), .C(_1908_), .Y(_1912_) );
NAND2X1 NAND2X1_257 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_x_4_), .B(_1854_), .Y(_1913_) );
NOR2X1 NOR2X1_373 ( .gnd(gnd), .vdd(vdd), .A(_1395_), .B(_474__bF_buf2), .Y(_1914_) );
NOR2X1 NOR2X1_374 ( .gnd(gnd), .vdd(vdd), .A(_1911_), .B(_1914_), .Y(_1915_) );
AOI21X1 AOI21X1_372 ( .gnd(gnd), .vdd(vdd), .A(_1915_), .B(_1853_), .C(_1868_), .Y(_1916_) );
AOI22X1 AOI22X1_23 ( .gnd(gnd), .vdd(vdd), .A(_1868_), .B(_1911_), .C(_1913_), .D(_1916_), .Y(_1917_) );
OAI21X1 OAI21X1_511 ( .gnd(gnd), .vdd(vdd), .A(_1917_), .B(_1864_), .C(_1912_), .Y(_1918_) );
INVX1 INVX1_111 ( .gnd(gnd), .vdd(vdd), .A(_1911_), .Y(_1919_) );
AOI21X1 AOI21X1_373 ( .gnd(gnd), .vdd(vdd), .A(_1862_), .B(_1919_), .C(micro_hash_ucr_pipe69), .Y(_1920_) );
OAI21X1 OAI21X1_512 ( .gnd(gnd), .vdd(vdd), .A(_876__bF_buf0), .B(_1919_), .C(_302__bF_buf3), .Y(_1921_) );
AOI21X1 AOI21X1_374 ( .gnd(gnd), .vdd(vdd), .A(_1920_), .B(_1918_), .C(_1921_), .Y(_375__4_) );
AOI21X1 AOI21X1_375 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_5_bF_buf0_), .B(micro_hash_ucr_a_5_bF_buf3_), .C(_1854_), .Y(_1922_) );
OAI22X1 OAI22X1_41 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_5_bF_buf3_), .B(micro_hash_ucr_a_5_bF_buf2_), .C(_1922_), .D(_1892_), .Y(_1923_) );
NAND3X1 NAND3X1_89 ( .gnd(gnd), .vdd(vdd), .A(_910_), .B(_911__bF_buf4), .C(_915__bF_buf3), .Y(_1924_) );
NAND2X1 NAND2X1_258 ( .gnd(gnd), .vdd(vdd), .A(_1850_), .B(_1891_), .Y(_1925_) );
NOR2X1 NOR2X1_375 ( .gnd(gnd), .vdd(vdd), .A(_1924_), .B(_1925_), .Y(_1926_) );
NAND2X1 NAND2X1_259 ( .gnd(gnd), .vdd(vdd), .A(_1848_), .B(_1843_), .Y(_1927_) );
NAND3X1 NAND3X1_90 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_x_5_), .B(_971_), .C(_1844_), .Y(_1928_) );
NOR2X1 NOR2X1_376 ( .gnd(gnd), .vdd(vdd), .A(_1928_), .B(_1927_), .Y(_1929_) );
NAND3X1 NAND3X1_91 ( .gnd(gnd), .vdd(vdd), .A(_1926_), .B(_1929_), .C(_1869_), .Y(_1930_) );
AOI21X1 AOI21X1_376 ( .gnd(gnd), .vdd(vdd), .A(_1930_), .B(_1923_), .C(_400__bF_buf9), .Y(_375__5_) );
AOI21X1 AOI21X1_377 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_6_bF_buf0_), .B(micro_hash_ucr_a_6_bF_buf2_), .C(_1854_), .Y(_1931_) );
OAI22X1 OAI22X1_42 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_6_bF_buf3_), .B(micro_hash_ucr_a_6_bF_buf1_), .C(_1931_), .D(_1892_), .Y(_1932_) );
NAND3X1 NAND3X1_92 ( .gnd(gnd), .vdd(vdd), .A(_876__bF_buf3), .B(micro_hash_ucr_x_6_), .C(_1844_), .Y(_1933_) );
NOR2X1 NOR2X1_377 ( .gnd(gnd), .vdd(vdd), .A(_1924_), .B(_1933_), .Y(_1934_) );
NAND2X1 NAND2X1_260 ( .gnd(gnd), .vdd(vdd), .A(_971_), .B(_1850_), .Y(_1935_) );
OR2X2 OR2X2_29 ( .gnd(gnd), .vdd(vdd), .A(_1908_), .B(_1927_), .Y(_1936_) );
NOR2X1 NOR2X1_378 ( .gnd(gnd), .vdd(vdd), .A(_1935_), .B(_1936_), .Y(_1937_) );
NAND3X1 NAND3X1_93 ( .gnd(gnd), .vdd(vdd), .A(_1860_), .B(_1934_), .C(_1937_), .Y(_1938_) );
AOI21X1 AOI21X1_378 ( .gnd(gnd), .vdd(vdd), .A(_1938_), .B(_1932_), .C(_400__bF_buf8), .Y(_375__6_) );
NAND2X1 NAND2X1_261 ( .gnd(gnd), .vdd(vdd), .A(_1721__bF_buf3), .B(_1717__bF_buf1), .Y(_1939_) );
AOI21X1 AOI21X1_379 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_7_), .B(micro_hash_ucr_a_7_), .C(_1854_), .Y(_1940_) );
OAI21X1 OAI21X1_513 ( .gnd(gnd), .vdd(vdd), .A(_1940_), .B(_1866_), .C(_1939_), .Y(_1941_) );
AND2X2 AND2X2_195 ( .gnd(gnd), .vdd(vdd), .A(_1874_), .B(_910_), .Y(_1942_) );
NAND3X1 NAND3X1_94 ( .gnd(gnd), .vdd(vdd), .A(_1876_), .B(_1942_), .C(_1895_), .Y(_1943_) );
NOR2X1 NOR2X1_379 ( .gnd(gnd), .vdd(vdd), .A(_1935_), .B(_1943_), .Y(_1944_) );
NAND3X1 NAND3X1_95 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_x_7_), .B(_1861_), .C(_1870_), .Y(_1945_) );
NOR2X1 NOR2X1_380 ( .gnd(gnd), .vdd(vdd), .A(_1945_), .B(_1885_), .Y(_1946_) );
AOI21X1 AOI21X1_380 ( .gnd(gnd), .vdd(vdd), .A(_1944_), .B(_1946_), .C(micro_hash_ucr_pipe69), .Y(_1947_) );
OAI21X1 OAI21X1_514 ( .gnd(gnd), .vdd(vdd), .A(_876__bF_buf2), .B(_1939_), .C(_302__bF_buf2), .Y(_1948_) );
AOI21X1 AOI21X1_381 ( .gnd(gnd), .vdd(vdd), .A(_1947_), .B(_1941_), .C(_1948_), .Y(_375__7_) );
NOR2X1 NOR2X1_381 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe69), .B(_400__bF_buf7), .Y(_1949_) );
INVX4 INVX4_54 ( .gnd(gnd), .vdd(vdd), .A(_1949_), .Y(_1950_) );
INVX1 INVX1_112 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_232_), .Y(_1951_) );
NOR2X1 NOR2X1_382 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_k_0_), .B(micro_hash_ucr_x_0_), .Y(_1952_) );
NAND2X1 NAND2X1_262 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_k_0_), .B(micro_hash_ucr_x_0_), .Y(_1953_) );
INVX4 INVX4_55 ( .gnd(gnd), .vdd(vdd), .A(_1953_), .Y(_1954_) );
OAI21X1 OAI21X1_515 ( .gnd(gnd), .vdd(vdd), .A(_1954_), .B(_1952_), .C(_1951_), .Y(_1955_) );
NOR2X1 NOR2X1_383 ( .gnd(gnd), .vdd(vdd), .A(_1952_), .B(_1954_), .Y(_1956_) );
INVX8 INVX8_87 ( .gnd(gnd), .vdd(vdd), .A(_1956__bF_buf5), .Y(_1957_) );
NOR2X1 NOR2X1_384 ( .gnd(gnd), .vdd(vdd), .A(_1951_), .B(_1957__bF_buf3), .Y(_1958_) );
INVX2 INVX2_98 ( .gnd(gnd), .vdd(vdd), .A(_1958_), .Y(_1959_) );
NAND2X1 NAND2X1_263 ( .gnd(gnd), .vdd(vdd), .A(_1955_), .B(_1959_), .Y(_1960_) );
XNOR2X1 XNOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_1956__bF_buf4), .B(micro_hash_ucr_Wx_72_), .Y(_1961_) );
NOR2X1 NOR2X1_385 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_32_), .B(_1956__bF_buf3), .Y(_1962_) );
AND2X2 AND2X2_196 ( .gnd(gnd), .vdd(vdd), .A(_1956__bF_buf2), .B(micro_hash_ucr_Wx_32_), .Y(_1963_) );
OAI21X1 OAI21X1_516 ( .gnd(gnd), .vdd(vdd), .A(_1963_), .B(_1962_), .C(micro_hash_ucr_pipe16_bF_buf3), .Y(_1964_) );
NOR2X1 NOR2X1_386 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_8_), .B(_1956__bF_buf1), .Y(_1965_) );
NAND2X1 NAND2X1_264 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_8_), .B(_1956__bF_buf0), .Y(_1966_) );
INVX2 INVX2_99 ( .gnd(gnd), .vdd(vdd), .A(_1966_), .Y(_1967_) );
OAI21X1 OAI21X1_517 ( .gnd(gnd), .vdd(vdd), .A(_1967_), .B(_1965_), .C(micro_hash_ucr_pipe10), .Y(_1968_) );
INVX1 INVX1_113 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_0_), .Y(_1969_) );
NOR2X1 NOR2X1_387 ( .gnd(gnd), .vdd(vdd), .A(_1969_), .B(_1957__bF_buf2), .Y(_1970_) );
OAI21X1 OAI21X1_518 ( .gnd(gnd), .vdd(vdd), .A(_1956__bF_buf5), .B(micro_hash_ucr_Wx_0_), .C(micro_hash_ucr_pipe8), .Y(_1971_) );
NOR2X1 NOR2X1_388 ( .gnd(gnd), .vdd(vdd), .A(_1971_), .B(_1970_), .Y(_1972_) );
NOR2X1 NOR2X1_389 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_0_bF_buf0_), .B(micro_hash_ucr_pipe6), .Y(_1973_) );
OAI21X1 OAI21X1_519 ( .gnd(gnd), .vdd(vdd), .A(_937_), .B(H_16_), .C(_938_), .Y(_1974_) );
OAI21X1 OAI21X1_520 ( .gnd(gnd), .vdd(vdd), .A(_1974_), .B(_1973_), .C(_936_), .Y(_1975_) );
OAI21X1 OAI21X1_521 ( .gnd(gnd), .vdd(vdd), .A(_1972_), .B(_1975_), .C(_1968_), .Y(_1976_) );
XOR2X1 XOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_1956__bF_buf4), .B(micro_hash_ucr_Wx_16_), .Y(_1977_) );
AOI21X1 AOI21X1_382 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe12), .B(_1977_), .C(micro_hash_ucr_pipe14_bF_buf3), .Y(_1978_) );
OAI21X1 OAI21X1_522 ( .gnd(gnd), .vdd(vdd), .A(_1976_), .B(micro_hash_ucr_pipe12), .C(_1978_), .Y(_1979_) );
XOR2X1 XOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_1956__bF_buf3), .B(micro_hash_ucr_Wx_24_), .Y(_1980_) );
OAI21X1 OAI21X1_523 ( .gnd(gnd), .vdd(vdd), .A(_932_), .B(_1980_), .C(_1979_), .Y(_1981_) );
NAND2X1 NAND2X1_265 ( .gnd(gnd), .vdd(vdd), .A(_930__bF_buf2), .B(_1981_), .Y(_1982_) );
AND2X2 AND2X2_197 ( .gnd(gnd), .vdd(vdd), .A(_1982_), .B(_1964_), .Y(_1983_) );
NOR2X1 NOR2X1_390 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_40_), .B(_1956__bF_buf2), .Y(_1984_) );
AND2X2 AND2X2_198 ( .gnd(gnd), .vdd(vdd), .A(_1956__bF_buf1), .B(micro_hash_ucr_Wx_40_), .Y(_1985_) );
OAI21X1 OAI21X1_524 ( .gnd(gnd), .vdd(vdd), .A(_1985_), .B(_1984_), .C(micro_hash_ucr_pipe18_bF_buf3), .Y(_1986_) );
OAI21X1 OAI21X1_525 ( .gnd(gnd), .vdd(vdd), .A(_1983_), .B(micro_hash_ucr_pipe18_bF_buf2), .C(_1986_), .Y(_1987_) );
NOR2X1 NOR2X1_391 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe20_bF_buf0), .B(_1987_), .Y(_1988_) );
AND2X2 AND2X2_199 ( .gnd(gnd), .vdd(vdd), .A(_1956__bF_buf0), .B(micro_hash_ucr_Wx_48_), .Y(_1989_) );
OAI21X1 OAI21X1_526 ( .gnd(gnd), .vdd(vdd), .A(_1956__bF_buf5), .B(micro_hash_ucr_Wx_48_), .C(micro_hash_ucr_pipe20_bF_buf4), .Y(_1990_) );
OAI21X1 OAI21X1_527 ( .gnd(gnd), .vdd(vdd), .A(_1989_), .B(_1990_), .C(_924__bF_buf0), .Y(_1991_) );
NOR2X1 NOR2X1_392 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_56_), .B(_1956__bF_buf4), .Y(_1992_) );
NOR2X1 NOR2X1_393 ( .gnd(gnd), .vdd(vdd), .A(_807_), .B(_1957__bF_buf1), .Y(_1993_) );
OAI21X1 OAI21X1_528 ( .gnd(gnd), .vdd(vdd), .A(_1993_), .B(_1992_), .C(micro_hash_ucr_pipe22_bF_buf4), .Y(_1994_) );
OAI21X1 OAI21X1_529 ( .gnd(gnd), .vdd(vdd), .A(_1988_), .B(_1991_), .C(_1994_), .Y(_1995_) );
NAND2X1 NAND2X1_266 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_64_), .B(_1956__bF_buf3), .Y(_1996_) );
OAI21X1 OAI21X1_530 ( .gnd(gnd), .vdd(vdd), .A(_1954_), .B(_1952_), .C(_853_), .Y(_1997_) );
AOI21X1 AOI21X1_383 ( .gnd(gnd), .vdd(vdd), .A(_1997_), .B(_1996_), .C(_919__bF_buf4), .Y(_1998_) );
AOI21X1 AOI21X1_384 ( .gnd(gnd), .vdd(vdd), .A(_919__bF_buf3), .B(_1995_), .C(_1998_), .Y(_1999_) );
NAND2X1 NAND2X1_267 ( .gnd(gnd), .vdd(vdd), .A(_920__bF_buf4), .B(_1999_), .Y(_2000_) );
OAI21X1 OAI21X1_531 ( .gnd(gnd), .vdd(vdd), .A(_920__bF_buf3), .B(_1961_), .C(_2000_), .Y(_2001_) );
NOR2X1 NOR2X1_394 ( .gnd(gnd), .vdd(vdd), .A(_740_), .B(_1957__bF_buf0), .Y(_2002_) );
NOR2X1 NOR2X1_395 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_80_), .B(_1956__bF_buf2), .Y(_2003_) );
OAI21X1 OAI21X1_532 ( .gnd(gnd), .vdd(vdd), .A(_2002_), .B(_2003_), .C(micro_hash_ucr_pipe28_bF_buf1), .Y(_2004_) );
OAI21X1 OAI21X1_533 ( .gnd(gnd), .vdd(vdd), .A(_2001_), .B(micro_hash_ucr_pipe28_bF_buf0), .C(_2004_), .Y(_2005_) );
OAI21X1 OAI21X1_534 ( .gnd(gnd), .vdd(vdd), .A(_1954_), .B(_1952_), .C(_778_), .Y(_2006_) );
NOR2X1 NOR2X1_396 ( .gnd(gnd), .vdd(vdd), .A(_778_), .B(_1957__bF_buf3), .Y(_2007_) );
NOR2X1 NOR2X1_397 ( .gnd(gnd), .vdd(vdd), .A(_913__bF_buf1), .B(_2007_), .Y(_2008_) );
AOI21X1 AOI21X1_385 ( .gnd(gnd), .vdd(vdd), .A(_2006_), .B(_2008_), .C(micro_hash_ucr_pipe32_bF_buf2), .Y(_2009_) );
OAI21X1 OAI21X1_535 ( .gnd(gnd), .vdd(vdd), .A(_2005_), .B(micro_hash_ucr_pipe30_bF_buf1), .C(_2009_), .Y(_2010_) );
NOR2X1 NOR2X1_398 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_96_), .B(_1956__bF_buf1), .Y(_2011_) );
NOR2X1 NOR2X1_399 ( .gnd(gnd), .vdd(vdd), .A(_640_), .B(_1957__bF_buf2), .Y(_2012_) );
OAI21X1 OAI21X1_536 ( .gnd(gnd), .vdd(vdd), .A(_2012_), .B(_2011_), .C(micro_hash_ucr_pipe32_bF_buf1), .Y(_2013_) );
NAND3X1 NAND3X1_96 ( .gnd(gnd), .vdd(vdd), .A(_912__bF_buf4), .B(_2013_), .C(_2010_), .Y(_2014_) );
NOR2X1 NOR2X1_400 ( .gnd(gnd), .vdd(vdd), .A(_670_), .B(_1957__bF_buf1), .Y(_2015_) );
OAI21X1 OAI21X1_537 ( .gnd(gnd), .vdd(vdd), .A(_1956__bF_buf0), .B(micro_hash_ucr_Wx_104_), .C(micro_hash_ucr_pipe34_bF_buf3), .Y(_2016_) );
OAI21X1 OAI21X1_538 ( .gnd(gnd), .vdd(vdd), .A(_2015_), .B(_2016_), .C(_2014_), .Y(_2017_) );
XNOR2X1 XNOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_1956__bF_buf5), .B(micro_hash_ucr_Wx_112_), .Y(_2018_) );
AOI21X1 AOI21X1_386 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe36_bF_buf3), .B(_2018_), .C(micro_hash_ucr_pipe38_bF_buf3), .Y(_2019_) );
OAI21X1 OAI21X1_539 ( .gnd(gnd), .vdd(vdd), .A(_2017_), .B(micro_hash_ucr_pipe36_bF_buf2), .C(_2019_), .Y(_2020_) );
NOR2X1 NOR2X1_401 ( .gnd(gnd), .vdd(vdd), .A(_560_), .B(_1957__bF_buf0), .Y(_2021_) );
OAI21X1 OAI21X1_540 ( .gnd(gnd), .vdd(vdd), .A(_1956__bF_buf4), .B(micro_hash_ucr_Wx_120_), .C(micro_hash_ucr_pipe38_bF_buf2), .Y(_2022_) );
OAI21X1 OAI21X1_541 ( .gnd(gnd), .vdd(vdd), .A(_2021_), .B(_2022_), .C(_2020_), .Y(_2023_) );
NOR2X1 NOR2X1_402 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_128_), .B(_1956__bF_buf3), .Y(_2024_) );
NOR2X1 NOR2X1_403 ( .gnd(gnd), .vdd(vdd), .A(_531_), .B(_1957__bF_buf3), .Y(_2025_) );
OAI21X1 OAI21X1_542 ( .gnd(gnd), .vdd(vdd), .A(_2025_), .B(_2024_), .C(micro_hash_ucr_pipe40_bF_buf0), .Y(_2026_) );
OAI21X1 OAI21X1_543 ( .gnd(gnd), .vdd(vdd), .A(_2023_), .B(micro_hash_ucr_pipe40_bF_buf4), .C(_2026_), .Y(_2027_) );
NOR2X1 NOR2X1_404 ( .gnd(gnd), .vdd(vdd), .A(_779_), .B(_1957__bF_buf2), .Y(_2028_) );
OAI21X1 OAI21X1_544 ( .gnd(gnd), .vdd(vdd), .A(_1956__bF_buf2), .B(micro_hash_ucr_Wx_136_), .C(micro_hash_ucr_pipe42_bF_buf0), .Y(_2029_) );
OAI22X1 OAI22X1_43 ( .gnd(gnd), .vdd(vdd), .A(_2028_), .B(_2029_), .C(_2027_), .D(micro_hash_ucr_pipe42_bF_buf3), .Y(_2030_) );
NOR2X1 NOR2X1_405 ( .gnd(gnd), .vdd(vdd), .A(_611_), .B(_1957__bF_buf1), .Y(_2031_) );
OAI21X1 OAI21X1_545 ( .gnd(gnd), .vdd(vdd), .A(_1956__bF_buf1), .B(micro_hash_ucr_Wx_144_), .C(micro_hash_ucr_pipe44), .Y(_2032_) );
OAI21X1 OAI21X1_546 ( .gnd(gnd), .vdd(vdd), .A(_2031_), .B(_2032_), .C(_900__bF_buf3), .Y(_2033_) );
AOI21X1 AOI21X1_387 ( .gnd(gnd), .vdd(vdd), .A(_902__bF_buf1), .B(_2030_), .C(_2033_), .Y(_2034_) );
NOR2X1 NOR2X1_406 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_152_), .B(_1956__bF_buf0), .Y(_2035_) );
NAND2X1 NAND2X1_268 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_152_), .B(_1956__bF_buf5), .Y(_2036_) );
INVX2 INVX2_100 ( .gnd(gnd), .vdd(vdd), .A(_2036_), .Y(_2037_) );
OAI21X1 OAI21X1_547 ( .gnd(gnd), .vdd(vdd), .A(_2037_), .B(_2035_), .C(micro_hash_ucr_pipe46_bF_buf4), .Y(_2038_) );
NAND2X1 NAND2X1_269 ( .gnd(gnd), .vdd(vdd), .A(_895__bF_buf4), .B(_2038_), .Y(_2039_) );
NOR2X1 NOR2X1_407 ( .gnd(gnd), .vdd(vdd), .A(_719_), .B(_1957__bF_buf0), .Y(_2040_) );
OAI21X1 OAI21X1_548 ( .gnd(gnd), .vdd(vdd), .A(_1956__bF_buf4), .B(micro_hash_ucr_Wx_160_), .C(micro_hash_ucr_pipe48_bF_buf3), .Y(_2041_) );
OAI22X1 OAI22X1_44 ( .gnd(gnd), .vdd(vdd), .A(_2040_), .B(_2041_), .C(_2034_), .D(_2039_), .Y(_2042_) );
NOR2X1 NOR2X1_408 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_168_), .B(_1956__bF_buf3), .Y(_2043_) );
NAND2X1 NAND2X1_270 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_168_), .B(_1956__bF_buf2), .Y(_2044_) );
INVX2 INVX2_101 ( .gnd(gnd), .vdd(vdd), .A(_2044_), .Y(_2045_) );
OAI21X1 OAI21X1_549 ( .gnd(gnd), .vdd(vdd), .A(_2045_), .B(_2043_), .C(micro_hash_ucr_pipe50_bF_buf1), .Y(_2046_) );
OAI21X1 OAI21X1_550 ( .gnd(gnd), .vdd(vdd), .A(_2042_), .B(micro_hash_ucr_pipe50_bF_buf0), .C(_2046_), .Y(_2047_) );
OAI21X1 OAI21X1_551 ( .gnd(gnd), .vdd(vdd), .A(_1954_), .B(_1952_), .C(_587_), .Y(_2048_) );
NOR2X1 NOR2X1_409 ( .gnd(gnd), .vdd(vdd), .A(_587_), .B(_1957__bF_buf3), .Y(_2049_) );
NOR2X1 NOR2X1_410 ( .gnd(gnd), .vdd(vdd), .A(_894__bF_buf2), .B(_2049_), .Y(_2050_) );
AOI21X1 AOI21X1_388 ( .gnd(gnd), .vdd(vdd), .A(_2048_), .B(_2050_), .C(micro_hash_ucr_pipe54_bF_buf1), .Y(_2051_) );
OAI21X1 OAI21X1_552 ( .gnd(gnd), .vdd(vdd), .A(_2047_), .B(micro_hash_ucr_pipe52_bF_buf0), .C(_2051_), .Y(_2052_) );
NOR2X1 NOR2X1_411 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_184_), .B(_1956__bF_buf1), .Y(_2053_) );
NOR2X1 NOR2X1_412 ( .gnd(gnd), .vdd(vdd), .A(_641_), .B(_1957__bF_buf2), .Y(_2054_) );
OAI21X1 OAI21X1_553 ( .gnd(gnd), .vdd(vdd), .A(_2054_), .B(_2053_), .C(micro_hash_ucr_pipe54_bF_buf0), .Y(_2055_) );
NAND3X1 NAND3X1_97 ( .gnd(gnd), .vdd(vdd), .A(_890__bF_buf4), .B(_2055_), .C(_2052_), .Y(_2056_) );
NOR2X1 NOR2X1_413 ( .gnd(gnd), .vdd(vdd), .A(_612_), .B(_1957__bF_buf1), .Y(_2057_) );
OAI21X1 OAI21X1_554 ( .gnd(gnd), .vdd(vdd), .A(_1956__bF_buf0), .B(micro_hash_ucr_Wx_192_), .C(micro_hash_ucr_pipe56_bF_buf3), .Y(_2058_) );
OAI21X1 OAI21X1_555 ( .gnd(gnd), .vdd(vdd), .A(_2057_), .B(_2058_), .C(_2056_), .Y(_2059_) );
XNOR2X1 XNOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_1956__bF_buf5), .B(micro_hash_ucr_Wx_200_), .Y(_2060_) );
AOI21X1 AOI21X1_389 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe58_bF_buf2), .B(_2060_), .C(micro_hash_ucr_pipe60_bF_buf4), .Y(_2061_) );
OAI21X1 OAI21X1_556 ( .gnd(gnd), .vdd(vdd), .A(_2059_), .B(micro_hash_ucr_pipe58_bF_buf1), .C(_2061_), .Y(_2062_) );
AND2X2 AND2X2_200 ( .gnd(gnd), .vdd(vdd), .A(_1956__bF_buf4), .B(micro_hash_ucr_Wx_208_), .Y(_2063_) );
OAI21X1 OAI21X1_557 ( .gnd(gnd), .vdd(vdd), .A(_1956__bF_buf3), .B(micro_hash_ucr_Wx_208_), .C(micro_hash_ucr_pipe60_bF_buf3), .Y(_2064_) );
OAI21X1 OAI21X1_558 ( .gnd(gnd), .vdd(vdd), .A(_2063_), .B(_2064_), .C(_2062_), .Y(_2065_) );
NOR2X1 NOR2X1_414 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_216_), .B(_1956__bF_buf2), .Y(_2066_) );
NAND2X1 NAND2X1_271 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_216_), .B(_1956__bF_buf1), .Y(_2067_) );
INVX2 INVX2_102 ( .gnd(gnd), .vdd(vdd), .A(_2067_), .Y(_2068_) );
OAI21X1 OAI21X1_559 ( .gnd(gnd), .vdd(vdd), .A(_2068_), .B(_2066_), .C(micro_hash_ucr_pipe62_bF_buf1), .Y(_2069_) );
OAI21X1 OAI21X1_560 ( .gnd(gnd), .vdd(vdd), .A(_2065_), .B(micro_hash_ucr_pipe62_bF_buf0), .C(_2069_), .Y(_2070_) );
AND2X2 AND2X2_201 ( .gnd(gnd), .vdd(vdd), .A(_1956__bF_buf0), .B(micro_hash_ucr_Wx_224_), .Y(_2071_) );
OAI21X1 OAI21X1_561 ( .gnd(gnd), .vdd(vdd), .A(_1956__bF_buf5), .B(micro_hash_ucr_Wx_224_), .C(micro_hash_ucr_pipe64_bF_buf2), .Y(_2072_) );
OAI22X1 OAI22X1_45 ( .gnd(gnd), .vdd(vdd), .A(_2071_), .B(_2072_), .C(_2070_), .D(micro_hash_ucr_pipe64_bF_buf1), .Y(_2073_) );
NAND2X1 NAND2X1_272 ( .gnd(gnd), .vdd(vdd), .A(_877__bF_buf3), .B(_2073_), .Y(_2074_) );
OAI21X1 OAI21X1_562 ( .gnd(gnd), .vdd(vdd), .A(_877__bF_buf2), .B(_1960_), .C(_2074_), .Y(_2075_) );
NOR2X1 NOR2X1_415 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_240_), .B(_1956__bF_buf4), .Y(_2076_) );
AND2X2 AND2X2_202 ( .gnd(gnd), .vdd(vdd), .A(_1956__bF_buf3), .B(micro_hash_ucr_Wx_240_), .Y(_2077_) );
OAI21X1 OAI21X1_563 ( .gnd(gnd), .vdd(vdd), .A(_2077_), .B(_2076_), .C(micro_hash_ucr_pipe68), .Y(_2078_) );
OAI21X1 OAI21X1_564 ( .gnd(gnd), .vdd(vdd), .A(_2075_), .B(micro_hash_ucr_pipe68), .C(_2078_), .Y(_2079_) );
INVX2 INVX2_103 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_248_), .Y(_2080_) );
AOI21X1 AOI21X1_390 ( .gnd(gnd), .vdd(vdd), .A(_2080_), .B(_1957__bF_buf0), .C(_400__bF_buf6), .Y(_2081_) );
OAI21X1 OAI21X1_565 ( .gnd(gnd), .vdd(vdd), .A(_2080_), .B(_1957__bF_buf3), .C(_2081_), .Y(_2082_) );
AOI22X1 AOI22X1_24 ( .gnd(gnd), .vdd(vdd), .A(_1950_), .B(_2082_), .C(_2079_), .D(_876__bF_buf1), .Y(_299__0_) );
NOR2X1 NOR2X1_416 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_k_1_), .B(micro_hash_ucr_x_1_), .Y(_2083_) );
NAND2X1 NAND2X1_273 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_k_1_), .B(micro_hash_ucr_x_1_), .Y(_2084_) );
INVX1 INVX1_114 ( .gnd(gnd), .vdd(vdd), .A(_2084_), .Y(_2085_) );
NOR2X1 NOR2X1_417 ( .gnd(gnd), .vdd(vdd), .A(_2083_), .B(_2085_), .Y(_2086_) );
NAND2X1 NAND2X1_274 ( .gnd(gnd), .vdd(vdd), .A(_1954_), .B(_2086_), .Y(_2087_) );
OAI21X1 OAI21X1_566 ( .gnd(gnd), .vdd(vdd), .A(_2085_), .B(_2083_), .C(_1953_), .Y(_2088_) );
NAND2X1 NAND2X1_275 ( .gnd(gnd), .vdd(vdd), .A(_2088_), .B(_2087_), .Y(_2089_) );
INVX8 INVX8_88 ( .gnd(gnd), .vdd(vdd), .A(_2089__bF_buf5), .Y(_2090_) );
NOR2X1 NOR2X1_418 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_9_), .B(_2090__bF_buf4), .Y(_2091_) );
NAND2X1 NAND2X1_276 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_9_), .B(_2090__bF_buf3), .Y(_2092_) );
INVX1 INVX1_115 ( .gnd(gnd), .vdd(vdd), .A(_2092_), .Y(_2093_) );
NOR2X1 NOR2X1_419 ( .gnd(gnd), .vdd(vdd), .A(_2091_), .B(_2093_), .Y(_2094_) );
XNOR2X1 XNOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_2094_), .B(_1967_), .Y(_2095_) );
NAND2X1 NAND2X1_277 ( .gnd(gnd), .vdd(vdd), .A(H_17_), .B(micro_hash_ucr_pipe6), .Y(_2096_) );
OAI21X1 OAI21X1_567 ( .gnd(gnd), .vdd(vdd), .A(_1058__bF_buf2), .B(micro_hash_ucr_pipe6), .C(_2096_), .Y(_2097_) );
INVX1 INVX1_116 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_1_), .Y(_2098_) );
NAND2X1 NAND2X1_278 ( .gnd(gnd), .vdd(vdd), .A(_2098_), .B(_2089__bF_buf4), .Y(_2099_) );
INVX1 INVX1_117 ( .gnd(gnd), .vdd(vdd), .A(_2099_), .Y(_2100_) );
NOR2X1 NOR2X1_420 ( .gnd(gnd), .vdd(vdd), .A(_2098_), .B(_2089__bF_buf3), .Y(_2101_) );
NOR2X1 NOR2X1_421 ( .gnd(gnd), .vdd(vdd), .A(_2101_), .B(_2100_), .Y(_2102_) );
AND2X2 AND2X2_203 ( .gnd(gnd), .vdd(vdd), .A(_2102_), .B(_1970_), .Y(_2103_) );
NOR2X1 NOR2X1_422 ( .gnd(gnd), .vdd(vdd), .A(_1970_), .B(_2102_), .Y(_2104_) );
OAI21X1 OAI21X1_568 ( .gnd(gnd), .vdd(vdd), .A(_2104_), .B(_2103_), .C(micro_hash_ucr_pipe8), .Y(_2105_) );
OAI21X1 OAI21X1_569 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe8), .B(_2097_), .C(_2105_), .Y(_2106_) );
MUX2X1 MUX2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_2106_), .B(_2095_), .S(_936_), .Y(_2107_) );
NAND2X1 NAND2X1_279 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_16_), .B(_1956__bF_buf2), .Y(_2108_) );
NOR2X1 NOR2X1_423 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_17_), .B(_2090__bF_buf2), .Y(_2109_) );
INVX1 INVX1_118 ( .gnd(gnd), .vdd(vdd), .A(_2109_), .Y(_2110_) );
NAND2X1 NAND2X1_280 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_17_), .B(_2090__bF_buf1), .Y(_2111_) );
NAND2X1 NAND2X1_281 ( .gnd(gnd), .vdd(vdd), .A(_2111_), .B(_2110_), .Y(_2112_) );
XOR2X1 XOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_2112_), .B(_2108_), .Y(_2113_) );
MUX2X1 MUX2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_2107_), .B(_2113_), .S(_931_), .Y(_2114_) );
NAND2X1 NAND2X1_282 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_24_), .B(_1956__bF_buf1), .Y(_2115_) );
NOR2X1 NOR2X1_424 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_25_), .B(_2090__bF_buf0), .Y(_2116_) );
INVX1 INVX1_119 ( .gnd(gnd), .vdd(vdd), .A(_2116_), .Y(_2117_) );
NAND2X1 NAND2X1_283 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_25_), .B(_2090__bF_buf4), .Y(_2118_) );
NAND2X1 NAND2X1_284 ( .gnd(gnd), .vdd(vdd), .A(_2118_), .B(_2117_), .Y(_2119_) );
XNOR2X1 XNOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_2119_), .B(_2115_), .Y(_2120_) );
MUX2X1 MUX2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_2114_), .B(_2120_), .S(_932_), .Y(_2121_) );
XNOR2X1 XNOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_2089__bF_buf2), .B(micro_hash_ucr_Wx_33_), .Y(_2122_) );
XOR2X1 XOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_2122_), .B(_1963_), .Y(_2123_) );
MUX2X1 MUX2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_2121_), .B(_2123_), .S(_930__bF_buf1), .Y(_2124_) );
XNOR2X1 XNOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_2089__bF_buf1), .B(micro_hash_ucr_Wx_41_), .Y(_2125_) );
NAND2X1 NAND2X1_285 ( .gnd(gnd), .vdd(vdd), .A(_1985_), .B(_2125_), .Y(_2126_) );
OR2X2 OR2X2_30 ( .gnd(gnd), .vdd(vdd), .A(_2125_), .B(_1985_), .Y(_2127_) );
NAND3X1 NAND3X1_98 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe18_bF_buf1), .B(_2126_), .C(_2127_), .Y(_2128_) );
OAI21X1 OAI21X1_570 ( .gnd(gnd), .vdd(vdd), .A(_2124_), .B(micro_hash_ucr_pipe18_bF_buf0), .C(_2128_), .Y(_2129_) );
NOR2X1 NOR2X1_425 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_49_), .B(_2090__bF_buf3), .Y(_2130_) );
AND2X2 AND2X2_204 ( .gnd(gnd), .vdd(vdd), .A(_2090__bF_buf2), .B(micro_hash_ucr_Wx_49_), .Y(_2131_) );
NOR2X1 NOR2X1_426 ( .gnd(gnd), .vdd(vdd), .A(_2130_), .B(_2131_), .Y(_2132_) );
AND2X2 AND2X2_205 ( .gnd(gnd), .vdd(vdd), .A(_2132_), .B(_1989_), .Y(_2133_) );
OAI21X1 OAI21X1_571 ( .gnd(gnd), .vdd(vdd), .A(_2132_), .B(_1989_), .C(micro_hash_ucr_pipe20_bF_buf3), .Y(_2134_) );
OAI21X1 OAI21X1_572 ( .gnd(gnd), .vdd(vdd), .A(_2133_), .B(_2134_), .C(_924__bF_buf4), .Y(_2135_) );
AOI21X1 AOI21X1_391 ( .gnd(gnd), .vdd(vdd), .A(_926__bF_buf4), .B(_2129_), .C(_2135_), .Y(_2136_) );
NOR2X1 NOR2X1_427 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_57_), .B(_2090__bF_buf1), .Y(_2137_) );
NOR2X1 NOR2X1_428 ( .gnd(gnd), .vdd(vdd), .A(_810_), .B(_2089__bF_buf0), .Y(_2138_) );
NOR2X1 NOR2X1_429 ( .gnd(gnd), .vdd(vdd), .A(_2138_), .B(_2137_), .Y(_2139_) );
AND2X2 AND2X2_206 ( .gnd(gnd), .vdd(vdd), .A(_2139_), .B(_1993_), .Y(_2140_) );
NOR2X1 NOR2X1_430 ( .gnd(gnd), .vdd(vdd), .A(_1993_), .B(_2139_), .Y(_2141_) );
OAI21X1 OAI21X1_573 ( .gnd(gnd), .vdd(vdd), .A(_2140_), .B(_2141_), .C(micro_hash_ucr_pipe22_bF_buf3), .Y(_2142_) );
NAND2X1 NAND2X1_286 ( .gnd(gnd), .vdd(vdd), .A(_919__bF_buf2), .B(_2142_), .Y(_2143_) );
NOR2X1 NOR2X1_431 ( .gnd(gnd), .vdd(vdd), .A(_2143_), .B(_2136_), .Y(_2144_) );
XNOR2X1 XNOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_2089__bF_buf5), .B(_856_), .Y(_2145_) );
NOR2X1 NOR2X1_432 ( .gnd(gnd), .vdd(vdd), .A(_1996_), .B(_2145_), .Y(_2146_) );
INVX1 INVX1_120 ( .gnd(gnd), .vdd(vdd), .A(_2146_), .Y(_2147_) );
AOI21X1 AOI21X1_392 ( .gnd(gnd), .vdd(vdd), .A(_1996_), .B(_2145_), .C(_919__bF_buf1), .Y(_2148_) );
AOI21X1 AOI21X1_393 ( .gnd(gnd), .vdd(vdd), .A(_2147_), .B(_2148_), .C(_2144_), .Y(_2149_) );
NOR2X1 NOR2X1_433 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_73_), .B(_2090__bF_buf0), .Y(_2150_) );
NOR2X1 NOR2X1_434 ( .gnd(gnd), .vdd(vdd), .A(_832_), .B(_2089__bF_buf4), .Y(_2151_) );
NOR2X1 NOR2X1_435 ( .gnd(gnd), .vdd(vdd), .A(_2151_), .B(_2150_), .Y(_2152_) );
NAND3X1 NAND3X1_99 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_72_), .B(_1956__bF_buf0), .C(_2152_), .Y(_2153_) );
INVX1 INVX1_121 ( .gnd(gnd), .vdd(vdd), .A(_2152_), .Y(_2154_) );
OAI21X1 OAI21X1_574 ( .gnd(gnd), .vdd(vdd), .A(_829_), .B(_1957__bF_buf2), .C(_2154_), .Y(_2155_) );
NAND3X1 NAND3X1_100 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe26_bF_buf3), .B(_2153_), .C(_2155_), .Y(_2156_) );
OAI21X1 OAI21X1_575 ( .gnd(gnd), .vdd(vdd), .A(_2149_), .B(micro_hash_ucr_pipe26_bF_buf2), .C(_2156_), .Y(_2157_) );
XNOR2X1 XNOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_2089__bF_buf3), .B(micro_hash_ucr_Wx_81_), .Y(_2158_) );
NOR2X1 NOR2X1_436 ( .gnd(gnd), .vdd(vdd), .A(_2002_), .B(_2158_), .Y(_2159_) );
NAND2X1 NAND2X1_287 ( .gnd(gnd), .vdd(vdd), .A(_2002_), .B(_2158_), .Y(_2160_) );
NAND2X1 NAND2X1_288 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe28_bF_buf3), .B(_2160_), .Y(_2161_) );
OAI21X1 OAI21X1_576 ( .gnd(gnd), .vdd(vdd), .A(_2161_), .B(_2159_), .C(_913__bF_buf0), .Y(_2162_) );
AOI21X1 AOI21X1_394 ( .gnd(gnd), .vdd(vdd), .A(_918__bF_buf2), .B(_2157_), .C(_2162_), .Y(_2163_) );
NOR2X1 NOR2X1_437 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_89_), .B(_2090__bF_buf4), .Y(_2164_) );
NOR2X1 NOR2X1_438 ( .gnd(gnd), .vdd(vdd), .A(_782_), .B(_2089__bF_buf2), .Y(_2165_) );
NOR2X1 NOR2X1_439 ( .gnd(gnd), .vdd(vdd), .A(_2165_), .B(_2164_), .Y(_2166_) );
AND2X2 AND2X2_207 ( .gnd(gnd), .vdd(vdd), .A(_2166_), .B(_2007_), .Y(_2167_) );
NOR2X1 NOR2X1_440 ( .gnd(gnd), .vdd(vdd), .A(_2007_), .B(_2166_), .Y(_2168_) );
OAI21X1 OAI21X1_577 ( .gnd(gnd), .vdd(vdd), .A(_2167_), .B(_2168_), .C(micro_hash_ucr_pipe30_bF_buf0), .Y(_2169_) );
NAND2X1 NAND2X1_289 ( .gnd(gnd), .vdd(vdd), .A(_914__bF_buf1), .B(_2169_), .Y(_2170_) );
XNOR2X1 XNOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_2089__bF_buf1), .B(micro_hash_ucr_Wx_97_), .Y(_2171_) );
OAI21X1 OAI21X1_578 ( .gnd(gnd), .vdd(vdd), .A(_2171_), .B(_2012_), .C(micro_hash_ucr_pipe32_bF_buf0), .Y(_2172_) );
AOI21X1 AOI21X1_395 ( .gnd(gnd), .vdd(vdd), .A(_2012_), .B(_2171_), .C(_2172_), .Y(_2173_) );
NOR2X1 NOR2X1_441 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe34_bF_buf2), .B(_2173_), .Y(_2174_) );
OAI21X1 OAI21X1_579 ( .gnd(gnd), .vdd(vdd), .A(_2163_), .B(_2170_), .C(_2174_), .Y(_2175_) );
NOR2X1 NOR2X1_442 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_105_), .B(_2090__bF_buf3), .Y(_2176_) );
NOR2X1 NOR2X1_443 ( .gnd(gnd), .vdd(vdd), .A(_673_), .B(_2089__bF_buf0), .Y(_2177_) );
NOR2X1 NOR2X1_444 ( .gnd(gnd), .vdd(vdd), .A(_2177_), .B(_2176_), .Y(_2178_) );
XOR2X1 XOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_2178_), .B(_2015_), .Y(_2179_) );
OAI21X1 OAI21X1_580 ( .gnd(gnd), .vdd(vdd), .A(_912__bF_buf3), .B(_2179_), .C(_2175_), .Y(_2180_) );
NOR2X1 NOR2X1_445 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe36_bF_buf1), .B(_2180_), .Y(_2181_) );
NOR2X1 NOR2X1_446 ( .gnd(gnd), .vdd(vdd), .A(_503_), .B(_1957__bF_buf1), .Y(_2182_) );
XNOR2X1 XNOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_2089__bF_buf5), .B(micro_hash_ucr_Wx_113_), .Y(_2183_) );
NOR2X1 NOR2X1_447 ( .gnd(gnd), .vdd(vdd), .A(_2182_), .B(_2183_), .Y(_2184_) );
NAND2X1 NAND2X1_290 ( .gnd(gnd), .vdd(vdd), .A(_2182_), .B(_2183_), .Y(_2185_) );
NAND2X1 NAND2X1_291 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe36_bF_buf0), .B(_2185_), .Y(_2186_) );
OAI21X1 OAI21X1_581 ( .gnd(gnd), .vdd(vdd), .A(_2186_), .B(_2184_), .C(_908__bF_buf4), .Y(_2187_) );
NOR2X1 NOR2X1_448 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_121_), .B(_2090__bF_buf2), .Y(_2188_) );
NOR2X1 NOR2X1_449 ( .gnd(gnd), .vdd(vdd), .A(_563_), .B(_2089__bF_buf4), .Y(_2189_) );
NOR2X1 NOR2X1_450 ( .gnd(gnd), .vdd(vdd), .A(_2189_), .B(_2188_), .Y(_2190_) );
XOR2X1 XOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_2190_), .B(_2021_), .Y(_2191_) );
OAI22X1 OAI22X1_46 ( .gnd(gnd), .vdd(vdd), .A(_908__bF_buf3), .B(_2191_), .C(_2181_), .D(_2187_), .Y(_2192_) );
XNOR2X1 XNOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_2089__bF_buf3), .B(micro_hash_ucr_Wx_129_), .Y(_2193_) );
XOR2X1 XOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_2193_), .B(_2025_), .Y(_2194_) );
AOI21X1 AOI21X1_396 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe40_bF_buf3), .B(_2194_), .C(micro_hash_ucr_pipe42_bF_buf2), .Y(_2195_) );
OAI21X1 OAI21X1_582 ( .gnd(gnd), .vdd(vdd), .A(_2192_), .B(micro_hash_ucr_pipe40_bF_buf2), .C(_2195_), .Y(_2196_) );
INVX1 INVX1_122 ( .gnd(gnd), .vdd(vdd), .A(_2028_), .Y(_2197_) );
NOR2X1 NOR2X1_451 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_137_), .B(_2090__bF_buf1), .Y(_2198_) );
INVX1 INVX1_123 ( .gnd(gnd), .vdd(vdd), .A(_2198_), .Y(_2199_) );
NOR2X1 NOR2X1_452 ( .gnd(gnd), .vdd(vdd), .A(_783_), .B(_2089__bF_buf2), .Y(_2200_) );
INVX2 INVX2_104 ( .gnd(gnd), .vdd(vdd), .A(_2200_), .Y(_2201_) );
NAND2X1 NAND2X1_292 ( .gnd(gnd), .vdd(vdd), .A(_2201_), .B(_2199_), .Y(_2202_) );
NOR2X1 NOR2X1_453 ( .gnd(gnd), .vdd(vdd), .A(_2197_), .B(_2202_), .Y(_2203_) );
AOI21X1 AOI21X1_397 ( .gnd(gnd), .vdd(vdd), .A(_2201_), .B(_2199_), .C(_2028_), .Y(_2204_) );
OAI21X1 OAI21X1_583 ( .gnd(gnd), .vdd(vdd), .A(_2203_), .B(_2204_), .C(micro_hash_ucr_pipe42_bF_buf1), .Y(_2205_) );
NAND3X1 NAND3X1_101 ( .gnd(gnd), .vdd(vdd), .A(_902__bF_buf0), .B(_2205_), .C(_2196_), .Y(_2206_) );
NOR2X1 NOR2X1_454 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_145_), .B(_2090__bF_buf0), .Y(_2207_) );
NOR2X1 NOR2X1_455 ( .gnd(gnd), .vdd(vdd), .A(_615_), .B(_2089__bF_buf1), .Y(_2208_) );
NOR2X1 NOR2X1_456 ( .gnd(gnd), .vdd(vdd), .A(_2208_), .B(_2207_), .Y(_2209_) );
NAND2X1 NAND2X1_293 ( .gnd(gnd), .vdd(vdd), .A(_2031_), .B(_2209_), .Y(_2210_) );
INVX1 INVX1_124 ( .gnd(gnd), .vdd(vdd), .A(_2210_), .Y(_2211_) );
OAI21X1 OAI21X1_584 ( .gnd(gnd), .vdd(vdd), .A(_2209_), .B(_2031_), .C(micro_hash_ucr_pipe44), .Y(_2212_) );
OAI21X1 OAI21X1_585 ( .gnd(gnd), .vdd(vdd), .A(_2211_), .B(_2212_), .C(_2206_), .Y(_2213_) );
NOR2X1 NOR2X1_457 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe46_bF_buf3), .B(_2213_), .Y(_2214_) );
NOR2X1 NOR2X1_458 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_153_), .B(_2090__bF_buf4), .Y(_2215_) );
INVX1 INVX1_125 ( .gnd(gnd), .vdd(vdd), .A(_2215_), .Y(_2216_) );
NAND2X1 NAND2X1_294 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_153_), .B(_2090__bF_buf3), .Y(_2217_) );
NAND2X1 NAND2X1_295 ( .gnd(gnd), .vdd(vdd), .A(_2217_), .B(_2216_), .Y(_2218_) );
XNOR2X1 XNOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(_2218_), .B(_2037_), .Y(_2219_) );
OAI21X1 OAI21X1_586 ( .gnd(gnd), .vdd(vdd), .A(_2219_), .B(_900__bF_buf2), .C(_895__bF_buf3), .Y(_2220_) );
NOR2X1 NOR2X1_459 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_161_), .B(_2090__bF_buf2), .Y(_2221_) );
NOR2X1 NOR2X1_460 ( .gnd(gnd), .vdd(vdd), .A(_722_), .B(_2089__bF_buf0), .Y(_2222_) );
NOR2X1 NOR2X1_461 ( .gnd(gnd), .vdd(vdd), .A(_2222_), .B(_2221_), .Y(_2223_) );
NAND2X1 NAND2X1_296 ( .gnd(gnd), .vdd(vdd), .A(_2040_), .B(_2223_), .Y(_2224_) );
INVX1 INVX1_126 ( .gnd(gnd), .vdd(vdd), .A(_2224_), .Y(_2225_) );
OAI21X1 OAI21X1_587 ( .gnd(gnd), .vdd(vdd), .A(_2223_), .B(_2040_), .C(micro_hash_ucr_pipe48_bF_buf2), .Y(_2226_) );
OAI22X1 OAI22X1_47 ( .gnd(gnd), .vdd(vdd), .A(_2225_), .B(_2226_), .C(_2214_), .D(_2220_), .Y(_2227_) );
NOR2X1 NOR2X1_462 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_169_), .B(_2090__bF_buf1), .Y(_2228_) );
NOR2X1 NOR2X1_463 ( .gnd(gnd), .vdd(vdd), .A(_699_), .B(_2089__bF_buf5), .Y(_2229_) );
NOR2X1 NOR2X1_464 ( .gnd(gnd), .vdd(vdd), .A(_2229_), .B(_2228_), .Y(_2230_) );
NAND2X1 NAND2X1_297 ( .gnd(gnd), .vdd(vdd), .A(_2045_), .B(_2230_), .Y(_2231_) );
INVX1 INVX1_127 ( .gnd(gnd), .vdd(vdd), .A(_2231_), .Y(_2232_) );
NOR2X1 NOR2X1_465 ( .gnd(gnd), .vdd(vdd), .A(_2045_), .B(_2230_), .Y(_2233_) );
OAI21X1 OAI21X1_588 ( .gnd(gnd), .vdd(vdd), .A(_2232_), .B(_2233_), .C(micro_hash_ucr_pipe50_bF_buf3), .Y(_2234_) );
OAI21X1 OAI21X1_589 ( .gnd(gnd), .vdd(vdd), .A(_2227_), .B(micro_hash_ucr_pipe50_bF_buf2), .C(_2234_), .Y(_2235_) );
NOR2X1 NOR2X1_466 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_177_), .B(_2090__bF_buf0), .Y(_2236_) );
NOR2X1 NOR2X1_467 ( .gnd(gnd), .vdd(vdd), .A(_590_), .B(_2089__bF_buf4), .Y(_2237_) );
NOR2X1 NOR2X1_468 ( .gnd(gnd), .vdd(vdd), .A(_2237_), .B(_2236_), .Y(_2238_) );
NOR2X1 NOR2X1_469 ( .gnd(gnd), .vdd(vdd), .A(_2049_), .B(_2238_), .Y(_2239_) );
NAND2X1 NAND2X1_298 ( .gnd(gnd), .vdd(vdd), .A(_2049_), .B(_2238_), .Y(_2240_) );
INVX1 INVX1_128 ( .gnd(gnd), .vdd(vdd), .A(_2240_), .Y(_2241_) );
NOR2X1 NOR2X1_470 ( .gnd(gnd), .vdd(vdd), .A(_2239_), .B(_2241_), .Y(_2242_) );
AOI21X1 AOI21X1_398 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe52_bF_buf4), .B(_2242_), .C(micro_hash_ucr_pipe54_bF_buf3), .Y(_2243_) );
OAI21X1 OAI21X1_590 ( .gnd(gnd), .vdd(vdd), .A(_2235_), .B(micro_hash_ucr_pipe52_bF_buf3), .C(_2243_), .Y(_2244_) );
XNOR2X1 XNOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_2089__bF_buf3), .B(micro_hash_ucr_Wx_185_), .Y(_2245_) );
XNOR2X1 XNOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_2245_), .B(_2054_), .Y(_2246_) );
AOI21X1 AOI21X1_399 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe54_bF_buf2), .B(_2246_), .C(micro_hash_ucr_pipe56_bF_buf2), .Y(_2247_) );
NOR2X1 NOR2X1_471 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_193_), .B(_2090__bF_buf4), .Y(_2248_) );
NOR2X1 NOR2X1_472 ( .gnd(gnd), .vdd(vdd), .A(_616_), .B(_2089__bF_buf2), .Y(_2249_) );
NOR2X1 NOR2X1_473 ( .gnd(gnd), .vdd(vdd), .A(_2249_), .B(_2248_), .Y(_2250_) );
NAND2X1 NAND2X1_299 ( .gnd(gnd), .vdd(vdd), .A(_2057_), .B(_2250_), .Y(_2251_) );
INVX1 INVX1_129 ( .gnd(gnd), .vdd(vdd), .A(_2251_), .Y(_2252_) );
NOR2X1 NOR2X1_474 ( .gnd(gnd), .vdd(vdd), .A(_2057_), .B(_2250_), .Y(_2253_) );
NOR2X1 NOR2X1_475 ( .gnd(gnd), .vdd(vdd), .A(_2253_), .B(_2252_), .Y(_2254_) );
AOI22X1 AOI22X1_25 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe56_bF_buf1), .B(_2254_), .C(_2244_), .D(_2247_), .Y(_2255_) );
NAND2X1 NAND2X1_300 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_200_), .B(_1956__bF_buf5), .Y(_2256_) );
XNOR2X1 XNOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_2089__bF_buf1), .B(_507_), .Y(_2257_) );
NOR2X1 NOR2X1_476 ( .gnd(gnd), .vdd(vdd), .A(_2256_), .B(_2257_), .Y(_2258_) );
INVX1 INVX1_130 ( .gnd(gnd), .vdd(vdd), .A(_2258_), .Y(_2259_) );
AOI21X1 AOI21X1_400 ( .gnd(gnd), .vdd(vdd), .A(_2256_), .B(_2257_), .C(_888__bF_buf1), .Y(_2260_) );
AOI21X1 AOI21X1_401 ( .gnd(gnd), .vdd(vdd), .A(_2260_), .B(_2259_), .C(micro_hash_ucr_pipe60_bF_buf2), .Y(_2261_) );
OAI21X1 OAI21X1_591 ( .gnd(gnd), .vdd(vdd), .A(_2255_), .B(micro_hash_ucr_pipe58_bF_buf0), .C(_2261_), .Y(_2262_) );
NAND2X1 NAND2X1_301 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_208_), .B(_1956__bF_buf4), .Y(_2263_) );
NOR2X1 NOR2X1_477 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_209_), .B(_2090__bF_buf3), .Y(_2264_) );
INVX1 INVX1_131 ( .gnd(gnd), .vdd(vdd), .A(_2264_), .Y(_2265_) );
NAND2X1 NAND2X1_302 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_209_), .B(_2090__bF_buf2), .Y(_2266_) );
NAND2X1 NAND2X1_303 ( .gnd(gnd), .vdd(vdd), .A(_2266_), .B(_2265_), .Y(_2267_) );
XNOR2X1 XNOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(_2267_), .B(_2263_), .Y(_2268_) );
AOI21X1 AOI21X1_402 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe60_bF_buf1), .B(_2268_), .C(micro_hash_ucr_pipe62_bF_buf4), .Y(_2269_) );
NOR2X1 NOR2X1_478 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_217_), .B(_2090__bF_buf1), .Y(_2270_) );
NOR2X1 NOR2X1_479 ( .gnd(gnd), .vdd(vdd), .A(_535_), .B(_2089__bF_buf0), .Y(_2271_) );
NOR2X1 NOR2X1_480 ( .gnd(gnd), .vdd(vdd), .A(_2271_), .B(_2270_), .Y(_2272_) );
NAND2X1 NAND2X1_304 ( .gnd(gnd), .vdd(vdd), .A(_2068_), .B(_2272_), .Y(_2273_) );
INVX1 INVX1_132 ( .gnd(gnd), .vdd(vdd), .A(_2273_), .Y(_2274_) );
NOR2X1 NOR2X1_481 ( .gnd(gnd), .vdd(vdd), .A(_2068_), .B(_2272_), .Y(_2275_) );
NOR2X1 NOR2X1_482 ( .gnd(gnd), .vdd(vdd), .A(_2275_), .B(_2274_), .Y(_2276_) );
AOI22X1 AOI22X1_26 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe62_bF_buf3), .B(_2276_), .C(_2262_), .D(_2269_), .Y(_2277_) );
XNOR2X1 XNOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_2089__bF_buf5), .B(micro_hash_ucr_Wx_225_), .Y(_2278_) );
XOR2X1 XOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_2278_), .B(_2071_), .Y(_2279_) );
AOI21X1 AOI21X1_403 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe64_bF_buf0), .B(_2279_), .C(micro_hash_ucr_pipe66_bF_buf4), .Y(_2280_) );
OAI21X1 OAI21X1_592 ( .gnd(gnd), .vdd(vdd), .A(_2277_), .B(micro_hash_ucr_pipe64_bF_buf4), .C(_2280_), .Y(_2281_) );
NOR2X1 NOR2X1_483 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_233_), .B(_2090__bF_buf0), .Y(_2282_) );
INVX1 INVX1_133 ( .gnd(gnd), .vdd(vdd), .A(_2282_), .Y(_2283_) );
NAND2X1 NAND2X1_305 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_233_), .B(_2090__bF_buf4), .Y(_2284_) );
NAND2X1 NAND2X1_306 ( .gnd(gnd), .vdd(vdd), .A(_2284_), .B(_2283_), .Y(_2285_) );
NOR2X1 NOR2X1_484 ( .gnd(gnd), .vdd(vdd), .A(_1959_), .B(_2285_), .Y(_2286_) );
AOI21X1 AOI21X1_404 ( .gnd(gnd), .vdd(vdd), .A(_2284_), .B(_2283_), .C(_1958_), .Y(_2287_) );
OAI21X1 OAI21X1_593 ( .gnd(gnd), .vdd(vdd), .A(_2286_), .B(_2287_), .C(micro_hash_ucr_pipe66_bF_buf3), .Y(_2288_) );
NAND3X1 NAND3X1_102 ( .gnd(gnd), .vdd(vdd), .A(_878__bF_buf4), .B(_2288_), .C(_2281_), .Y(_2289_) );
XNOR2X1 XNOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(_2089__bF_buf4), .B(micro_hash_ucr_Wx_241_), .Y(_2290_) );
XOR2X1 XOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_2290_), .B(_2077_), .Y(_2291_) );
AOI21X1 AOI21X1_405 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe68), .B(_2291_), .C(micro_hash_ucr_pipe69), .Y(_2292_) );
NOR2X1 NOR2X1_485 ( .gnd(gnd), .vdd(vdd), .A(_2080_), .B(_1957__bF_buf0), .Y(_2293_) );
NOR2X1 NOR2X1_486 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_249_), .B(_2090__bF_buf3), .Y(_2294_) );
INVX1 INVX1_134 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_249_), .Y(_2295_) );
NOR2X1 NOR2X1_487 ( .gnd(gnd), .vdd(vdd), .A(_2295_), .B(_2089__bF_buf3), .Y(_2296_) );
NOR2X1 NOR2X1_488 ( .gnd(gnd), .vdd(vdd), .A(_2296_), .B(_2294_), .Y(_2297_) );
AOI21X1 AOI21X1_406 ( .gnd(gnd), .vdd(vdd), .A(_2293_), .B(_2297_), .C(_400__bF_buf5), .Y(_2298_) );
OAI21X1 OAI21X1_594 ( .gnd(gnd), .vdd(vdd), .A(_2293_), .B(_2297_), .C(_2298_), .Y(_2299_) );
AOI22X1 AOI22X1_27 ( .gnd(gnd), .vdd(vdd), .A(_1950_), .B(_2299_), .C(_2289_), .D(_2292_), .Y(_299__1_) );
NOR2X1 NOR2X1_489 ( .gnd(gnd), .vdd(vdd), .A(_2101_), .B(_2103_), .Y(_2300_) );
OAI21X1 OAI21X1_595 ( .gnd(gnd), .vdd(vdd), .A(_2083_), .B(_1953_), .C(_2084_), .Y(_2301_) );
XOR2X1 XOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_k_2_), .B(micro_hash_ucr_x_2_), .Y(_2302_) );
NAND2X1 NAND2X1_307 ( .gnd(gnd), .vdd(vdd), .A(_2302_), .B(_2301_), .Y(_2303_) );
INVX8 INVX8_89 ( .gnd(gnd), .vdd(vdd), .A(_2303_), .Y(_2304_) );
NOR2X1 NOR2X1_490 ( .gnd(gnd), .vdd(vdd), .A(_2302_), .B(_2301_), .Y(_2305_) );
NOR2X1 NOR2X1_491 ( .gnd(gnd), .vdd(vdd), .A(_2305__bF_buf3), .B(_2304__bF_buf3), .Y(_2306_) );
XNOR2X1 XNOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_2306__bF_buf3), .B(micro_hash_ucr_Wx_2_), .Y(_2307_) );
NOR2X1 NOR2X1_492 ( .gnd(gnd), .vdd(vdd), .A(_2307_), .B(_2300_), .Y(_2308_) );
AND2X2 AND2X2_208 ( .gnd(gnd), .vdd(vdd), .A(_2300_), .B(_2307_), .Y(_2309_) );
OAI21X1 OAI21X1_596 ( .gnd(gnd), .vdd(vdd), .A(_2309_), .B(_2308_), .C(micro_hash_ucr_pipe8), .Y(_2310_) );
OAI21X1 OAI21X1_597 ( .gnd(gnd), .vdd(vdd), .A(_2091_), .B(_1966_), .C(_2092_), .Y(_2311_) );
XNOR2X1 XNOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(_2306__bF_buf2), .B(micro_hash_ucr_Wx_10_), .Y(_2312_) );
XNOR2X1 XNOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_2311_), .B(_2312_), .Y(_2313_) );
NAND2X1 NAND2X1_308 ( .gnd(gnd), .vdd(vdd), .A(_1174_), .B(_937_), .Y(_2314_) );
OAI21X1 OAI21X1_598 ( .gnd(gnd), .vdd(vdd), .A(H_18_), .B(_937_), .C(_2314_), .Y(_2315_) );
AOI21X1 AOI21X1_407 ( .gnd(gnd), .vdd(vdd), .A(_938_), .B(_2315_), .C(micro_hash_ucr_pipe10), .Y(_2316_) );
AOI22X1 AOI22X1_28 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe10), .B(_2313_), .C(_2310_), .D(_2316_), .Y(_2317_) );
OAI21X1 OAI21X1_599 ( .gnd(gnd), .vdd(vdd), .A(_2109_), .B(_2108_), .C(_2111_), .Y(_2318_) );
INVX1 INVX1_135 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_18_), .Y(_2319_) );
OAI21X1 OAI21X1_600 ( .gnd(gnd), .vdd(vdd), .A(_2304__bF_buf2), .B(_2305__bF_buf2), .C(_2319_), .Y(_2320_) );
INVX1 INVX1_136 ( .gnd(gnd), .vdd(vdd), .A(_2320_), .Y(_2321_) );
INVX8 INVX8_90 ( .gnd(gnd), .vdd(vdd), .A(_2306__bF_buf1), .Y(_2322_) );
NOR2X1 NOR2X1_493 ( .gnd(gnd), .vdd(vdd), .A(_2319_), .B(_2322__bF_buf5), .Y(_2323_) );
NOR2X1 NOR2X1_494 ( .gnd(gnd), .vdd(vdd), .A(_2321_), .B(_2323_), .Y(_2324_) );
XOR2X1 XOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_2324_), .B(_2318_), .Y(_2325_) );
AOI21X1 AOI21X1_408 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe12), .B(_2325_), .C(micro_hash_ucr_pipe14_bF_buf2), .Y(_2326_) );
OAI21X1 OAI21X1_601 ( .gnd(gnd), .vdd(vdd), .A(_2317_), .B(micro_hash_ucr_pipe12), .C(_2326_), .Y(_2327_) );
OAI21X1 OAI21X1_602 ( .gnd(gnd), .vdd(vdd), .A(_2116_), .B(_2115_), .C(_2118_), .Y(_2328_) );
INVX2 INVX2_105 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_26_), .Y(_2329_) );
XNOR2X1 XNOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_2306__bF_buf0), .B(_2329_), .Y(_2330_) );
NAND2X1 NAND2X1_309 ( .gnd(gnd), .vdd(vdd), .A(_2330_), .B(_2328_), .Y(_2331_) );
INVX1 INVX1_137 ( .gnd(gnd), .vdd(vdd), .A(_2331_), .Y(_2332_) );
NOR2X1 NOR2X1_495 ( .gnd(gnd), .vdd(vdd), .A(_2330_), .B(_2328_), .Y(_2333_) );
OAI21X1 OAI21X1_603 ( .gnd(gnd), .vdd(vdd), .A(_2332_), .B(_2333_), .C(micro_hash_ucr_pipe14_bF_buf1), .Y(_2334_) );
AOI21X1 AOI21X1_409 ( .gnd(gnd), .vdd(vdd), .A(_2334_), .B(_2327_), .C(micro_hash_ucr_pipe16_bF_buf2), .Y(_2335_) );
INVX1 INVX1_138 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_33_), .Y(_2336_) );
NAND2X1 NAND2X1_310 ( .gnd(gnd), .vdd(vdd), .A(_1963_), .B(_2122_), .Y(_2337_) );
OAI21X1 OAI21X1_604 ( .gnd(gnd), .vdd(vdd), .A(_2336_), .B(_2089__bF_buf2), .C(_2337_), .Y(_2338_) );
INVX2 INVX2_106 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_34_), .Y(_2339_) );
OAI21X1 OAI21X1_605 ( .gnd(gnd), .vdd(vdd), .A(_2304__bF_buf1), .B(_2305__bF_buf1), .C(_2339_), .Y(_2340_) );
NOR2X1 NOR2X1_496 ( .gnd(gnd), .vdd(vdd), .A(_2339_), .B(_2322__bF_buf4), .Y(_2341_) );
INVX1 INVX1_139 ( .gnd(gnd), .vdd(vdd), .A(_2341_), .Y(_2342_) );
NAND2X1 NAND2X1_311 ( .gnd(gnd), .vdd(vdd), .A(_2340_), .B(_2342_), .Y(_2343_) );
XNOR2X1 XNOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_2343_), .B(_2338_), .Y(_2344_) );
OAI21X1 OAI21X1_606 ( .gnd(gnd), .vdd(vdd), .A(_2344_), .B(_930__bF_buf0), .C(_925__bF_buf1), .Y(_2345_) );
INVX1 INVX1_140 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_41_), .Y(_2346_) );
OAI21X1 OAI21X1_607 ( .gnd(gnd), .vdd(vdd), .A(_2346_), .B(_2089__bF_buf1), .C(_2126_), .Y(_2347_) );
INVX2 INVX2_107 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_42_), .Y(_2348_) );
XNOR2X1 XNOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(_2306__bF_buf3), .B(_2348_), .Y(_2349_) );
XOR2X1 XOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_2347_), .B(_2349_), .Y(_2350_) );
AOI21X1 AOI21X1_410 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe18_bF_buf4), .B(_2350_), .C(micro_hash_ucr_pipe20_bF_buf2), .Y(_2351_) );
OAI21X1 OAI21X1_608 ( .gnd(gnd), .vdd(vdd), .A(_2335_), .B(_2345_), .C(_2351_), .Y(_2352_) );
OR2X2 OR2X2_31 ( .gnd(gnd), .vdd(vdd), .A(_2133_), .B(_2131_), .Y(_2353_) );
INVX1 INVX1_141 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_50_), .Y(_2354_) );
OAI21X1 OAI21X1_609 ( .gnd(gnd), .vdd(vdd), .A(_2304__bF_buf0), .B(_2305__bF_buf0), .C(_2354_), .Y(_2355_) );
NOR2X1 NOR2X1_497 ( .gnd(gnd), .vdd(vdd), .A(_2354_), .B(_2322__bF_buf3), .Y(_2356_) );
INVX1 INVX1_142 ( .gnd(gnd), .vdd(vdd), .A(_2356_), .Y(_2357_) );
NAND2X1 NAND2X1_312 ( .gnd(gnd), .vdd(vdd), .A(_2355_), .B(_2357_), .Y(_2358_) );
XOR2X1 XOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_2353_), .B(_2358_), .Y(_2359_) );
AOI21X1 AOI21X1_411 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe20_bF_buf1), .B(_2359_), .C(micro_hash_ucr_pipe22_bF_buf2), .Y(_2360_) );
NAND2X1 NAND2X1_313 ( .gnd(gnd), .vdd(vdd), .A(_2360_), .B(_2352_), .Y(_2361_) );
OAI21X1 OAI21X1_610 ( .gnd(gnd), .vdd(vdd), .A(_2304__bF_buf3), .B(_2305__bF_buf3), .C(_813_), .Y(_2362_) );
INVX1 INVX1_143 ( .gnd(gnd), .vdd(vdd), .A(_2362_), .Y(_2363_) );
NOR2X1 NOR2X1_498 ( .gnd(gnd), .vdd(vdd), .A(_813_), .B(_2322__bF_buf2), .Y(_2364_) );
NOR2X1 NOR2X1_499 ( .gnd(gnd), .vdd(vdd), .A(_2363_), .B(_2364_), .Y(_2365_) );
OAI21X1 OAI21X1_611 ( .gnd(gnd), .vdd(vdd), .A(_2140_), .B(_2138_), .C(_2365_), .Y(_2366_) );
NOR2X1 NOR2X1_500 ( .gnd(gnd), .vdd(vdd), .A(_2138_), .B(_2140_), .Y(_2367_) );
OAI21X1 OAI21X1_612 ( .gnd(gnd), .vdd(vdd), .A(_2363_), .B(_2364_), .C(_2367_), .Y(_2368_) );
NAND2X1 NAND2X1_314 ( .gnd(gnd), .vdd(vdd), .A(_2366_), .B(_2368_), .Y(_2369_) );
OAI21X1 OAI21X1_613 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf3), .B(_2369_), .C(_2361_), .Y(_2370_) );
OAI21X1 OAI21X1_614 ( .gnd(gnd), .vdd(vdd), .A(_856_), .B(_2089__bF_buf0), .C(_2147_), .Y(_2371_) );
XNOR2X1 XNOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_2306__bF_buf2), .B(_859_), .Y(_2372_) );
NAND2X1 NAND2X1_315 ( .gnd(gnd), .vdd(vdd), .A(_2372_), .B(_2371_), .Y(_2373_) );
INVX1 INVX1_144 ( .gnd(gnd), .vdd(vdd), .A(_2373_), .Y(_2374_) );
NOR2X1 NOR2X1_501 ( .gnd(gnd), .vdd(vdd), .A(_2372_), .B(_2371_), .Y(_2375_) );
OAI21X1 OAI21X1_615 ( .gnd(gnd), .vdd(vdd), .A(_2374_), .B(_2375_), .C(micro_hash_ucr_pipe24_bF_buf0), .Y(_2376_) );
OAI21X1 OAI21X1_616 ( .gnd(gnd), .vdd(vdd), .A(_2370_), .B(micro_hash_ucr_pipe24_bF_buf4), .C(_2376_), .Y(_2377_) );
NOR2X1 NOR2X1_502 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe26_bF_buf1), .B(_2377_), .Y(_2378_) );
OAI21X1 OAI21X1_617 ( .gnd(gnd), .vdd(vdd), .A(_832_), .B(_2089__bF_buf5), .C(_2153_), .Y(_2379_) );
XNOR2X1 XNOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(_2306__bF_buf1), .B(_835_), .Y(_2380_) );
NOR2X1 NOR2X1_503 ( .gnd(gnd), .vdd(vdd), .A(_2380_), .B(_2379_), .Y(_2381_) );
NAND2X1 NAND2X1_316 ( .gnd(gnd), .vdd(vdd), .A(_2380_), .B(_2379_), .Y(_2382_) );
NAND2X1 NAND2X1_317 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe26_bF_buf0), .B(_2382_), .Y(_2383_) );
OAI21X1 OAI21X1_618 ( .gnd(gnd), .vdd(vdd), .A(_2383_), .B(_2381_), .C(_918__bF_buf1), .Y(_2384_) );
OAI21X1 OAI21X1_619 ( .gnd(gnd), .vdd(vdd), .A(_743_), .B(_2089__bF_buf4), .C(_2160_), .Y(_2385_) );
OAI21X1 OAI21X1_620 ( .gnd(gnd), .vdd(vdd), .A(_2304__bF_buf2), .B(_2305__bF_buf2), .C(_746_), .Y(_2386_) );
NOR2X1 NOR2X1_504 ( .gnd(gnd), .vdd(vdd), .A(_746_), .B(_2322__bF_buf1), .Y(_2387_) );
INVX1 INVX1_145 ( .gnd(gnd), .vdd(vdd), .A(_2387_), .Y(_2388_) );
NAND2X1 NAND2X1_318 ( .gnd(gnd), .vdd(vdd), .A(_2386_), .B(_2388_), .Y(_2389_) );
XOR2X1 XOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_2389_), .B(_2385_), .Y(_2390_) );
AOI21X1 AOI21X1_412 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe28_bF_buf2), .B(_2390_), .C(micro_hash_ucr_pipe30_bF_buf3), .Y(_2391_) );
OAI21X1 OAI21X1_621 ( .gnd(gnd), .vdd(vdd), .A(_2378_), .B(_2384_), .C(_2391_), .Y(_2392_) );
OAI21X1 OAI21X1_622 ( .gnd(gnd), .vdd(vdd), .A(_2304__bF_buf1), .B(_2305__bF_buf1), .C(_786_), .Y(_2393_) );
INVX1 INVX1_146 ( .gnd(gnd), .vdd(vdd), .A(_2393_), .Y(_2394_) );
NOR2X1 NOR2X1_505 ( .gnd(gnd), .vdd(vdd), .A(_786_), .B(_2322__bF_buf0), .Y(_2395_) );
NOR2X1 NOR2X1_506 ( .gnd(gnd), .vdd(vdd), .A(_2394_), .B(_2395_), .Y(_2396_) );
OAI21X1 OAI21X1_623 ( .gnd(gnd), .vdd(vdd), .A(_2167_), .B(_2165_), .C(_2396_), .Y(_2397_) );
NOR2X1 NOR2X1_507 ( .gnd(gnd), .vdd(vdd), .A(_2165_), .B(_2167_), .Y(_2398_) );
OAI21X1 OAI21X1_624 ( .gnd(gnd), .vdd(vdd), .A(_2394_), .B(_2395_), .C(_2398_), .Y(_2399_) );
NAND2X1 NAND2X1_319 ( .gnd(gnd), .vdd(vdd), .A(_2397_), .B(_2399_), .Y(_2400_) );
OAI21X1 OAI21X1_625 ( .gnd(gnd), .vdd(vdd), .A(_913__bF_buf4), .B(_2400_), .C(_2392_), .Y(_2401_) );
NAND2X1 NAND2X1_320 ( .gnd(gnd), .vdd(vdd), .A(_2012_), .B(_2171_), .Y(_2402_) );
OAI21X1 OAI21X1_626 ( .gnd(gnd), .vdd(vdd), .A(_644_), .B(_2089__bF_buf3), .C(_2402_), .Y(_2403_) );
OAI21X1 OAI21X1_627 ( .gnd(gnd), .vdd(vdd), .A(_2304__bF_buf0), .B(_2305__bF_buf0), .C(_648_), .Y(_2404_) );
NOR2X1 NOR2X1_508 ( .gnd(gnd), .vdd(vdd), .A(_648_), .B(_2322__bF_buf5), .Y(_2405_) );
INVX1 INVX1_147 ( .gnd(gnd), .vdd(vdd), .A(_2405_), .Y(_2406_) );
NAND2X1 NAND2X1_321 ( .gnd(gnd), .vdd(vdd), .A(_2404_), .B(_2406_), .Y(_2407_) );
XNOR2X1 XNOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_2407_), .B(_2403_), .Y(_2408_) );
MUX2X1 MUX2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_2401_), .B(_2408_), .S(_914__bF_buf0), .Y(_2409_) );
AOI21X1 AOI21X1_413 ( .gnd(gnd), .vdd(vdd), .A(_2015_), .B(_2178_), .C(_2177_), .Y(_2410_) );
OAI21X1 OAI21X1_628 ( .gnd(gnd), .vdd(vdd), .A(_2304__bF_buf3), .B(_2305__bF_buf3), .C(_676_), .Y(_2411_) );
INVX1 INVX1_148 ( .gnd(gnd), .vdd(vdd), .A(_2411_), .Y(_2412_) );
NOR2X1 NOR2X1_509 ( .gnd(gnd), .vdd(vdd), .A(_676_), .B(_2322__bF_buf4), .Y(_2413_) );
OAI21X1 OAI21X1_629 ( .gnd(gnd), .vdd(vdd), .A(_2413_), .B(_2412_), .C(_2410_), .Y(_2414_) );
INVX1 INVX1_149 ( .gnd(gnd), .vdd(vdd), .A(_2410_), .Y(_2415_) );
NOR2X1 NOR2X1_510 ( .gnd(gnd), .vdd(vdd), .A(_2412_), .B(_2413_), .Y(_2416_) );
NAND2X1 NAND2X1_322 ( .gnd(gnd), .vdd(vdd), .A(_2416_), .B(_2415_), .Y(_2417_) );
AOI21X1 AOI21X1_414 ( .gnd(gnd), .vdd(vdd), .A(_2414_), .B(_2417_), .C(_912__bF_buf2), .Y(_2418_) );
AOI21X1 AOI21X1_415 ( .gnd(gnd), .vdd(vdd), .A(_912__bF_buf1), .B(_2409_), .C(_2418_), .Y(_2419_) );
OAI21X1 OAI21X1_630 ( .gnd(gnd), .vdd(vdd), .A(_506_), .B(_2089__bF_buf2), .C(_2185_), .Y(_2420_) );
OAI21X1 OAI21X1_631 ( .gnd(gnd), .vdd(vdd), .A(_2304__bF_buf2), .B(_2305__bF_buf2), .C(_510_), .Y(_2421_) );
NOR2X1 NOR2X1_511 ( .gnd(gnd), .vdd(vdd), .A(_510_), .B(_2322__bF_buf3), .Y(_2422_) );
INVX1 INVX1_150 ( .gnd(gnd), .vdd(vdd), .A(_2422_), .Y(_2423_) );
NAND2X1 NAND2X1_323 ( .gnd(gnd), .vdd(vdd), .A(_2421_), .B(_2423_), .Y(_2424_) );
XOR2X1 XOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_2424_), .B(_2420_), .Y(_2425_) );
AOI21X1 AOI21X1_416 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe36_bF_buf3), .B(_2425_), .C(micro_hash_ucr_pipe38_bF_buf1), .Y(_2426_) );
OAI21X1 OAI21X1_632 ( .gnd(gnd), .vdd(vdd), .A(_2419_), .B(micro_hash_ucr_pipe36_bF_buf2), .C(_2426_), .Y(_2427_) );
AOI21X1 AOI21X1_417 ( .gnd(gnd), .vdd(vdd), .A(_2021_), .B(_2190_), .C(_2189_), .Y(_2428_) );
OAI21X1 OAI21X1_633 ( .gnd(gnd), .vdd(vdd), .A(_2304__bF_buf1), .B(_2305__bF_buf1), .C(_566_), .Y(_2429_) );
INVX1 INVX1_151 ( .gnd(gnd), .vdd(vdd), .A(_2429_), .Y(_2430_) );
NOR2X1 NOR2X1_512 ( .gnd(gnd), .vdd(vdd), .A(_566_), .B(_2322__bF_buf2), .Y(_2431_) );
NOR2X1 NOR2X1_513 ( .gnd(gnd), .vdd(vdd), .A(_2430_), .B(_2431_), .Y(_2432_) );
INVX1 INVX1_152 ( .gnd(gnd), .vdd(vdd), .A(_2432_), .Y(_2433_) );
NOR2X1 NOR2X1_514 ( .gnd(gnd), .vdd(vdd), .A(_2433_), .B(_2428_), .Y(_2434_) );
INVX1 INVX1_153 ( .gnd(gnd), .vdd(vdd), .A(_2434_), .Y(_2435_) );
OAI21X1 OAI21X1_634 ( .gnd(gnd), .vdd(vdd), .A(_2431_), .B(_2430_), .C(_2428_), .Y(_2436_) );
NAND2X1 NAND2X1_324 ( .gnd(gnd), .vdd(vdd), .A(_2436_), .B(_2435_), .Y(_2437_) );
OAI21X1 OAI21X1_635 ( .gnd(gnd), .vdd(vdd), .A(_908__bF_buf2), .B(_2437_), .C(_2427_), .Y(_2438_) );
NOR2X1 NOR2X1_515 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe40_bF_buf1), .B(_2438_), .Y(_2439_) );
NAND2X1 NAND2X1_325 ( .gnd(gnd), .vdd(vdd), .A(_2025_), .B(_2193_), .Y(_2440_) );
OAI21X1 OAI21X1_636 ( .gnd(gnd), .vdd(vdd), .A(_534_), .B(_2089__bF_buf1), .C(_2440_), .Y(_2441_) );
OAI21X1 OAI21X1_637 ( .gnd(gnd), .vdd(vdd), .A(_2304__bF_buf0), .B(_2305__bF_buf0), .C(_538_), .Y(_2442_) );
NOR2X1 NOR2X1_516 ( .gnd(gnd), .vdd(vdd), .A(_538_), .B(_2322__bF_buf1), .Y(_2443_) );
INVX1 INVX1_154 ( .gnd(gnd), .vdd(vdd), .A(_2443_), .Y(_2444_) );
NAND2X1 NAND2X1_326 ( .gnd(gnd), .vdd(vdd), .A(_2442_), .B(_2444_), .Y(_2445_) );
XNOR2X1 XNOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(_2445_), .B(_2441_), .Y(_2446_) );
OAI21X1 OAI21X1_638 ( .gnd(gnd), .vdd(vdd), .A(_2446_), .B(_906__bF_buf1), .C(_901__bF_buf3), .Y(_2447_) );
XNOR2X1 XNOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(_2306__bF_buf0), .B(_787_), .Y(_2448_) );
OAI21X1 OAI21X1_639 ( .gnd(gnd), .vdd(vdd), .A(_2203_), .B(_2200_), .C(_2448_), .Y(_2449_) );
INVX1 INVX1_155 ( .gnd(gnd), .vdd(vdd), .A(_2449_), .Y(_2450_) );
OAI21X1 OAI21X1_640 ( .gnd(gnd), .vdd(vdd), .A(_2198_), .B(_2197_), .C(_2201_), .Y(_2451_) );
OAI21X1 OAI21X1_641 ( .gnd(gnd), .vdd(vdd), .A(_2451_), .B(_2448_), .C(micro_hash_ucr_pipe42_bF_buf0), .Y(_2452_) );
OAI22X1 OAI22X1_48 ( .gnd(gnd), .vdd(vdd), .A(_2450_), .B(_2452_), .C(_2439_), .D(_2447_), .Y(_2453_) );
OAI21X1 OAI21X1_642 ( .gnd(gnd), .vdd(vdd), .A(_615_), .B(_2089__bF_buf0), .C(_2210_), .Y(_2454_) );
XNOR2X1 XNOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(_2306__bF_buf3), .B(_619_), .Y(_2455_) );
NOR2X1 NOR2X1_517 ( .gnd(gnd), .vdd(vdd), .A(_2455_), .B(_2454_), .Y(_2456_) );
OAI21X1 OAI21X1_643 ( .gnd(gnd), .vdd(vdd), .A(_2211_), .B(_2208_), .C(_2455_), .Y(_2457_) );
INVX1 INVX1_156 ( .gnd(gnd), .vdd(vdd), .A(_2457_), .Y(_2458_) );
OAI21X1 OAI21X1_644 ( .gnd(gnd), .vdd(vdd), .A(_2458_), .B(_2456_), .C(micro_hash_ucr_pipe44), .Y(_2459_) );
OAI21X1 OAI21X1_645 ( .gnd(gnd), .vdd(vdd), .A(_2453_), .B(micro_hash_ucr_pipe44), .C(_2459_), .Y(_2460_) );
OAI21X1 OAI21X1_646 ( .gnd(gnd), .vdd(vdd), .A(_2215_), .B(_2036_), .C(_2217_), .Y(_2461_) );
OAI21X1 OAI21X1_647 ( .gnd(gnd), .vdd(vdd), .A(_2304__bF_buf3), .B(_2305__bF_buf3), .C(_677_), .Y(_2462_) );
NOR2X1 NOR2X1_518 ( .gnd(gnd), .vdd(vdd), .A(_677_), .B(_2322__bF_buf0), .Y(_2463_) );
INVX1 INVX1_157 ( .gnd(gnd), .vdd(vdd), .A(_2463_), .Y(_2464_) );
NAND2X1 NAND2X1_327 ( .gnd(gnd), .vdd(vdd), .A(_2462_), .B(_2464_), .Y(_2465_) );
XNOR2X1 XNOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_2465_), .B(_2461_), .Y(_2466_) );
OAI21X1 OAI21X1_648 ( .gnd(gnd), .vdd(vdd), .A(_2466_), .B(_900__bF_buf1), .C(_895__bF_buf2), .Y(_2467_) );
AOI21X1 AOI21X1_418 ( .gnd(gnd), .vdd(vdd), .A(_900__bF_buf0), .B(_2460_), .C(_2467_), .Y(_2468_) );
XNOR2X1 XNOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(_2306__bF_buf2), .B(_725_), .Y(_2469_) );
OAI21X1 OAI21X1_649 ( .gnd(gnd), .vdd(vdd), .A(_2225_), .B(_2222_), .C(_2469_), .Y(_2470_) );
INVX1 INVX1_158 ( .gnd(gnd), .vdd(vdd), .A(_2470_), .Y(_2471_) );
OAI21X1 OAI21X1_650 ( .gnd(gnd), .vdd(vdd), .A(_722_), .B(_2089__bF_buf5), .C(_2224_), .Y(_2472_) );
OAI21X1 OAI21X1_651 ( .gnd(gnd), .vdd(vdd), .A(_2472_), .B(_2469_), .C(micro_hash_ucr_pipe48_bF_buf1), .Y(_2473_) );
OAI21X1 OAI21X1_652 ( .gnd(gnd), .vdd(vdd), .A(_2471_), .B(_2473_), .C(_896__bF_buf1), .Y(_2474_) );
XNOR2X1 XNOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(_2306__bF_buf1), .B(_702_), .Y(_2475_) );
OAI21X1 OAI21X1_653 ( .gnd(gnd), .vdd(vdd), .A(_2232_), .B(_2229_), .C(_2475_), .Y(_2476_) );
INVX1 INVX1_159 ( .gnd(gnd), .vdd(vdd), .A(_2476_), .Y(_2477_) );
OAI21X1 OAI21X1_654 ( .gnd(gnd), .vdd(vdd), .A(_699_), .B(_2089__bF_buf4), .C(_2231_), .Y(_2478_) );
NOR2X1 NOR2X1_519 ( .gnd(gnd), .vdd(vdd), .A(_2475_), .B(_2478_), .Y(_2479_) );
OAI21X1 OAI21X1_655 ( .gnd(gnd), .vdd(vdd), .A(_2477_), .B(_2479_), .C(micro_hash_ucr_pipe50_bF_buf1), .Y(_2480_) );
OAI21X1 OAI21X1_656 ( .gnd(gnd), .vdd(vdd), .A(_2468_), .B(_2474_), .C(_2480_), .Y(_2481_) );
XNOR2X1 XNOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_2306__bF_buf0), .B(_593_), .Y(_2482_) );
OAI21X1 OAI21X1_657 ( .gnd(gnd), .vdd(vdd), .A(_2241_), .B(_2237_), .C(_2482_), .Y(_2483_) );
INVX1 INVX1_160 ( .gnd(gnd), .vdd(vdd), .A(_2483_), .Y(_2484_) );
OAI21X1 OAI21X1_658 ( .gnd(gnd), .vdd(vdd), .A(_590_), .B(_2089__bF_buf3), .C(_2240_), .Y(_2485_) );
OAI21X1 OAI21X1_659 ( .gnd(gnd), .vdd(vdd), .A(_2485_), .B(_2482_), .C(micro_hash_ucr_pipe52_bF_buf2), .Y(_2486_) );
OAI22X1 OAI22X1_49 ( .gnd(gnd), .vdd(vdd), .A(_2484_), .B(_2486_), .C(_2481_), .D(micro_hash_ucr_pipe52_bF_buf1), .Y(_2487_) );
NOR2X1 NOR2X1_520 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe54_bF_buf1), .B(_2487_), .Y(_2488_) );
NAND2X1 NAND2X1_328 ( .gnd(gnd), .vdd(vdd), .A(_2054_), .B(_2245_), .Y(_2489_) );
OAI21X1 OAI21X1_660 ( .gnd(gnd), .vdd(vdd), .A(_645_), .B(_2089__bF_buf2), .C(_2489_), .Y(_2490_) );
OAI21X1 OAI21X1_661 ( .gnd(gnd), .vdd(vdd), .A(_2304__bF_buf2), .B(_2305__bF_buf2), .C(_649_), .Y(_2491_) );
NOR2X1 NOR2X1_521 ( .gnd(gnd), .vdd(vdd), .A(_649_), .B(_2322__bF_buf5), .Y(_2492_) );
INVX1 INVX1_161 ( .gnd(gnd), .vdd(vdd), .A(_2492_), .Y(_2493_) );
NAND2X1 NAND2X1_329 ( .gnd(gnd), .vdd(vdd), .A(_2491_), .B(_2493_), .Y(_2494_) );
XNOR2X1 XNOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(_2494_), .B(_2490_), .Y(_2495_) );
OAI21X1 OAI21X1_662 ( .gnd(gnd), .vdd(vdd), .A(_2495_), .B(_889__bF_buf1), .C(_890__bF_buf3), .Y(_2496_) );
XNOR2X1 XNOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(_2306__bF_buf3), .B(_620_), .Y(_2497_) );
OAI21X1 OAI21X1_663 ( .gnd(gnd), .vdd(vdd), .A(_2252_), .B(_2249_), .C(_2497_), .Y(_2498_) );
INVX1 INVX1_162 ( .gnd(gnd), .vdd(vdd), .A(_2498_), .Y(_2499_) );
OAI21X1 OAI21X1_664 ( .gnd(gnd), .vdd(vdd), .A(_616_), .B(_2089__bF_buf1), .C(_2251_), .Y(_2500_) );
OAI21X1 OAI21X1_665 ( .gnd(gnd), .vdd(vdd), .A(_2500_), .B(_2497_), .C(micro_hash_ucr_pipe56_bF_buf0), .Y(_2501_) );
OAI22X1 OAI22X1_50 ( .gnd(gnd), .vdd(vdd), .A(_2499_), .B(_2501_), .C(_2488_), .D(_2496_), .Y(_2502_) );
OAI21X1 OAI21X1_666 ( .gnd(gnd), .vdd(vdd), .A(_507_), .B(_2089__bF_buf0), .C(_2259_), .Y(_2503_) );
XNOR2X1 XNOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(_2306__bF_buf2), .B(_511_), .Y(_2504_) );
NOR2X1 NOR2X1_522 ( .gnd(gnd), .vdd(vdd), .A(_2504_), .B(_2503_), .Y(_2505_) );
NAND2X1 NAND2X1_330 ( .gnd(gnd), .vdd(vdd), .A(_2504_), .B(_2503_), .Y(_2506_) );
INVX1 INVX1_163 ( .gnd(gnd), .vdd(vdd), .A(_2506_), .Y(_2507_) );
OAI21X1 OAI21X1_667 ( .gnd(gnd), .vdd(vdd), .A(_2507_), .B(_2505_), .C(micro_hash_ucr_pipe58_bF_buf4), .Y(_2508_) );
OAI21X1 OAI21X1_668 ( .gnd(gnd), .vdd(vdd), .A(_2502_), .B(micro_hash_ucr_pipe58_bF_buf3), .C(_2508_), .Y(_2509_) );
OAI21X1 OAI21X1_669 ( .gnd(gnd), .vdd(vdd), .A(_2264_), .B(_2263_), .C(_2266_), .Y(_2510_) );
OAI21X1 OAI21X1_670 ( .gnd(gnd), .vdd(vdd), .A(_2304__bF_buf1), .B(_2305__bF_buf1), .C(_567_), .Y(_2511_) );
NOR2X1 NOR2X1_523 ( .gnd(gnd), .vdd(vdd), .A(_567_), .B(_2322__bF_buf4), .Y(_2512_) );
INVX1 INVX1_164 ( .gnd(gnd), .vdd(vdd), .A(_2512_), .Y(_2513_) );
NAND2X1 NAND2X1_331 ( .gnd(gnd), .vdd(vdd), .A(_2511_), .B(_2513_), .Y(_2514_) );
XOR2X1 XOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(_2514_), .B(_2510_), .Y(_2515_) );
MUX2X1 MUX2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_2509_), .B(_2515_), .S(_883__bF_buf3), .Y(_2516_) );
XNOR2X1 XNOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(_2306__bF_buf1), .B(_539_), .Y(_2517_) );
OAI21X1 OAI21X1_671 ( .gnd(gnd), .vdd(vdd), .A(_2274_), .B(_2271_), .C(_2517_), .Y(_2518_) );
INVX1 INVX1_165 ( .gnd(gnd), .vdd(vdd), .A(_2518_), .Y(_2519_) );
OAI21X1 OAI21X1_672 ( .gnd(gnd), .vdd(vdd), .A(_535_), .B(_2089__bF_buf5), .C(_2273_), .Y(_2520_) );
NOR2X1 NOR2X1_524 ( .gnd(gnd), .vdd(vdd), .A(_2517_), .B(_2520_), .Y(_2521_) );
OAI21X1 OAI21X1_673 ( .gnd(gnd), .vdd(vdd), .A(_2519_), .B(_2521_), .C(micro_hash_ucr_pipe62_bF_buf2), .Y(_2522_) );
OAI21X1 OAI21X1_674 ( .gnd(gnd), .vdd(vdd), .A(_2516_), .B(micro_hash_ucr_pipe62_bF_buf1), .C(_2522_), .Y(_2523_) );
INVX1 INVX1_166 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_225_), .Y(_2524_) );
NAND2X1 NAND2X1_332 ( .gnd(gnd), .vdd(vdd), .A(_2071_), .B(_2278_), .Y(_2525_) );
OAI21X1 OAI21X1_675 ( .gnd(gnd), .vdd(vdd), .A(_2524_), .B(_2089__bF_buf4), .C(_2525_), .Y(_2526_) );
INVX2 INVX2_108 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_226_), .Y(_2527_) );
OAI21X1 OAI21X1_676 ( .gnd(gnd), .vdd(vdd), .A(_2304__bF_buf0), .B(_2305__bF_buf0), .C(_2527_), .Y(_2528_) );
NOR2X1 NOR2X1_525 ( .gnd(gnd), .vdd(vdd), .A(_2527_), .B(_2322__bF_buf3), .Y(_2529_) );
INVX1 INVX1_167 ( .gnd(gnd), .vdd(vdd), .A(_2529_), .Y(_2530_) );
NAND2X1 NAND2X1_333 ( .gnd(gnd), .vdd(vdd), .A(_2528_), .B(_2530_), .Y(_2531_) );
XOR2X1 XOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_2531_), .B(_2526_), .Y(_2532_) );
MUX2X1 MUX2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_2523_), .B(_2532_), .S(_882__bF_buf0), .Y(_2533_) );
OAI21X1 OAI21X1_677 ( .gnd(gnd), .vdd(vdd), .A(_2282_), .B(_1959_), .C(_2284_), .Y(_2534_) );
INVX2 INVX2_109 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_234_), .Y(_2535_) );
XNOR2X1 XNOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(_2306__bF_buf0), .B(_2535_), .Y(_2536_) );
NOR2X1 NOR2X1_526 ( .gnd(gnd), .vdd(vdd), .A(_2536_), .B(_2534_), .Y(_2537_) );
NAND2X1 NAND2X1_334 ( .gnd(gnd), .vdd(vdd), .A(_2536_), .B(_2534_), .Y(_2538_) );
NAND2X1 NAND2X1_335 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe66_bF_buf2), .B(_2538_), .Y(_2539_) );
OAI21X1 OAI21X1_678 ( .gnd(gnd), .vdd(vdd), .A(_2539_), .B(_2537_), .C(_878__bF_buf3), .Y(_2540_) );
AOI21X1 AOI21X1_419 ( .gnd(gnd), .vdd(vdd), .A(_877__bF_buf1), .B(_2533_), .C(_2540_), .Y(_2541_) );
INVX1 INVX1_168 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_241_), .Y(_2542_) );
NAND2X1 NAND2X1_336 ( .gnd(gnd), .vdd(vdd), .A(_2077_), .B(_2290_), .Y(_2543_) );
OAI21X1 OAI21X1_679 ( .gnd(gnd), .vdd(vdd), .A(_2542_), .B(_2089__bF_buf3), .C(_2543_), .Y(_2544_) );
INVX2 INVX2_110 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_242_), .Y(_2545_) );
OAI21X1 OAI21X1_680 ( .gnd(gnd), .vdd(vdd), .A(_2304__bF_buf3), .B(_2305__bF_buf3), .C(_2545_), .Y(_2546_) );
NOR2X1 NOR2X1_527 ( .gnd(gnd), .vdd(vdd), .A(_2545_), .B(_2322__bF_buf2), .Y(_2547_) );
INVX1 INVX1_169 ( .gnd(gnd), .vdd(vdd), .A(_2547_), .Y(_2548_) );
NAND2X1 NAND2X1_337 ( .gnd(gnd), .vdd(vdd), .A(_2546_), .B(_2548_), .Y(_2549_) );
XNOR2X1 XNOR2X1_61 ( .gnd(gnd), .vdd(vdd), .A(_2549_), .B(_2544_), .Y(_2550_) );
OAI21X1 OAI21X1_681 ( .gnd(gnd), .vdd(vdd), .A(_2550_), .B(_878__bF_buf2), .C(_1949_), .Y(_2551_) );
NAND2X1 NAND2X1_338 ( .gnd(gnd), .vdd(vdd), .A(_2293_), .B(_2297_), .Y(_2552_) );
OAI21X1 OAI21X1_682 ( .gnd(gnd), .vdd(vdd), .A(_2295_), .B(_2089__bF_buf2), .C(_2552_), .Y(_2553_) );
INVX1 INVX1_170 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_250_), .Y(_2554_) );
OAI21X1 OAI21X1_683 ( .gnd(gnd), .vdd(vdd), .A(_2304__bF_buf2), .B(_2305__bF_buf2), .C(_2554_), .Y(_2555_) );
INVX1 INVX1_171 ( .gnd(gnd), .vdd(vdd), .A(_2555_), .Y(_2556_) );
NOR2X1 NOR2X1_528 ( .gnd(gnd), .vdd(vdd), .A(_2554_), .B(_2322__bF_buf1), .Y(_2557_) );
NOR2X1 NOR2X1_529 ( .gnd(gnd), .vdd(vdd), .A(_2556_), .B(_2557_), .Y(_2558_) );
AND2X2 AND2X2_209 ( .gnd(gnd), .vdd(vdd), .A(_2553_), .B(_2558_), .Y(_2559_) );
OAI21X1 OAI21X1_684 ( .gnd(gnd), .vdd(vdd), .A(_2553_), .B(_2558_), .C(_369_), .Y(_2560_) );
OAI22X1 OAI22X1_51 ( .gnd(gnd), .vdd(vdd), .A(_2559_), .B(_2560_), .C(_2541_), .D(_2551_), .Y(_299__2_) );
NAND2X1 NAND2X1_339 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_2_), .B(_2306__bF_buf3), .Y(_2561_) );
OAI21X1 OAI21X1_685 ( .gnd(gnd), .vdd(vdd), .A(_2300_), .B(_2307_), .C(_2561_), .Y(_2562_) );
INVX1 INVX1_172 ( .gnd(gnd), .vdd(vdd), .A(_2562_), .Y(_2563_) );
INVX1 INVX1_173 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_3_), .Y(_2564_) );
INVX1 INVX1_174 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_k_2_), .Y(_2565_) );
INVX1 INVX1_175 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_x_2_), .Y(_2566_) );
OAI21X1 OAI21X1_686 ( .gnd(gnd), .vdd(vdd), .A(_2565_), .B(_2566_), .C(_2303_), .Y(_2567_) );
XOR2X1 XOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_k_3_), .B(micro_hash_ucr_x_3_), .Y(_2568_) );
AND2X2 AND2X2_210 ( .gnd(gnd), .vdd(vdd), .A(_2567_), .B(_2568_), .Y(_2569_) );
NOR2X1 NOR2X1_530 ( .gnd(gnd), .vdd(vdd), .A(_2568_), .B(_2567_), .Y(_2570_) );
OAI21X1 OAI21X1_687 ( .gnd(gnd), .vdd(vdd), .A(_2569__bF_buf4), .B(_2570__bF_buf4), .C(_2564_), .Y(_2571_) );
INVX1 INVX1_176 ( .gnd(gnd), .vdd(vdd), .A(_2571_), .Y(_2572_) );
NOR2X1 NOR2X1_531 ( .gnd(gnd), .vdd(vdd), .A(_2570__bF_buf3), .B(_2569__bF_buf3), .Y(_2573_) );
INVX8 INVX8_91 ( .gnd(gnd), .vdd(vdd), .A(_2573_), .Y(_2574_) );
NOR2X1 NOR2X1_532 ( .gnd(gnd), .vdd(vdd), .A(_2564_), .B(_2574__bF_buf4), .Y(_2575_) );
NOR2X1 NOR2X1_533 ( .gnd(gnd), .vdd(vdd), .A(_2572_), .B(_2575_), .Y(_2576_) );
OAI21X1 OAI21X1_688 ( .gnd(gnd), .vdd(vdd), .A(_2563_), .B(_2576_), .C(micro_hash_ucr_pipe8), .Y(_2577_) );
AOI21X1 AOI21X1_420 ( .gnd(gnd), .vdd(vdd), .A(_2563_), .B(_2576_), .C(_2577_), .Y(_2578_) );
NOR2X1 NOR2X1_534 ( .gnd(gnd), .vdd(vdd), .A(_4444_), .B(_937_), .Y(_2579_) );
OAI21X1 OAI21X1_689 ( .gnd(gnd), .vdd(vdd), .A(_4445_), .B(micro_hash_ucr_pipe6), .C(_938_), .Y(_2580_) );
OAI21X1 OAI21X1_690 ( .gnd(gnd), .vdd(vdd), .A(_2580_), .B(_2579_), .C(_936_), .Y(_2581_) );
INVX1 INVX1_177 ( .gnd(gnd), .vdd(vdd), .A(_2311_), .Y(_2582_) );
NAND2X1 NAND2X1_340 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_10_), .B(_2306__bF_buf2), .Y(_2583_) );
OAI21X1 OAI21X1_691 ( .gnd(gnd), .vdd(vdd), .A(_2582_), .B(_2312_), .C(_2583_), .Y(_2584_) );
INVX1 INVX1_178 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_11_), .Y(_2585_) );
OAI21X1 OAI21X1_692 ( .gnd(gnd), .vdd(vdd), .A(_2569__bF_buf2), .B(_2570__bF_buf2), .C(_2585_), .Y(_2586_) );
INVX1 INVX1_179 ( .gnd(gnd), .vdd(vdd), .A(_2586_), .Y(_2587_) );
NOR2X1 NOR2X1_535 ( .gnd(gnd), .vdd(vdd), .A(_2585_), .B(_2574__bF_buf3), .Y(_2588_) );
NOR2X1 NOR2X1_536 ( .gnd(gnd), .vdd(vdd), .A(_2587_), .B(_2588_), .Y(_2589_) );
XOR2X1 XOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_2584_), .B(_2589_), .Y(_2590_) );
AOI21X1 AOI21X1_421 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe10), .B(_2590_), .C(micro_hash_ucr_pipe12), .Y(_2591_) );
OAI21X1 OAI21X1_693 ( .gnd(gnd), .vdd(vdd), .A(_2578_), .B(_2581_), .C(_2591_), .Y(_2592_) );
AOI21X1 AOI21X1_422 ( .gnd(gnd), .vdd(vdd), .A(_2320_), .B(_2318_), .C(_2323_), .Y(_2593_) );
INVX2 INVX2_111 ( .gnd(gnd), .vdd(vdd), .A(_2593_), .Y(_2594_) );
INVX1 INVX1_180 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_19_), .Y(_2595_) );
OAI21X1 OAI21X1_694 ( .gnd(gnd), .vdd(vdd), .A(_2569__bF_buf1), .B(_2570__bF_buf1), .C(_2595_), .Y(_2596_) );
NOR2X1 NOR2X1_537 ( .gnd(gnd), .vdd(vdd), .A(_2595_), .B(_2574__bF_buf2), .Y(_2597_) );
INVX1 INVX1_181 ( .gnd(gnd), .vdd(vdd), .A(_2597_), .Y(_2598_) );
NAND2X1 NAND2X1_341 ( .gnd(gnd), .vdd(vdd), .A(_2596_), .B(_2598_), .Y(_2599_) );
AOI21X1 AOI21X1_423 ( .gnd(gnd), .vdd(vdd), .A(_2594_), .B(_2599_), .C(_931_), .Y(_2600_) );
OAI21X1 OAI21X1_695 ( .gnd(gnd), .vdd(vdd), .A(_2594_), .B(_2599_), .C(_2600_), .Y(_2601_) );
AOI21X1 AOI21X1_424 ( .gnd(gnd), .vdd(vdd), .A(_2601_), .B(_2592_), .C(micro_hash_ucr_pipe14_bF_buf0), .Y(_2602_) );
OAI21X1 OAI21X1_696 ( .gnd(gnd), .vdd(vdd), .A(_2329_), .B(_2322__bF_buf0), .C(_2331_), .Y(_2603_) );
INVX1 INVX1_182 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_27_), .Y(_2604_) );
OAI21X1 OAI21X1_697 ( .gnd(gnd), .vdd(vdd), .A(_2569__bF_buf0), .B(_2570__bF_buf0), .C(_2604_), .Y(_2605_) );
INVX1 INVX1_183 ( .gnd(gnd), .vdd(vdd), .A(_2605_), .Y(_2606_) );
NOR2X1 NOR2X1_538 ( .gnd(gnd), .vdd(vdd), .A(_2604_), .B(_2574__bF_buf1), .Y(_2607_) );
NOR2X1 NOR2X1_539 ( .gnd(gnd), .vdd(vdd), .A(_2606_), .B(_2607_), .Y(_2608_) );
XOR2X1 XOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(_2603_), .B(_2608_), .Y(_2609_) );
NOR2X1 NOR2X1_540 ( .gnd(gnd), .vdd(vdd), .A(_932_), .B(_2609_), .Y(_2610_) );
OAI21X1 OAI21X1_698 ( .gnd(gnd), .vdd(vdd), .A(_2602_), .B(_2610_), .C(_930__bF_buf4), .Y(_2611_) );
NAND3X1 NAND3X1_103 ( .gnd(gnd), .vdd(vdd), .A(_2340_), .B(_2342_), .C(_2338_), .Y(_2612_) );
OAI21X1 OAI21X1_699 ( .gnd(gnd), .vdd(vdd), .A(_2339_), .B(_2322__bF_buf5), .C(_2612_), .Y(_2613_) );
INVX1 INVX1_184 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_35_), .Y(_2614_) );
OAI21X1 OAI21X1_700 ( .gnd(gnd), .vdd(vdd), .A(_2569__bF_buf4), .B(_2570__bF_buf4), .C(_2614_), .Y(_2615_) );
NOR2X1 NOR2X1_541 ( .gnd(gnd), .vdd(vdd), .A(_2614_), .B(_2574__bF_buf0), .Y(_2616_) );
INVX1 INVX1_185 ( .gnd(gnd), .vdd(vdd), .A(_2616_), .Y(_2617_) );
NAND2X1 NAND2X1_342 ( .gnd(gnd), .vdd(vdd), .A(_2615_), .B(_2617_), .Y(_2618_) );
AOI21X1 AOI21X1_425 ( .gnd(gnd), .vdd(vdd), .A(_2618_), .B(_2613_), .C(_930__bF_buf3), .Y(_2619_) );
OAI21X1 OAI21X1_701 ( .gnd(gnd), .vdd(vdd), .A(_2613_), .B(_2618_), .C(_2619_), .Y(_2620_) );
AND2X2 AND2X2_211 ( .gnd(gnd), .vdd(vdd), .A(_2620_), .B(_925__bF_buf0), .Y(_2621_) );
NAND2X1 NAND2X1_343 ( .gnd(gnd), .vdd(vdd), .A(_2349_), .B(_2347_), .Y(_2622_) );
OAI21X1 OAI21X1_702 ( .gnd(gnd), .vdd(vdd), .A(_2348_), .B(_2322__bF_buf4), .C(_2622_), .Y(_2623_) );
INVX1 INVX1_186 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_43_), .Y(_2624_) );
OAI21X1 OAI21X1_703 ( .gnd(gnd), .vdd(vdd), .A(_2569__bF_buf3), .B(_2570__bF_buf3), .C(_2624_), .Y(_2625_) );
NOR2X1 NOR2X1_542 ( .gnd(gnd), .vdd(vdd), .A(_2624_), .B(_2574__bF_buf4), .Y(_2626_) );
INVX1 INVX1_187 ( .gnd(gnd), .vdd(vdd), .A(_2626_), .Y(_2627_) );
NAND2X1 NAND2X1_344 ( .gnd(gnd), .vdd(vdd), .A(_2625_), .B(_2627_), .Y(_2628_) );
XOR2X1 XOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_2623_), .B(_2628_), .Y(_2629_) );
OAI21X1 OAI21X1_704 ( .gnd(gnd), .vdd(vdd), .A(_2629_), .B(_925__bF_buf4), .C(_926__bF_buf3), .Y(_2630_) );
AOI21X1 AOI21X1_426 ( .gnd(gnd), .vdd(vdd), .A(_2621_), .B(_2611_), .C(_2630_), .Y(_2631_) );
NOR2X1 NOR2X1_543 ( .gnd(gnd), .vdd(vdd), .A(_2131_), .B(_2133_), .Y(_2632_) );
OAI21X1 OAI21X1_705 ( .gnd(gnd), .vdd(vdd), .A(_2632_), .B(_2358_), .C(_2357_), .Y(_2633_) );
INVX1 INVX1_188 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_51_), .Y(_2634_) );
OAI21X1 OAI21X1_706 ( .gnd(gnd), .vdd(vdd), .A(_2569__bF_buf2), .B(_2570__bF_buf2), .C(_2634_), .Y(_2635_) );
NOR2X1 NOR2X1_544 ( .gnd(gnd), .vdd(vdd), .A(_2634_), .B(_2574__bF_buf3), .Y(_2636_) );
INVX1 INVX1_189 ( .gnd(gnd), .vdd(vdd), .A(_2636_), .Y(_2637_) );
NAND2X1 NAND2X1_345 ( .gnd(gnd), .vdd(vdd), .A(_2635_), .B(_2637_), .Y(_2638_) );
XNOR2X1 XNOR2X1_62 ( .gnd(gnd), .vdd(vdd), .A(_2633_), .B(_2638_), .Y(_2639_) );
OAI21X1 OAI21X1_707 ( .gnd(gnd), .vdd(vdd), .A(_2639_), .B(_926__bF_buf2), .C(_924__bF_buf2), .Y(_2640_) );
OAI21X1 OAI21X1_708 ( .gnd(gnd), .vdd(vdd), .A(_813_), .B(_2322__bF_buf3), .C(_2366_), .Y(_2641_) );
OAI21X1 OAI21X1_709 ( .gnd(gnd), .vdd(vdd), .A(_2569__bF_buf1), .B(_2570__bF_buf1), .C(_816_), .Y(_2642_) );
INVX1 INVX1_190 ( .gnd(gnd), .vdd(vdd), .A(_2642_), .Y(_2643_) );
NOR2X1 NOR2X1_545 ( .gnd(gnd), .vdd(vdd), .A(_816_), .B(_2574__bF_buf2), .Y(_2644_) );
NOR2X1 NOR2X1_546 ( .gnd(gnd), .vdd(vdd), .A(_2643_), .B(_2644_), .Y(_2645_) );
XOR2X1 XOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(_2641_), .B(_2645_), .Y(_2646_) );
AOI21X1 AOI21X1_427 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe22_bF_buf1), .B(_2646_), .C(micro_hash_ucr_pipe24_bF_buf3), .Y(_2647_) );
OAI21X1 OAI21X1_710 ( .gnd(gnd), .vdd(vdd), .A(_2631_), .B(_2640_), .C(_2647_), .Y(_2648_) );
OAI21X1 OAI21X1_711 ( .gnd(gnd), .vdd(vdd), .A(_859_), .B(_2322__bF_buf2), .C(_2373_), .Y(_2649_) );
OAI21X1 OAI21X1_712 ( .gnd(gnd), .vdd(vdd), .A(_2569__bF_buf0), .B(_2570__bF_buf0), .C(_862_), .Y(_2650_) );
NOR2X1 NOR2X1_547 ( .gnd(gnd), .vdd(vdd), .A(_862_), .B(_2574__bF_buf1), .Y(_2651_) );
INVX1 INVX1_191 ( .gnd(gnd), .vdd(vdd), .A(_2651_), .Y(_2652_) );
NAND2X1 NAND2X1_346 ( .gnd(gnd), .vdd(vdd), .A(_2650_), .B(_2652_), .Y(_2653_) );
AOI21X1 AOI21X1_428 ( .gnd(gnd), .vdd(vdd), .A(_2653_), .B(_2649_), .C(_919__bF_buf0), .Y(_2654_) );
OAI21X1 OAI21X1_713 ( .gnd(gnd), .vdd(vdd), .A(_2649_), .B(_2653_), .C(_2654_), .Y(_2655_) );
AND2X2 AND2X2_212 ( .gnd(gnd), .vdd(vdd), .A(_2655_), .B(_920__bF_buf2), .Y(_2656_) );
OAI21X1 OAI21X1_714 ( .gnd(gnd), .vdd(vdd), .A(_835_), .B(_2322__bF_buf1), .C(_2382_), .Y(_2657_) );
OAI21X1 OAI21X1_715 ( .gnd(gnd), .vdd(vdd), .A(_2569__bF_buf4), .B(_2570__bF_buf4), .C(_838_), .Y(_2658_) );
NOR2X1 NOR2X1_548 ( .gnd(gnd), .vdd(vdd), .A(_838_), .B(_2574__bF_buf0), .Y(_2659_) );
INVX1 INVX1_192 ( .gnd(gnd), .vdd(vdd), .A(_2659_), .Y(_2660_) );
NAND2X1 NAND2X1_347 ( .gnd(gnd), .vdd(vdd), .A(_2658_), .B(_2660_), .Y(_2661_) );
XOR2X1 XOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_2657_), .B(_2661_), .Y(_2662_) );
OAI21X1 OAI21X1_716 ( .gnd(gnd), .vdd(vdd), .A(_2662_), .B(_920__bF_buf1), .C(_918__bF_buf0), .Y(_2663_) );
AOI21X1 AOI21X1_429 ( .gnd(gnd), .vdd(vdd), .A(_2656_), .B(_2648_), .C(_2663_), .Y(_2664_) );
NAND3X1 NAND3X1_104 ( .gnd(gnd), .vdd(vdd), .A(_2386_), .B(_2388_), .C(_2385_), .Y(_2665_) );
OAI21X1 OAI21X1_717 ( .gnd(gnd), .vdd(vdd), .A(_746_), .B(_2322__bF_buf0), .C(_2665_), .Y(_2666_) );
OAI21X1 OAI21X1_718 ( .gnd(gnd), .vdd(vdd), .A(_2569__bF_buf3), .B(_2570__bF_buf3), .C(_749_), .Y(_2667_) );
NOR2X1 NOR2X1_549 ( .gnd(gnd), .vdd(vdd), .A(_749_), .B(_2574__bF_buf4), .Y(_2668_) );
INVX1 INVX1_193 ( .gnd(gnd), .vdd(vdd), .A(_2668_), .Y(_2669_) );
NAND2X1 NAND2X1_348 ( .gnd(gnd), .vdd(vdd), .A(_2667_), .B(_2669_), .Y(_2670_) );
XNOR2X1 XNOR2X1_63 ( .gnd(gnd), .vdd(vdd), .A(_2666_), .B(_2670_), .Y(_2671_) );
OAI21X1 OAI21X1_719 ( .gnd(gnd), .vdd(vdd), .A(_2671_), .B(_918__bF_buf4), .C(_913__bF_buf3), .Y(_2672_) );
OAI21X1 OAI21X1_720 ( .gnd(gnd), .vdd(vdd), .A(_786_), .B(_2322__bF_buf5), .C(_2397_), .Y(_2673_) );
OAI21X1 OAI21X1_721 ( .gnd(gnd), .vdd(vdd), .A(_2569__bF_buf2), .B(_2570__bF_buf2), .C(_790_), .Y(_2674_) );
INVX1 INVX1_194 ( .gnd(gnd), .vdd(vdd), .A(_2674_), .Y(_2675_) );
NOR2X1 NOR2X1_550 ( .gnd(gnd), .vdd(vdd), .A(_790_), .B(_2574__bF_buf3), .Y(_2676_) );
NOR2X1 NOR2X1_551 ( .gnd(gnd), .vdd(vdd), .A(_2675_), .B(_2676_), .Y(_2677_) );
XOR2X1 XOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(_2673_), .B(_2677_), .Y(_2678_) );
AOI21X1 AOI21X1_430 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe30_bF_buf2), .B(_2678_), .C(micro_hash_ucr_pipe32_bF_buf3), .Y(_2679_) );
OAI21X1 OAI21X1_722 ( .gnd(gnd), .vdd(vdd), .A(_2664_), .B(_2672_), .C(_2679_), .Y(_2680_) );
NAND3X1 NAND3X1_105 ( .gnd(gnd), .vdd(vdd), .A(_2404_), .B(_2406_), .C(_2403_), .Y(_2681_) );
OAI21X1 OAI21X1_723 ( .gnd(gnd), .vdd(vdd), .A(_648_), .B(_2322__bF_buf4), .C(_2681_), .Y(_2682_) );
OAI21X1 OAI21X1_724 ( .gnd(gnd), .vdd(vdd), .A(_2569__bF_buf1), .B(_2570__bF_buf1), .C(_652_), .Y(_2683_) );
NOR2X1 NOR2X1_552 ( .gnd(gnd), .vdd(vdd), .A(_652_), .B(_2574__bF_buf2), .Y(_2684_) );
INVX1 INVX1_195 ( .gnd(gnd), .vdd(vdd), .A(_2684_), .Y(_2685_) );
NAND2X1 NAND2X1_349 ( .gnd(gnd), .vdd(vdd), .A(_2683_), .B(_2685_), .Y(_2686_) );
AOI21X1 AOI21X1_431 ( .gnd(gnd), .vdd(vdd), .A(_2686_), .B(_2682_), .C(_914__bF_buf4), .Y(_2687_) );
OAI21X1 OAI21X1_725 ( .gnd(gnd), .vdd(vdd), .A(_2682_), .B(_2686_), .C(_2687_), .Y(_2688_) );
AND2X2 AND2X2_213 ( .gnd(gnd), .vdd(vdd), .A(_2688_), .B(_912__bF_buf0), .Y(_2689_) );
OAI21X1 OAI21X1_726 ( .gnd(gnd), .vdd(vdd), .A(_676_), .B(_2322__bF_buf3), .C(_2417_), .Y(_2690_) );
OAI21X1 OAI21X1_727 ( .gnd(gnd), .vdd(vdd), .A(_2569__bF_buf0), .B(_2570__bF_buf0), .C(_680_), .Y(_2691_) );
NOR2X1 NOR2X1_553 ( .gnd(gnd), .vdd(vdd), .A(_680_), .B(_2574__bF_buf1), .Y(_2692_) );
INVX1 INVX1_196 ( .gnd(gnd), .vdd(vdd), .A(_2692_), .Y(_2693_) );
NAND2X1 NAND2X1_350 ( .gnd(gnd), .vdd(vdd), .A(_2691_), .B(_2693_), .Y(_2694_) );
XOR2X1 XOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_2690_), .B(_2694_), .Y(_2695_) );
OAI21X1 OAI21X1_728 ( .gnd(gnd), .vdd(vdd), .A(_2695_), .B(_912__bF_buf4), .C(_907__bF_buf4), .Y(_2696_) );
AOI21X1 AOI21X1_432 ( .gnd(gnd), .vdd(vdd), .A(_2689_), .B(_2680_), .C(_2696_), .Y(_2697_) );
NAND3X1 NAND3X1_106 ( .gnd(gnd), .vdd(vdd), .A(_2421_), .B(_2423_), .C(_2420_), .Y(_2698_) );
OAI21X1 OAI21X1_729 ( .gnd(gnd), .vdd(vdd), .A(_510_), .B(_2322__bF_buf2), .C(_2698_), .Y(_2699_) );
OAI21X1 OAI21X1_730 ( .gnd(gnd), .vdd(vdd), .A(_2569__bF_buf4), .B(_2570__bF_buf4), .C(_514_), .Y(_2700_) );
NOR2X1 NOR2X1_554 ( .gnd(gnd), .vdd(vdd), .A(_514_), .B(_2574__bF_buf0), .Y(_2701_) );
INVX1 INVX1_197 ( .gnd(gnd), .vdd(vdd), .A(_2701_), .Y(_2702_) );
NAND2X1 NAND2X1_351 ( .gnd(gnd), .vdd(vdd), .A(_2700_), .B(_2702_), .Y(_2703_) );
XNOR2X1 XNOR2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_2699_), .B(_2703_), .Y(_2704_) );
OAI21X1 OAI21X1_731 ( .gnd(gnd), .vdd(vdd), .A(_2704_), .B(_907__bF_buf3), .C(_908__bF_buf1), .Y(_2705_) );
OAI21X1 OAI21X1_732 ( .gnd(gnd), .vdd(vdd), .A(_566_), .B(_2322__bF_buf1), .C(_2435_), .Y(_2706_) );
OAI21X1 OAI21X1_733 ( .gnd(gnd), .vdd(vdd), .A(_2569__bF_buf3), .B(_2570__bF_buf3), .C(_570_), .Y(_2707_) );
NOR2X1 NOR2X1_555 ( .gnd(gnd), .vdd(vdd), .A(_570_), .B(_2574__bF_buf4), .Y(_2708_) );
INVX1 INVX1_198 ( .gnd(gnd), .vdd(vdd), .A(_2708_), .Y(_2709_) );
NAND2X1 NAND2X1_352 ( .gnd(gnd), .vdd(vdd), .A(_2707_), .B(_2709_), .Y(_2710_) );
XNOR2X1 XNOR2X1_65 ( .gnd(gnd), .vdd(vdd), .A(_2706_), .B(_2710_), .Y(_2711_) );
AOI21X1 AOI21X1_433 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe38_bF_buf0), .B(_2711_), .C(micro_hash_ucr_pipe40_bF_buf0), .Y(_2712_) );
OAI21X1 OAI21X1_734 ( .gnd(gnd), .vdd(vdd), .A(_2697_), .B(_2705_), .C(_2712_), .Y(_2713_) );
NAND3X1 NAND3X1_107 ( .gnd(gnd), .vdd(vdd), .A(_2442_), .B(_2444_), .C(_2441_), .Y(_2714_) );
OAI21X1 OAI21X1_735 ( .gnd(gnd), .vdd(vdd), .A(_538_), .B(_2322__bF_buf0), .C(_2714_), .Y(_2715_) );
OAI21X1 OAI21X1_736 ( .gnd(gnd), .vdd(vdd), .A(_2569__bF_buf2), .B(_2570__bF_buf2), .C(_542_), .Y(_2716_) );
NOR2X1 NOR2X1_556 ( .gnd(gnd), .vdd(vdd), .A(_542_), .B(_2574__bF_buf3), .Y(_2717_) );
INVX1 INVX1_199 ( .gnd(gnd), .vdd(vdd), .A(_2717_), .Y(_2718_) );
NAND2X1 NAND2X1_353 ( .gnd(gnd), .vdd(vdd), .A(_2716_), .B(_2718_), .Y(_2719_) );
AOI21X1 AOI21X1_434 ( .gnd(gnd), .vdd(vdd), .A(_2719_), .B(_2715_), .C(_906__bF_buf0), .Y(_2720_) );
OAI21X1 OAI21X1_737 ( .gnd(gnd), .vdd(vdd), .A(_2715_), .B(_2719_), .C(_2720_), .Y(_2721_) );
AND2X2 AND2X2_214 ( .gnd(gnd), .vdd(vdd), .A(_2721_), .B(_901__bF_buf2), .Y(_2722_) );
OAI21X1 OAI21X1_738 ( .gnd(gnd), .vdd(vdd), .A(_787_), .B(_2322__bF_buf5), .C(_2449_), .Y(_2723_) );
OAI21X1 OAI21X1_739 ( .gnd(gnd), .vdd(vdd), .A(_2569__bF_buf1), .B(_2570__bF_buf1), .C(_791_), .Y(_2724_) );
NOR2X1 NOR2X1_557 ( .gnd(gnd), .vdd(vdd), .A(_791_), .B(_2574__bF_buf2), .Y(_2725_) );
INVX1 INVX1_200 ( .gnd(gnd), .vdd(vdd), .A(_2725_), .Y(_2726_) );
NAND2X1 NAND2X1_354 ( .gnd(gnd), .vdd(vdd), .A(_2724_), .B(_2726_), .Y(_2727_) );
XOR2X1 XOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_2723_), .B(_2727_), .Y(_2728_) );
OAI21X1 OAI21X1_740 ( .gnd(gnd), .vdd(vdd), .A(_2728_), .B(_901__bF_buf1), .C(_902__bF_buf4), .Y(_2729_) );
AOI21X1 AOI21X1_435 ( .gnd(gnd), .vdd(vdd), .A(_2722_), .B(_2713_), .C(_2729_), .Y(_2730_) );
OAI21X1 OAI21X1_741 ( .gnd(gnd), .vdd(vdd), .A(_619_), .B(_2322__bF_buf4), .C(_2457_), .Y(_2731_) );
OAI21X1 OAI21X1_742 ( .gnd(gnd), .vdd(vdd), .A(_2569__bF_buf0), .B(_2570__bF_buf0), .C(_623_), .Y(_2732_) );
NOR2X1 NOR2X1_558 ( .gnd(gnd), .vdd(vdd), .A(_623_), .B(_2574__bF_buf1), .Y(_2733_) );
INVX1 INVX1_201 ( .gnd(gnd), .vdd(vdd), .A(_2733_), .Y(_2734_) );
NAND2X1 NAND2X1_355 ( .gnd(gnd), .vdd(vdd), .A(_2732_), .B(_2734_), .Y(_2735_) );
XNOR2X1 XNOR2X1_66 ( .gnd(gnd), .vdd(vdd), .A(_2731_), .B(_2735_), .Y(_2736_) );
OAI21X1 OAI21X1_743 ( .gnd(gnd), .vdd(vdd), .A(_2736_), .B(_902__bF_buf3), .C(_900__bF_buf3), .Y(_2737_) );
NAND3X1 NAND3X1_108 ( .gnd(gnd), .vdd(vdd), .A(_2462_), .B(_2464_), .C(_2461_), .Y(_2738_) );
OAI21X1 OAI21X1_744 ( .gnd(gnd), .vdd(vdd), .A(_677_), .B(_2322__bF_buf3), .C(_2738_), .Y(_2739_) );
OAI21X1 OAI21X1_745 ( .gnd(gnd), .vdd(vdd), .A(_2569__bF_buf4), .B(_2570__bF_buf4), .C(_681_), .Y(_2740_) );
INVX1 INVX1_202 ( .gnd(gnd), .vdd(vdd), .A(_2740_), .Y(_2741_) );
NOR2X1 NOR2X1_559 ( .gnd(gnd), .vdd(vdd), .A(_681_), .B(_2574__bF_buf0), .Y(_2742_) );
NOR2X1 NOR2X1_560 ( .gnd(gnd), .vdd(vdd), .A(_2741_), .B(_2742_), .Y(_2743_) );
XOR2X1 XOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_2739_), .B(_2743_), .Y(_2744_) );
AOI21X1 AOI21X1_436 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe46_bF_buf2), .B(_2744_), .C(micro_hash_ucr_pipe48_bF_buf0), .Y(_2745_) );
OAI21X1 OAI21X1_746 ( .gnd(gnd), .vdd(vdd), .A(_2730_), .B(_2737_), .C(_2745_), .Y(_2746_) );
OAI21X1 OAI21X1_747 ( .gnd(gnd), .vdd(vdd), .A(_725_), .B(_2322__bF_buf2), .C(_2470_), .Y(_2747_) );
OAI21X1 OAI21X1_748 ( .gnd(gnd), .vdd(vdd), .A(_2569__bF_buf3), .B(_2570__bF_buf3), .C(_728_), .Y(_2748_) );
NOR2X1 NOR2X1_561 ( .gnd(gnd), .vdd(vdd), .A(_728_), .B(_2574__bF_buf4), .Y(_2749_) );
INVX1 INVX1_203 ( .gnd(gnd), .vdd(vdd), .A(_2749_), .Y(_2750_) );
NAND2X1 NAND2X1_356 ( .gnd(gnd), .vdd(vdd), .A(_2748_), .B(_2750_), .Y(_2751_) );
AOI21X1 AOI21X1_437 ( .gnd(gnd), .vdd(vdd), .A(_2751_), .B(_2747_), .C(_895__bF_buf1), .Y(_2752_) );
OAI21X1 OAI21X1_749 ( .gnd(gnd), .vdd(vdd), .A(_2747_), .B(_2751_), .C(_2752_), .Y(_2753_) );
AND2X2 AND2X2_215 ( .gnd(gnd), .vdd(vdd), .A(_2753_), .B(_896__bF_buf0), .Y(_2754_) );
OAI21X1 OAI21X1_750 ( .gnd(gnd), .vdd(vdd), .A(_702_), .B(_2322__bF_buf1), .C(_2476_), .Y(_2755_) );
OAI21X1 OAI21X1_751 ( .gnd(gnd), .vdd(vdd), .A(_2569__bF_buf2), .B(_2570__bF_buf2), .C(_705_), .Y(_2756_) );
NOR2X1 NOR2X1_562 ( .gnd(gnd), .vdd(vdd), .A(_705_), .B(_2574__bF_buf3), .Y(_2757_) );
INVX1 INVX1_204 ( .gnd(gnd), .vdd(vdd), .A(_2757_), .Y(_2758_) );
NAND2X1 NAND2X1_357 ( .gnd(gnd), .vdd(vdd), .A(_2756_), .B(_2758_), .Y(_2759_) );
XOR2X1 XOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(_2755_), .B(_2759_), .Y(_2760_) );
OAI21X1 OAI21X1_752 ( .gnd(gnd), .vdd(vdd), .A(_2760_), .B(_896__bF_buf4), .C(_894__bF_buf1), .Y(_2761_) );
AOI21X1 AOI21X1_438 ( .gnd(gnd), .vdd(vdd), .A(_2754_), .B(_2746_), .C(_2761_), .Y(_2762_) );
OAI21X1 OAI21X1_753 ( .gnd(gnd), .vdd(vdd), .A(_593_), .B(_2322__bF_buf0), .C(_2483_), .Y(_2763_) );
OAI21X1 OAI21X1_754 ( .gnd(gnd), .vdd(vdd), .A(_2569__bF_buf1), .B(_2570__bF_buf1), .C(_596_), .Y(_2764_) );
NOR2X1 NOR2X1_563 ( .gnd(gnd), .vdd(vdd), .A(_596_), .B(_2574__bF_buf2), .Y(_2765_) );
INVX1 INVX1_205 ( .gnd(gnd), .vdd(vdd), .A(_2765_), .Y(_2766_) );
NAND2X1 NAND2X1_358 ( .gnd(gnd), .vdd(vdd), .A(_2764_), .B(_2766_), .Y(_2767_) );
XNOR2X1 XNOR2X1_67 ( .gnd(gnd), .vdd(vdd), .A(_2763_), .B(_2767_), .Y(_2768_) );
OAI21X1 OAI21X1_755 ( .gnd(gnd), .vdd(vdd), .A(_2768_), .B(_894__bF_buf0), .C(_889__bF_buf0), .Y(_2769_) );
NAND3X1 NAND3X1_109 ( .gnd(gnd), .vdd(vdd), .A(_2491_), .B(_2493_), .C(_2490_), .Y(_2770_) );
OAI21X1 OAI21X1_756 ( .gnd(gnd), .vdd(vdd), .A(_649_), .B(_2322__bF_buf5), .C(_2770_), .Y(_2771_) );
OAI21X1 OAI21X1_757 ( .gnd(gnd), .vdd(vdd), .A(_2569__bF_buf0), .B(_2570__bF_buf0), .C(_653_), .Y(_2772_) );
INVX1 INVX1_206 ( .gnd(gnd), .vdd(vdd), .A(_2772_), .Y(_2773_) );
NOR2X1 NOR2X1_564 ( .gnd(gnd), .vdd(vdd), .A(_653_), .B(_2574__bF_buf1), .Y(_2774_) );
NOR2X1 NOR2X1_565 ( .gnd(gnd), .vdd(vdd), .A(_2773_), .B(_2774_), .Y(_2775_) );
XOR2X1 XOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_2771_), .B(_2775_), .Y(_2776_) );
AOI21X1 AOI21X1_439 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe54_bF_buf0), .B(_2776_), .C(micro_hash_ucr_pipe56_bF_buf3), .Y(_2777_) );
OAI21X1 OAI21X1_758 ( .gnd(gnd), .vdd(vdd), .A(_2762_), .B(_2769_), .C(_2777_), .Y(_2778_) );
OAI21X1 OAI21X1_759 ( .gnd(gnd), .vdd(vdd), .A(_620_), .B(_2322__bF_buf4), .C(_2498_), .Y(_2779_) );
OAI21X1 OAI21X1_760 ( .gnd(gnd), .vdd(vdd), .A(_2569__bF_buf4), .B(_2570__bF_buf4), .C(_624_), .Y(_2780_) );
NOR2X1 NOR2X1_566 ( .gnd(gnd), .vdd(vdd), .A(_624_), .B(_2574__bF_buf0), .Y(_2781_) );
INVX1 INVX1_207 ( .gnd(gnd), .vdd(vdd), .A(_2781_), .Y(_2782_) );
NAND2X1 NAND2X1_359 ( .gnd(gnd), .vdd(vdd), .A(_2780_), .B(_2782_), .Y(_2783_) );
AOI21X1 AOI21X1_440 ( .gnd(gnd), .vdd(vdd), .A(_2783_), .B(_2779_), .C(_890__bF_buf2), .Y(_2784_) );
OAI21X1 OAI21X1_761 ( .gnd(gnd), .vdd(vdd), .A(_2779_), .B(_2783_), .C(_2784_), .Y(_2785_) );
AND2X2 AND2X2_216 ( .gnd(gnd), .vdd(vdd), .A(_2785_), .B(_888__bF_buf0), .Y(_2786_) );
OAI21X1 OAI21X1_762 ( .gnd(gnd), .vdd(vdd), .A(_511_), .B(_2322__bF_buf3), .C(_2506_), .Y(_2787_) );
OAI21X1 OAI21X1_763 ( .gnd(gnd), .vdd(vdd), .A(_2569__bF_buf3), .B(_2570__bF_buf3), .C(_515_), .Y(_2788_) );
NOR2X1 NOR2X1_567 ( .gnd(gnd), .vdd(vdd), .A(_515_), .B(_2574__bF_buf4), .Y(_2789_) );
INVX1 INVX1_208 ( .gnd(gnd), .vdd(vdd), .A(_2789_), .Y(_2790_) );
NAND2X1 NAND2X1_360 ( .gnd(gnd), .vdd(vdd), .A(_2788_), .B(_2790_), .Y(_2791_) );
XOR2X1 XOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(_2787_), .B(_2791_), .Y(_2792_) );
OAI21X1 OAI21X1_764 ( .gnd(gnd), .vdd(vdd), .A(_2792_), .B(_888__bF_buf3), .C(_883__bF_buf2), .Y(_2793_) );
AOI21X1 AOI21X1_441 ( .gnd(gnd), .vdd(vdd), .A(_2786_), .B(_2778_), .C(_2793_), .Y(_2794_) );
NAND3X1 NAND3X1_110 ( .gnd(gnd), .vdd(vdd), .A(_2511_), .B(_2513_), .C(_2510_), .Y(_2795_) );
OAI21X1 OAI21X1_765 ( .gnd(gnd), .vdd(vdd), .A(_567_), .B(_2322__bF_buf2), .C(_2795_), .Y(_2796_) );
OAI21X1 OAI21X1_766 ( .gnd(gnd), .vdd(vdd), .A(_2569__bF_buf2), .B(_2570__bF_buf2), .C(_571_), .Y(_2797_) );
NOR2X1 NOR2X1_568 ( .gnd(gnd), .vdd(vdd), .A(_571_), .B(_2574__bF_buf3), .Y(_2798_) );
INVX1 INVX1_209 ( .gnd(gnd), .vdd(vdd), .A(_2798_), .Y(_2799_) );
NAND2X1 NAND2X1_361 ( .gnd(gnd), .vdd(vdd), .A(_2797_), .B(_2799_), .Y(_2800_) );
XNOR2X1 XNOR2X1_68 ( .gnd(gnd), .vdd(vdd), .A(_2800_), .B(_2796_), .Y(_2801_) );
OAI21X1 OAI21X1_767 ( .gnd(gnd), .vdd(vdd), .A(_2801_), .B(_883__bF_buf1), .C(_884__bF_buf4), .Y(_2802_) );
OAI21X1 OAI21X1_768 ( .gnd(gnd), .vdd(vdd), .A(_539_), .B(_2322__bF_buf1), .C(_2518_), .Y(_2803_) );
OAI21X1 OAI21X1_769 ( .gnd(gnd), .vdd(vdd), .A(_2569__bF_buf1), .B(_2570__bF_buf1), .C(_543_), .Y(_2804_) );
INVX1 INVX1_210 ( .gnd(gnd), .vdd(vdd), .A(_2804_), .Y(_2805_) );
NOR2X1 NOR2X1_569 ( .gnd(gnd), .vdd(vdd), .A(_543_), .B(_2574__bF_buf2), .Y(_2806_) );
NOR2X1 NOR2X1_570 ( .gnd(gnd), .vdd(vdd), .A(_2805_), .B(_2806_), .Y(_2807_) );
XOR2X1 XOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_2803_), .B(_2807_), .Y(_2808_) );
AOI21X1 AOI21X1_442 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe62_bF_buf0), .B(_2808_), .C(micro_hash_ucr_pipe64_bF_buf3), .Y(_2809_) );
OAI21X1 OAI21X1_770 ( .gnd(gnd), .vdd(vdd), .A(_2794_), .B(_2802_), .C(_2809_), .Y(_2810_) );
NAND3X1 NAND3X1_111 ( .gnd(gnd), .vdd(vdd), .A(_2528_), .B(_2530_), .C(_2526_), .Y(_2811_) );
OAI21X1 OAI21X1_771 ( .gnd(gnd), .vdd(vdd), .A(_2527_), .B(_2322__bF_buf0), .C(_2811_), .Y(_2812_) );
INVX1 INVX1_211 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_227_), .Y(_2813_) );
OAI21X1 OAI21X1_772 ( .gnd(gnd), .vdd(vdd), .A(_2569__bF_buf0), .B(_2570__bF_buf0), .C(_2813_), .Y(_2814_) );
NOR2X1 NOR2X1_571 ( .gnd(gnd), .vdd(vdd), .A(_2813_), .B(_2574__bF_buf1), .Y(_2815_) );
INVX1 INVX1_212 ( .gnd(gnd), .vdd(vdd), .A(_2815_), .Y(_2816_) );
NAND2X1 NAND2X1_362 ( .gnd(gnd), .vdd(vdd), .A(_2814_), .B(_2816_), .Y(_2817_) );
AOI21X1 AOI21X1_443 ( .gnd(gnd), .vdd(vdd), .A(_2817_), .B(_2812_), .C(_882__bF_buf3), .Y(_2818_) );
OAI21X1 OAI21X1_773 ( .gnd(gnd), .vdd(vdd), .A(_2812_), .B(_2817_), .C(_2818_), .Y(_2819_) );
AND2X2 AND2X2_217 ( .gnd(gnd), .vdd(vdd), .A(_2819_), .B(_877__bF_buf0), .Y(_2820_) );
OAI21X1 OAI21X1_774 ( .gnd(gnd), .vdd(vdd), .A(_2535_), .B(_2322__bF_buf5), .C(_2538_), .Y(_2821_) );
INVX1 INVX1_213 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_235_), .Y(_2822_) );
OAI21X1 OAI21X1_775 ( .gnd(gnd), .vdd(vdd), .A(_2569__bF_buf4), .B(_2570__bF_buf4), .C(_2822_), .Y(_2823_) );
NOR2X1 NOR2X1_572 ( .gnd(gnd), .vdd(vdd), .A(_2822_), .B(_2574__bF_buf0), .Y(_2824_) );
INVX1 INVX1_214 ( .gnd(gnd), .vdd(vdd), .A(_2824_), .Y(_2825_) );
NAND2X1 NAND2X1_363 ( .gnd(gnd), .vdd(vdd), .A(_2823_), .B(_2825_), .Y(_2826_) );
XOR2X1 XOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(_2826_), .B(_2821_), .Y(_2827_) );
OAI21X1 OAI21X1_776 ( .gnd(gnd), .vdd(vdd), .A(_2827_), .B(_877__bF_buf3), .C(_878__bF_buf1), .Y(_2828_) );
AOI21X1 AOI21X1_444 ( .gnd(gnd), .vdd(vdd), .A(_2820_), .B(_2810_), .C(_2828_), .Y(_2829_) );
NAND3X1 NAND3X1_112 ( .gnd(gnd), .vdd(vdd), .A(_2546_), .B(_2548_), .C(_2544_), .Y(_2830_) );
OAI21X1 OAI21X1_777 ( .gnd(gnd), .vdd(vdd), .A(_2545_), .B(_2322__bF_buf4), .C(_2830_), .Y(_2831_) );
INVX1 INVX1_215 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_243_), .Y(_2832_) );
OAI21X1 OAI21X1_778 ( .gnd(gnd), .vdd(vdd), .A(_2569__bF_buf3), .B(_2570__bF_buf3), .C(_2832_), .Y(_2833_) );
INVX1 INVX1_216 ( .gnd(gnd), .vdd(vdd), .A(_2833_), .Y(_2834_) );
NOR2X1 NOR2X1_573 ( .gnd(gnd), .vdd(vdd), .A(_2832_), .B(_2574__bF_buf4), .Y(_2835_) );
NOR2X1 NOR2X1_574 ( .gnd(gnd), .vdd(vdd), .A(_2834_), .B(_2835_), .Y(_2836_) );
XOR2X1 XOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(_2831_), .B(_2836_), .Y(_2837_) );
OAI21X1 OAI21X1_779 ( .gnd(gnd), .vdd(vdd), .A(_2837_), .B(_878__bF_buf0), .C(_1949_), .Y(_2838_) );
NOR2X1 NOR2X1_575 ( .gnd(gnd), .vdd(vdd), .A(_2557_), .B(_2559_), .Y(_2839_) );
INVX2 INVX2_112 ( .gnd(gnd), .vdd(vdd), .A(_2839_), .Y(_2840_) );
INVX1 INVX1_217 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_251_), .Y(_2841_) );
OAI21X1 OAI21X1_780 ( .gnd(gnd), .vdd(vdd), .A(_2569__bF_buf2), .B(_2570__bF_buf2), .C(_2841_), .Y(_2842_) );
INVX1 INVX1_218 ( .gnd(gnd), .vdd(vdd), .A(_2842_), .Y(_2843_) );
NOR2X1 NOR2X1_576 ( .gnd(gnd), .vdd(vdd), .A(_2841_), .B(_2574__bF_buf3), .Y(_2844_) );
NOR2X1 NOR2X1_577 ( .gnd(gnd), .vdd(vdd), .A(_2843_), .B(_2844_), .Y(_2845_) );
AND2X2 AND2X2_218 ( .gnd(gnd), .vdd(vdd), .A(_2840_), .B(_2845_), .Y(_2846_) );
OAI21X1 OAI21X1_781 ( .gnd(gnd), .vdd(vdd), .A(_2840_), .B(_2845_), .C(_369_), .Y(_2847_) );
OAI22X1 OAI22X1_52 ( .gnd(gnd), .vdd(vdd), .A(_2846_), .B(_2847_), .C(_2829_), .D(_2838_), .Y(_299__3_) );
AOI21X1 AOI21X1_445 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_k_3_), .B(micro_hash_ucr_x_3_), .C(_2569__bF_buf1), .Y(_2848_) );
NOR2X1 NOR2X1_578 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_k_4_), .B(micro_hash_ucr_x_4_), .Y(_2849_) );
INVX1 INVX1_219 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_k_4_), .Y(_2850_) );
INVX1 INVX1_220 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_x_4_), .Y(_2851_) );
NOR2X1 NOR2X1_579 ( .gnd(gnd), .vdd(vdd), .A(_2850_), .B(_2851_), .Y(_2852_) );
NOR2X1 NOR2X1_580 ( .gnd(gnd), .vdd(vdd), .A(_2849_), .B(_2852_), .Y(_2853_) );
INVX1 INVX1_221 ( .gnd(gnd), .vdd(vdd), .A(_2853_), .Y(_2854_) );
OR2X2 OR2X2_32 ( .gnd(gnd), .vdd(vdd), .A(_2848_), .B(_2854_), .Y(_2855_) );
OAI21X1 OAI21X1_782 ( .gnd(gnd), .vdd(vdd), .A(_2849_), .B(_2852_), .C(_2848_), .Y(_2856_) );
NAND2X1 NAND2X1_364 ( .gnd(gnd), .vdd(vdd), .A(_2856_), .B(_2855_), .Y(_2857_) );
XOR2X1 XOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(_2857__bF_buf5), .B(micro_hash_ucr_Wx_4_), .Y(_2858_) );
AOI21X1 AOI21X1_446 ( .gnd(gnd), .vdd(vdd), .A(_2571_), .B(_2562_), .C(_2575_), .Y(_2859_) );
AND2X2 AND2X2_219 ( .gnd(gnd), .vdd(vdd), .A(_2859_), .B(_2858_), .Y(_2860_) );
NOR2X1 NOR2X1_581 ( .gnd(gnd), .vdd(vdd), .A(_2858_), .B(_2859_), .Y(_2861_) );
OAI21X1 OAI21X1_783 ( .gnd(gnd), .vdd(vdd), .A(_2860_), .B(_2861_), .C(micro_hash_ucr_pipe8), .Y(_2862_) );
XOR2X1 XOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_2857__bF_buf4), .B(micro_hash_ucr_Wx_12_), .Y(_2863_) );
AOI21X1 AOI21X1_447 ( .gnd(gnd), .vdd(vdd), .A(_2586_), .B(_2584_), .C(_2588_), .Y(_2864_) );
XOR2X1 XOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(_2864_), .B(_2863_), .Y(_2865_) );
NAND2X1 NAND2X1_365 ( .gnd(gnd), .vdd(vdd), .A(_1394_), .B(_937_), .Y(_2866_) );
OAI21X1 OAI21X1_784 ( .gnd(gnd), .vdd(vdd), .A(H_20_), .B(_937_), .C(_2866_), .Y(_2867_) );
AOI21X1 AOI21X1_448 ( .gnd(gnd), .vdd(vdd), .A(_938_), .B(_2867_), .C(micro_hash_ucr_pipe10), .Y(_2868_) );
AOI22X1 AOI22X1_29 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe10), .B(_2865_), .C(_2862_), .D(_2868_), .Y(_2869_) );
XNOR2X1 XNOR2X1_69 ( .gnd(gnd), .vdd(vdd), .A(_2857__bF_buf3), .B(micro_hash_ucr_Wx_20_), .Y(_2870_) );
INVX1 INVX1_222 ( .gnd(gnd), .vdd(vdd), .A(_2870_), .Y(_2871_) );
AOI21X1 AOI21X1_449 ( .gnd(gnd), .vdd(vdd), .A(_2596_), .B(_2594_), .C(_2597_), .Y(_2872_) );
NAND2X1 NAND2X1_366 ( .gnd(gnd), .vdd(vdd), .A(_2872_), .B(_2871_), .Y(_2873_) );
NOR2X1 NOR2X1_582 ( .gnd(gnd), .vdd(vdd), .A(_2872_), .B(_2871_), .Y(_2874_) );
INVX1 INVX1_223 ( .gnd(gnd), .vdd(vdd), .A(_2874_), .Y(_2875_) );
NAND3X1 NAND3X1_113 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe12), .B(_2873_), .C(_2875_), .Y(_2876_) );
OAI21X1 OAI21X1_785 ( .gnd(gnd), .vdd(vdd), .A(_2869_), .B(micro_hash_ucr_pipe12), .C(_2876_), .Y(_2877_) );
XNOR2X1 XNOR2X1_70 ( .gnd(gnd), .vdd(vdd), .A(_2857__bF_buf2), .B(micro_hash_ucr_Wx_28_), .Y(_2878_) );
AOI21X1 AOI21X1_450 ( .gnd(gnd), .vdd(vdd), .A(_2605_), .B(_2603_), .C(_2607_), .Y(_2879_) );
INVX1 INVX1_224 ( .gnd(gnd), .vdd(vdd), .A(_2879_), .Y(_2880_) );
AND2X2 AND2X2_220 ( .gnd(gnd), .vdd(vdd), .A(_2880_), .B(_2878_), .Y(_2881_) );
NOR2X1 NOR2X1_583 ( .gnd(gnd), .vdd(vdd), .A(_2878_), .B(_2880_), .Y(_2882_) );
OAI21X1 OAI21X1_786 ( .gnd(gnd), .vdd(vdd), .A(_2881_), .B(_2882_), .C(micro_hash_ucr_pipe14_bF_buf4), .Y(_2883_) );
OAI21X1 OAI21X1_787 ( .gnd(gnd), .vdd(vdd), .A(_2877_), .B(micro_hash_ucr_pipe14_bF_buf3), .C(_2883_), .Y(_2884_) );
AND2X2 AND2X2_221 ( .gnd(gnd), .vdd(vdd), .A(_2884_), .B(_930__bF_buf2), .Y(_2885_) );
XNOR2X1 XNOR2X1_71 ( .gnd(gnd), .vdd(vdd), .A(_2857__bF_buf1), .B(micro_hash_ucr_Wx_36_), .Y(_2886_) );
INVX1 INVX1_225 ( .gnd(gnd), .vdd(vdd), .A(_2886_), .Y(_2887_) );
AOI21X1 AOI21X1_451 ( .gnd(gnd), .vdd(vdd), .A(_2615_), .B(_2613_), .C(_2616_), .Y(_2888_) );
NAND2X1 NAND2X1_367 ( .gnd(gnd), .vdd(vdd), .A(_2887_), .B(_2888_), .Y(_2889_) );
NOR2X1 NOR2X1_584 ( .gnd(gnd), .vdd(vdd), .A(_2887_), .B(_2888_), .Y(_2890_) );
INVX1 INVX1_226 ( .gnd(gnd), .vdd(vdd), .A(_2890_), .Y(_2891_) );
AOI21X1 AOI21X1_452 ( .gnd(gnd), .vdd(vdd), .A(_2889_), .B(_2891_), .C(_930__bF_buf1), .Y(_2892_) );
OAI21X1 OAI21X1_788 ( .gnd(gnd), .vdd(vdd), .A(_2885_), .B(_2892_), .C(_925__bF_buf3), .Y(_2893_) );
XOR2X1 XOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(_2857__bF_buf0), .B(micro_hash_ucr_Wx_44_), .Y(_2894_) );
AOI21X1 AOI21X1_453 ( .gnd(gnd), .vdd(vdd), .A(_2625_), .B(_2623_), .C(_2626_), .Y(_2895_) );
NOR2X1 NOR2X1_585 ( .gnd(gnd), .vdd(vdd), .A(_2894_), .B(_2895_), .Y(_2896_) );
AND2X2 AND2X2_222 ( .gnd(gnd), .vdd(vdd), .A(_2895_), .B(_2894_), .Y(_2897_) );
OAI21X1 OAI21X1_789 ( .gnd(gnd), .vdd(vdd), .A(_2897_), .B(_2896_), .C(micro_hash_ucr_pipe18_bF_buf3), .Y(_2898_) );
NAND2X1 NAND2X1_368 ( .gnd(gnd), .vdd(vdd), .A(_2898_), .B(_2893_), .Y(_2899_) );
XNOR2X1 XNOR2X1_72 ( .gnd(gnd), .vdd(vdd), .A(_2857__bF_buf5), .B(micro_hash_ucr_Wx_52_), .Y(_2900_) );
INVX1 INVX1_227 ( .gnd(gnd), .vdd(vdd), .A(_2900_), .Y(_2901_) );
AOI21X1 AOI21X1_454 ( .gnd(gnd), .vdd(vdd), .A(_2635_), .B(_2633_), .C(_2636_), .Y(_2902_) );
NAND2X1 NAND2X1_369 ( .gnd(gnd), .vdd(vdd), .A(_2901_), .B(_2902_), .Y(_2903_) );
NOR2X1 NOR2X1_586 ( .gnd(gnd), .vdd(vdd), .A(_2901_), .B(_2902_), .Y(_2904_) );
INVX1 INVX1_228 ( .gnd(gnd), .vdd(vdd), .A(_2904_), .Y(_2905_) );
NAND3X1 NAND3X1_114 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe20_bF_buf0), .B(_2903_), .C(_2905_), .Y(_2906_) );
OAI21X1 OAI21X1_790 ( .gnd(gnd), .vdd(vdd), .A(_2899_), .B(micro_hash_ucr_pipe20_bF_buf4), .C(_2906_), .Y(_2907_) );
XNOR2X1 XNOR2X1_73 ( .gnd(gnd), .vdd(vdd), .A(_2857__bF_buf4), .B(micro_hash_ucr_Wx_60_), .Y(_2908_) );
INVX1 INVX1_229 ( .gnd(gnd), .vdd(vdd), .A(_2908_), .Y(_2909_) );
AOI21X1 AOI21X1_455 ( .gnd(gnd), .vdd(vdd), .A(_2642_), .B(_2641_), .C(_2644_), .Y(_2910_) );
NAND2X1 NAND2X1_370 ( .gnd(gnd), .vdd(vdd), .A(_2909_), .B(_2910_), .Y(_2911_) );
NOR2X1 NOR2X1_587 ( .gnd(gnd), .vdd(vdd), .A(_2909_), .B(_2910_), .Y(_2912_) );
INVX1 INVX1_230 ( .gnd(gnd), .vdd(vdd), .A(_2912_), .Y(_2913_) );
NAND2X1 NAND2X1_371 ( .gnd(gnd), .vdd(vdd), .A(_2911_), .B(_2913_), .Y(_2914_) );
OAI21X1 OAI21X1_791 ( .gnd(gnd), .vdd(vdd), .A(_2914_), .B(_924__bF_buf1), .C(_919__bF_buf4), .Y(_2915_) );
AOI21X1 AOI21X1_456 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf0), .B(_2907_), .C(_2915_), .Y(_2916_) );
XNOR2X1 XNOR2X1_74 ( .gnd(gnd), .vdd(vdd), .A(_2857__bF_buf3), .B(micro_hash_ucr_Wx_68_), .Y(_2917_) );
AOI21X1 AOI21X1_457 ( .gnd(gnd), .vdd(vdd), .A(_2650_), .B(_2649_), .C(_2651_), .Y(_2918_) );
INVX1 INVX1_231 ( .gnd(gnd), .vdd(vdd), .A(_2918_), .Y(_2919_) );
NOR2X1 NOR2X1_588 ( .gnd(gnd), .vdd(vdd), .A(_2917_), .B(_2919_), .Y(_2920_) );
NAND2X1 NAND2X1_372 ( .gnd(gnd), .vdd(vdd), .A(_2917_), .B(_2919_), .Y(_2921_) );
INVX1 INVX1_232 ( .gnd(gnd), .vdd(vdd), .A(_2921_), .Y(_2922_) );
OAI21X1 OAI21X1_792 ( .gnd(gnd), .vdd(vdd), .A(_2922_), .B(_2920_), .C(micro_hash_ucr_pipe24_bF_buf2), .Y(_2923_) );
NAND2X1 NAND2X1_373 ( .gnd(gnd), .vdd(vdd), .A(_920__bF_buf0), .B(_2923_), .Y(_2924_) );
NOR2X1 NOR2X1_589 ( .gnd(gnd), .vdd(vdd), .A(_2924_), .B(_2916_), .Y(_2925_) );
XNOR2X1 XNOR2X1_75 ( .gnd(gnd), .vdd(vdd), .A(_2857__bF_buf2), .B(micro_hash_ucr_Wx_76_), .Y(_2926_) );
INVX1 INVX1_233 ( .gnd(gnd), .vdd(vdd), .A(_2926_), .Y(_2927_) );
AOI21X1 AOI21X1_458 ( .gnd(gnd), .vdd(vdd), .A(_2658_), .B(_2657_), .C(_2659_), .Y(_2928_) );
NOR2X1 NOR2X1_590 ( .gnd(gnd), .vdd(vdd), .A(_2927_), .B(_2928_), .Y(_2929_) );
INVX1 INVX1_234 ( .gnd(gnd), .vdd(vdd), .A(_2929_), .Y(_2930_) );
AOI21X1 AOI21X1_459 ( .gnd(gnd), .vdd(vdd), .A(_2927_), .B(_2928_), .C(_920__bF_buf4), .Y(_2931_) );
AOI21X1 AOI21X1_460 ( .gnd(gnd), .vdd(vdd), .A(_2930_), .B(_2931_), .C(_2925_), .Y(_2932_) );
XNOR2X1 XNOR2X1_76 ( .gnd(gnd), .vdd(vdd), .A(_2857__bF_buf1), .B(micro_hash_ucr_Wx_84_), .Y(_2933_) );
INVX1 INVX1_235 ( .gnd(gnd), .vdd(vdd), .A(_2933_), .Y(_2934_) );
AOI21X1 AOI21X1_461 ( .gnd(gnd), .vdd(vdd), .A(_2667_), .B(_2666_), .C(_2668_), .Y(_2935_) );
NAND2X1 NAND2X1_374 ( .gnd(gnd), .vdd(vdd), .A(_2934_), .B(_2935_), .Y(_2936_) );
NOR2X1 NOR2X1_591 ( .gnd(gnd), .vdd(vdd), .A(_2934_), .B(_2935_), .Y(_2937_) );
INVX1 INVX1_236 ( .gnd(gnd), .vdd(vdd), .A(_2937_), .Y(_2938_) );
NAND3X1 NAND3X1_115 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe28_bF_buf1), .B(_2936_), .C(_2938_), .Y(_2939_) );
OAI21X1 OAI21X1_793 ( .gnd(gnd), .vdd(vdd), .A(_2932_), .B(micro_hash_ucr_pipe28_bF_buf0), .C(_2939_), .Y(_2940_) );
XNOR2X1 XNOR2X1_77 ( .gnd(gnd), .vdd(vdd), .A(_2857__bF_buf0), .B(micro_hash_ucr_Wx_92_), .Y(_2941_) );
INVX1 INVX1_237 ( .gnd(gnd), .vdd(vdd), .A(_2941_), .Y(_2942_) );
AOI21X1 AOI21X1_462 ( .gnd(gnd), .vdd(vdd), .A(_2674_), .B(_2673_), .C(_2676_), .Y(_2943_) );
NOR2X1 NOR2X1_592 ( .gnd(gnd), .vdd(vdd), .A(_2942_), .B(_2943_), .Y(_2944_) );
INVX1 INVX1_238 ( .gnd(gnd), .vdd(vdd), .A(_2944_), .Y(_2945_) );
AOI21X1 AOI21X1_463 ( .gnd(gnd), .vdd(vdd), .A(_2942_), .B(_2943_), .C(_913__bF_buf2), .Y(_2946_) );
AOI22X1 AOI22X1_30 ( .gnd(gnd), .vdd(vdd), .A(_2945_), .B(_2946_), .C(_2940_), .D(_913__bF_buf1), .Y(_2947_) );
NAND2X1 NAND2X1_375 ( .gnd(gnd), .vdd(vdd), .A(_914__bF_buf3), .B(_2947_), .Y(_2948_) );
XNOR2X1 XNOR2X1_78 ( .gnd(gnd), .vdd(vdd), .A(_2857__bF_buf5), .B(micro_hash_ucr_Wx_100_), .Y(_2949_) );
INVX1 INVX1_239 ( .gnd(gnd), .vdd(vdd), .A(_2949_), .Y(_2950_) );
AOI21X1 AOI21X1_464 ( .gnd(gnd), .vdd(vdd), .A(_2683_), .B(_2682_), .C(_2684_), .Y(_2951_) );
AND2X2 AND2X2_223 ( .gnd(gnd), .vdd(vdd), .A(_2951_), .B(_2950_), .Y(_2952_) );
NOR2X1 NOR2X1_593 ( .gnd(gnd), .vdd(vdd), .A(_2950_), .B(_2951_), .Y(_2953_) );
OAI21X1 OAI21X1_794 ( .gnd(gnd), .vdd(vdd), .A(_2952_), .B(_2953_), .C(micro_hash_ucr_pipe32_bF_buf2), .Y(_2954_) );
AOI21X1 AOI21X1_465 ( .gnd(gnd), .vdd(vdd), .A(_2954_), .B(_2948_), .C(micro_hash_ucr_pipe34_bF_buf1), .Y(_2955_) );
XNOR2X1 XNOR2X1_79 ( .gnd(gnd), .vdd(vdd), .A(_2857__bF_buf4), .B(micro_hash_ucr_Wx_108_), .Y(_2956_) );
INVX1 INVX1_240 ( .gnd(gnd), .vdd(vdd), .A(_2956_), .Y(_2957_) );
AOI21X1 AOI21X1_466 ( .gnd(gnd), .vdd(vdd), .A(_2691_), .B(_2690_), .C(_2692_), .Y(_2958_) );
NAND2X1 NAND2X1_376 ( .gnd(gnd), .vdd(vdd), .A(_2957_), .B(_2958_), .Y(_2959_) );
NOR2X1 NOR2X1_594 ( .gnd(gnd), .vdd(vdd), .A(_2957_), .B(_2958_), .Y(_2960_) );
INVX1 INVX1_241 ( .gnd(gnd), .vdd(vdd), .A(_2960_), .Y(_2961_) );
AOI21X1 AOI21X1_467 ( .gnd(gnd), .vdd(vdd), .A(_2959_), .B(_2961_), .C(_912__bF_buf3), .Y(_2962_) );
OAI21X1 OAI21X1_795 ( .gnd(gnd), .vdd(vdd), .A(_2955_), .B(_2962_), .C(_907__bF_buf2), .Y(_2963_) );
XNOR2X1 XNOR2X1_80 ( .gnd(gnd), .vdd(vdd), .A(_2857__bF_buf3), .B(_518_), .Y(_2964_) );
AOI21X1 AOI21X1_468 ( .gnd(gnd), .vdd(vdd), .A(_2700_), .B(_2699_), .C(_2701_), .Y(_2965_) );
AND2X2 AND2X2_224 ( .gnd(gnd), .vdd(vdd), .A(_2965_), .B(_2964_), .Y(_2966_) );
NOR2X1 NOR2X1_595 ( .gnd(gnd), .vdd(vdd), .A(_2964_), .B(_2965_), .Y(_2967_) );
OAI21X1 OAI21X1_796 ( .gnd(gnd), .vdd(vdd), .A(_2966_), .B(_2967_), .C(micro_hash_ucr_pipe36_bF_buf1), .Y(_2968_) );
NAND3X1 NAND3X1_116 ( .gnd(gnd), .vdd(vdd), .A(_908__bF_buf0), .B(_2968_), .C(_2963_), .Y(_2969_) );
XNOR2X1 XNOR2X1_81 ( .gnd(gnd), .vdd(vdd), .A(_2857__bF_buf2), .B(micro_hash_ucr_Wx_124_), .Y(_2970_) );
INVX1 INVX1_242 ( .gnd(gnd), .vdd(vdd), .A(_2970_), .Y(_2971_) );
AOI21X1 AOI21X1_469 ( .gnd(gnd), .vdd(vdd), .A(_2707_), .B(_2706_), .C(_2708_), .Y(_2972_) );
NOR2X1 NOR2X1_596 ( .gnd(gnd), .vdd(vdd), .A(_2971_), .B(_2972_), .Y(_2973_) );
INVX1 INVX1_243 ( .gnd(gnd), .vdd(vdd), .A(_2973_), .Y(_2974_) );
NAND2X1 NAND2X1_377 ( .gnd(gnd), .vdd(vdd), .A(_2971_), .B(_2972_), .Y(_2975_) );
NAND2X1 NAND2X1_378 ( .gnd(gnd), .vdd(vdd), .A(_2975_), .B(_2974_), .Y(_2976_) );
OAI21X1 OAI21X1_797 ( .gnd(gnd), .vdd(vdd), .A(_908__bF_buf4), .B(_2976_), .C(_2969_), .Y(_2977_) );
NOR2X1 NOR2X1_597 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe40_bF_buf4), .B(_2977_), .Y(_2978_) );
XNOR2X1 XNOR2X1_82 ( .gnd(gnd), .vdd(vdd), .A(_2857__bF_buf1), .B(micro_hash_ucr_Wx_132_), .Y(_2979_) );
INVX1 INVX1_244 ( .gnd(gnd), .vdd(vdd), .A(_2979_), .Y(_2980_) );
AOI21X1 AOI21X1_470 ( .gnd(gnd), .vdd(vdd), .A(_2716_), .B(_2715_), .C(_2717_), .Y(_2981_) );
NAND2X1 NAND2X1_379 ( .gnd(gnd), .vdd(vdd), .A(_2980_), .B(_2981_), .Y(_2982_) );
NOR2X1 NOR2X1_598 ( .gnd(gnd), .vdd(vdd), .A(_2980_), .B(_2981_), .Y(_2983_) );
INVX1 INVX1_245 ( .gnd(gnd), .vdd(vdd), .A(_2983_), .Y(_2984_) );
AOI21X1 AOI21X1_471 ( .gnd(gnd), .vdd(vdd), .A(_2982_), .B(_2984_), .C(_906__bF_buf4), .Y(_2985_) );
OAI21X1 OAI21X1_798 ( .gnd(gnd), .vdd(vdd), .A(_2978_), .B(_2985_), .C(_901__bF_buf0), .Y(_2986_) );
XNOR2X1 XNOR2X1_83 ( .gnd(gnd), .vdd(vdd), .A(_2857__bF_buf0), .B(micro_hash_ucr_Wx_140_), .Y(_2987_) );
INVX1 INVX1_246 ( .gnd(gnd), .vdd(vdd), .A(_2987_), .Y(_2988_) );
AOI21X1 AOI21X1_472 ( .gnd(gnd), .vdd(vdd), .A(_2724_), .B(_2723_), .C(_2725_), .Y(_2989_) );
AND2X2 AND2X2_225 ( .gnd(gnd), .vdd(vdd), .A(_2989_), .B(_2988_), .Y(_2990_) );
NOR2X1 NOR2X1_599 ( .gnd(gnd), .vdd(vdd), .A(_2988_), .B(_2989_), .Y(_2991_) );
OAI21X1 OAI21X1_799 ( .gnd(gnd), .vdd(vdd), .A(_2990_), .B(_2991_), .C(micro_hash_ucr_pipe42_bF_buf3), .Y(_2992_) );
NAND3X1 NAND3X1_117 ( .gnd(gnd), .vdd(vdd), .A(_902__bF_buf2), .B(_2992_), .C(_2986_), .Y(_2993_) );
XNOR2X1 XNOR2X1_84 ( .gnd(gnd), .vdd(vdd), .A(_2857__bF_buf5), .B(micro_hash_ucr_Wx_148_), .Y(_2994_) );
INVX1 INVX1_247 ( .gnd(gnd), .vdd(vdd), .A(_2994_), .Y(_2995_) );
AOI21X1 AOI21X1_473 ( .gnd(gnd), .vdd(vdd), .A(_2732_), .B(_2731_), .C(_2733_), .Y(_2996_) );
NOR2X1 NOR2X1_600 ( .gnd(gnd), .vdd(vdd), .A(_2995_), .B(_2996_), .Y(_2997_) );
INVX1 INVX1_248 ( .gnd(gnd), .vdd(vdd), .A(_2997_), .Y(_2998_) );
NAND2X1 NAND2X1_380 ( .gnd(gnd), .vdd(vdd), .A(_2995_), .B(_2996_), .Y(_2999_) );
NAND2X1 NAND2X1_381 ( .gnd(gnd), .vdd(vdd), .A(_2999_), .B(_2998_), .Y(_3000_) );
OAI21X1 OAI21X1_800 ( .gnd(gnd), .vdd(vdd), .A(_902__bF_buf1), .B(_3000_), .C(_2993_), .Y(_3001_) );
NOR2X1 NOR2X1_601 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe46_bF_buf1), .B(_3001_), .Y(_3002_) );
XNOR2X1 XNOR2X1_85 ( .gnd(gnd), .vdd(vdd), .A(_2857__bF_buf4), .B(micro_hash_ucr_Wx_156_), .Y(_3003_) );
INVX1 INVX1_249 ( .gnd(gnd), .vdd(vdd), .A(_3003_), .Y(_3004_) );
AOI21X1 AOI21X1_474 ( .gnd(gnd), .vdd(vdd), .A(_2740_), .B(_2739_), .C(_2742_), .Y(_3005_) );
NAND2X1 NAND2X1_382 ( .gnd(gnd), .vdd(vdd), .A(_3005_), .B(_3004_), .Y(_3006_) );
NOR2X1 NOR2X1_602 ( .gnd(gnd), .vdd(vdd), .A(_3005_), .B(_3004_), .Y(_3007_) );
INVX1 INVX1_250 ( .gnd(gnd), .vdd(vdd), .A(_3007_), .Y(_3008_) );
AOI21X1 AOI21X1_475 ( .gnd(gnd), .vdd(vdd), .A(_3006_), .B(_3008_), .C(_900__bF_buf2), .Y(_3009_) );
OAI21X1 OAI21X1_801 ( .gnd(gnd), .vdd(vdd), .A(_3002_), .B(_3009_), .C(_895__bF_buf0), .Y(_3010_) );
XNOR2X1 XNOR2X1_86 ( .gnd(gnd), .vdd(vdd), .A(_2857__bF_buf3), .B(micro_hash_ucr_Wx_164_), .Y(_3011_) );
INVX1 INVX1_251 ( .gnd(gnd), .vdd(vdd), .A(_3011_), .Y(_3012_) );
AOI21X1 AOI21X1_476 ( .gnd(gnd), .vdd(vdd), .A(_2748_), .B(_2747_), .C(_2749_), .Y(_3013_) );
AND2X2 AND2X2_226 ( .gnd(gnd), .vdd(vdd), .A(_3013_), .B(_3012_), .Y(_3014_) );
NOR2X1 NOR2X1_603 ( .gnd(gnd), .vdd(vdd), .A(_3012_), .B(_3013_), .Y(_3015_) );
OAI21X1 OAI21X1_802 ( .gnd(gnd), .vdd(vdd), .A(_3014_), .B(_3015_), .C(micro_hash_ucr_pipe48_bF_buf3), .Y(_3016_) );
NAND3X1 NAND3X1_118 ( .gnd(gnd), .vdd(vdd), .A(_896__bF_buf3), .B(_3016_), .C(_3010_), .Y(_3017_) );
XNOR2X1 XNOR2X1_87 ( .gnd(gnd), .vdd(vdd), .A(_2857__bF_buf2), .B(micro_hash_ucr_Wx_172_), .Y(_3018_) );
INVX1 INVX1_252 ( .gnd(gnd), .vdd(vdd), .A(_3018_), .Y(_3019_) );
AOI21X1 AOI21X1_477 ( .gnd(gnd), .vdd(vdd), .A(_2756_), .B(_2755_), .C(_2757_), .Y(_3020_) );
OR2X2 OR2X2_33 ( .gnd(gnd), .vdd(vdd), .A(_3020_), .B(_3019_), .Y(_3021_) );
NAND2X1 NAND2X1_383 ( .gnd(gnd), .vdd(vdd), .A(_3019_), .B(_3020_), .Y(_3022_) );
NAND2X1 NAND2X1_384 ( .gnd(gnd), .vdd(vdd), .A(_3022_), .B(_3021_), .Y(_3023_) );
OAI21X1 OAI21X1_803 ( .gnd(gnd), .vdd(vdd), .A(_896__bF_buf2), .B(_3023_), .C(_3017_), .Y(_3024_) );
XNOR2X1 XNOR2X1_88 ( .gnd(gnd), .vdd(vdd), .A(_2857__bF_buf1), .B(_599_), .Y(_3025_) );
AOI21X1 AOI21X1_478 ( .gnd(gnd), .vdd(vdd), .A(_2764_), .B(_2763_), .C(_2765_), .Y(_3026_) );
AND2X2 AND2X2_227 ( .gnd(gnd), .vdd(vdd), .A(_3026_), .B(_3025_), .Y(_3027_) );
NOR2X1 NOR2X1_604 ( .gnd(gnd), .vdd(vdd), .A(_3025_), .B(_3026_), .Y(_3028_) );
OAI21X1 OAI21X1_804 ( .gnd(gnd), .vdd(vdd), .A(_3027_), .B(_3028_), .C(micro_hash_ucr_pipe52_bF_buf0), .Y(_3029_) );
OAI21X1 OAI21X1_805 ( .gnd(gnd), .vdd(vdd), .A(_3024_), .B(micro_hash_ucr_pipe52_bF_buf4), .C(_3029_), .Y(_3030_) );
NAND2X1 NAND2X1_385 ( .gnd(gnd), .vdd(vdd), .A(_889__bF_buf4), .B(_3030_), .Y(_3031_) );
XNOR2X1 XNOR2X1_89 ( .gnd(gnd), .vdd(vdd), .A(_2857__bF_buf0), .B(micro_hash_ucr_Wx_188_), .Y(_3032_) );
INVX1 INVX1_253 ( .gnd(gnd), .vdd(vdd), .A(_3032_), .Y(_3033_) );
AOI21X1 AOI21X1_479 ( .gnd(gnd), .vdd(vdd), .A(_2772_), .B(_2771_), .C(_2774_), .Y(_3034_) );
AND2X2 AND2X2_228 ( .gnd(gnd), .vdd(vdd), .A(_3034_), .B(_3033_), .Y(_3035_) );
NOR2X1 NOR2X1_605 ( .gnd(gnd), .vdd(vdd), .A(_3033_), .B(_3034_), .Y(_3036_) );
OAI21X1 OAI21X1_806 ( .gnd(gnd), .vdd(vdd), .A(_3035_), .B(_3036_), .C(micro_hash_ucr_pipe54_bF_buf3), .Y(_3037_) );
AND2X2 AND2X2_229 ( .gnd(gnd), .vdd(vdd), .A(_3037_), .B(_890__bF_buf1), .Y(_3038_) );
XNOR2X1 XNOR2X1_90 ( .gnd(gnd), .vdd(vdd), .A(_2857__bF_buf5), .B(micro_hash_ucr_Wx_196_), .Y(_3039_) );
INVX1 INVX1_254 ( .gnd(gnd), .vdd(vdd), .A(_3039_), .Y(_3040_) );
AOI21X1 AOI21X1_480 ( .gnd(gnd), .vdd(vdd), .A(_2780_), .B(_2779_), .C(_2781_), .Y(_3041_) );
NOR2X1 NOR2X1_606 ( .gnd(gnd), .vdd(vdd), .A(_3040_), .B(_3041_), .Y(_3042_) );
INVX1 INVX1_255 ( .gnd(gnd), .vdd(vdd), .A(_3042_), .Y(_3043_) );
AOI21X1 AOI21X1_481 ( .gnd(gnd), .vdd(vdd), .A(_3040_), .B(_3041_), .C(_890__bF_buf0), .Y(_3044_) );
AOI22X1 AOI22X1_31 ( .gnd(gnd), .vdd(vdd), .A(_3043_), .B(_3044_), .C(_3031_), .D(_3038_), .Y(_3045_) );
XNOR2X1 XNOR2X1_91 ( .gnd(gnd), .vdd(vdd), .A(_2857__bF_buf4), .B(micro_hash_ucr_Wx_204_), .Y(_3046_) );
INVX1 INVX1_256 ( .gnd(gnd), .vdd(vdd), .A(_3046_), .Y(_3047_) );
AOI21X1 AOI21X1_482 ( .gnd(gnd), .vdd(vdd), .A(_2788_), .B(_2787_), .C(_2789_), .Y(_3048_) );
NAND2X1 NAND2X1_386 ( .gnd(gnd), .vdd(vdd), .A(_3047_), .B(_3048_), .Y(_3049_) );
NOR2X1 NOR2X1_607 ( .gnd(gnd), .vdd(vdd), .A(_3047_), .B(_3048_), .Y(_3050_) );
NOR2X1 NOR2X1_608 ( .gnd(gnd), .vdd(vdd), .A(_888__bF_buf2), .B(_3050_), .Y(_3051_) );
AOI21X1 AOI21X1_483 ( .gnd(gnd), .vdd(vdd), .A(_3049_), .B(_3051_), .C(micro_hash_ucr_pipe60_bF_buf0), .Y(_3052_) );
OAI21X1 OAI21X1_807 ( .gnd(gnd), .vdd(vdd), .A(_3045_), .B(micro_hash_ucr_pipe58_bF_buf2), .C(_3052_), .Y(_3053_) );
XOR2X1 XOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_2857__bF_buf3), .B(micro_hash_ucr_Wx_212_), .Y(_3054_) );
AOI21X1 AOI21X1_484 ( .gnd(gnd), .vdd(vdd), .A(_2797_), .B(_2796_), .C(_2798_), .Y(_3055_) );
AND2X2 AND2X2_230 ( .gnd(gnd), .vdd(vdd), .A(_3055_), .B(_3054_), .Y(_3056_) );
NOR2X1 NOR2X1_609 ( .gnd(gnd), .vdd(vdd), .A(_3054_), .B(_3055_), .Y(_3057_) );
OAI21X1 OAI21X1_808 ( .gnd(gnd), .vdd(vdd), .A(_3056_), .B(_3057_), .C(micro_hash_ucr_pipe60_bF_buf4), .Y(_3058_) );
AND2X2 AND2X2_231 ( .gnd(gnd), .vdd(vdd), .A(_3058_), .B(_884__bF_buf3), .Y(_3059_) );
XNOR2X1 XNOR2X1_92 ( .gnd(gnd), .vdd(vdd), .A(_2857__bF_buf2), .B(micro_hash_ucr_Wx_220_), .Y(_3060_) );
INVX1 INVX1_257 ( .gnd(gnd), .vdd(vdd), .A(_3060_), .Y(_3061_) );
AOI21X1 AOI21X1_485 ( .gnd(gnd), .vdd(vdd), .A(_2804_), .B(_2803_), .C(_2806_), .Y(_3062_) );
NOR2X1 NOR2X1_610 ( .gnd(gnd), .vdd(vdd), .A(_3061_), .B(_3062_), .Y(_3063_) );
INVX1 INVX1_258 ( .gnd(gnd), .vdd(vdd), .A(_3063_), .Y(_3064_) );
AOI21X1 AOI21X1_486 ( .gnd(gnd), .vdd(vdd), .A(_3061_), .B(_3062_), .C(_884__bF_buf2), .Y(_3065_) );
AOI22X1 AOI22X1_32 ( .gnd(gnd), .vdd(vdd), .A(_3064_), .B(_3065_), .C(_3053_), .D(_3059_), .Y(_3066_) );
XNOR2X1 XNOR2X1_93 ( .gnd(gnd), .vdd(vdd), .A(_2857__bF_buf1), .B(micro_hash_ucr_Wx_228_), .Y(_3067_) );
INVX1 INVX1_259 ( .gnd(gnd), .vdd(vdd), .A(_3067_), .Y(_3068_) );
AOI21X1 AOI21X1_487 ( .gnd(gnd), .vdd(vdd), .A(_2814_), .B(_2812_), .C(_2815_), .Y(_3069_) );
NAND2X1 NAND2X1_387 ( .gnd(gnd), .vdd(vdd), .A(_3068_), .B(_3069_), .Y(_3070_) );
NOR2X1 NOR2X1_611 ( .gnd(gnd), .vdd(vdd), .A(_3068_), .B(_3069_), .Y(_3071_) );
NOR2X1 NOR2X1_612 ( .gnd(gnd), .vdd(vdd), .A(_882__bF_buf2), .B(_3071_), .Y(_3072_) );
AOI21X1 AOI21X1_488 ( .gnd(gnd), .vdd(vdd), .A(_3070_), .B(_3072_), .C(micro_hash_ucr_pipe66_bF_buf1), .Y(_3073_) );
OAI21X1 OAI21X1_809 ( .gnd(gnd), .vdd(vdd), .A(_3066_), .B(micro_hash_ucr_pipe64_bF_buf2), .C(_3073_), .Y(_3074_) );
XNOR2X1 XNOR2X1_94 ( .gnd(gnd), .vdd(vdd), .A(_2857__bF_buf0), .B(micro_hash_ucr_Wx_236_), .Y(_3075_) );
INVX1 INVX1_260 ( .gnd(gnd), .vdd(vdd), .A(_3075_), .Y(_3076_) );
AOI21X1 AOI21X1_489 ( .gnd(gnd), .vdd(vdd), .A(_2823_), .B(_2821_), .C(_2824_), .Y(_3077_) );
AND2X2 AND2X2_232 ( .gnd(gnd), .vdd(vdd), .A(_3076_), .B(_3077_), .Y(_3078_) );
NOR2X1 NOR2X1_613 ( .gnd(gnd), .vdd(vdd), .A(_3077_), .B(_3076_), .Y(_3079_) );
OAI21X1 OAI21X1_810 ( .gnd(gnd), .vdd(vdd), .A(_3078_), .B(_3079_), .C(micro_hash_ucr_pipe66_bF_buf0), .Y(_3080_) );
AND2X2 AND2X2_233 ( .gnd(gnd), .vdd(vdd), .A(_3074_), .B(_3080_), .Y(_3081_) );
XNOR2X1 XNOR2X1_95 ( .gnd(gnd), .vdd(vdd), .A(_2857__bF_buf5), .B(micro_hash_ucr_Wx_244_), .Y(_3082_) );
INVX1 INVX1_261 ( .gnd(gnd), .vdd(vdd), .A(_3082_), .Y(_3083_) );
AOI21X1 AOI21X1_490 ( .gnd(gnd), .vdd(vdd), .A(_2833_), .B(_2831_), .C(_2835_), .Y(_3084_) );
AND2X2 AND2X2_234 ( .gnd(gnd), .vdd(vdd), .A(_3084_), .B(_3083_), .Y(_3085_) );
NOR2X1 NOR2X1_614 ( .gnd(gnd), .vdd(vdd), .A(_3083_), .B(_3084_), .Y(_3086_) );
OAI21X1 OAI21X1_811 ( .gnd(gnd), .vdd(vdd), .A(_3085_), .B(_3086_), .C(micro_hash_ucr_pipe68), .Y(_3087_) );
OAI21X1 OAI21X1_812 ( .gnd(gnd), .vdd(vdd), .A(_3081_), .B(micro_hash_ucr_pipe68), .C(_3087_), .Y(_3088_) );
XNOR2X1 XNOR2X1_96 ( .gnd(gnd), .vdd(vdd), .A(_2857__bF_buf4), .B(micro_hash_ucr_Wx_252_), .Y(_3089_) );
AOI21X1 AOI21X1_491 ( .gnd(gnd), .vdd(vdd), .A(_2842_), .B(_2840_), .C(_2844_), .Y(_3090_) );
XNOR2X1 XNOR2X1_97 ( .gnd(gnd), .vdd(vdd), .A(_3090_), .B(_3089_), .Y(_3091_) );
OAI21X1 OAI21X1_813 ( .gnd(gnd), .vdd(vdd), .A(_3091_), .B(_876__bF_buf0), .C(_302__bF_buf1), .Y(_3092_) );
AOI21X1 AOI21X1_492 ( .gnd(gnd), .vdd(vdd), .A(_876__bF_buf3), .B(_3088_), .C(_3092_), .Y(_299__4_) );
INVX2 INVX2_113 ( .gnd(gnd), .vdd(vdd), .A(_369_), .Y(_3093_) );
INVX8 INVX8_92 ( .gnd(gnd), .vdd(vdd), .A(_2857__bF_buf3), .Y(_3094_) );
AOI21X1 AOI21X1_493 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_220_), .B(_3094__bF_buf3), .C(_3063_), .Y(_3095_) );
OAI21X1 OAI21X1_814 ( .gnd(gnd), .vdd(vdd), .A(_2850_), .B(_2851_), .C(_2855_), .Y(_3096_) );
NOR2X1 NOR2X1_615 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_k_5_), .B(micro_hash_ucr_x_5_), .Y(_3097_) );
INVX1 INVX1_262 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_x_5_), .Y(_3098_) );
NOR2X1 NOR2X1_616 ( .gnd(gnd), .vdd(vdd), .A(_1834_), .B(_3098_), .Y(_3099_) );
NOR2X1 NOR2X1_617 ( .gnd(gnd), .vdd(vdd), .A(_3097_), .B(_3099_), .Y(_3100_) );
NAND2X1 NAND2X1_388 ( .gnd(gnd), .vdd(vdd), .A(_3100_), .B(_3096_), .Y(_3101_) );
INVX8 INVX8_93 ( .gnd(gnd), .vdd(vdd), .A(_3101_), .Y(_3102_) );
NOR2X1 NOR2X1_618 ( .gnd(gnd), .vdd(vdd), .A(_3100_), .B(_3096_), .Y(_3103_) );
OAI21X1 OAI21X1_815 ( .gnd(gnd), .vdd(vdd), .A(_3102_), .B(_3103_), .C(_550_), .Y(_3104_) );
INVX1 INVX1_263 ( .gnd(gnd), .vdd(vdd), .A(_3104_), .Y(_3105_) );
NOR2X1 NOR2X1_619 ( .gnd(gnd), .vdd(vdd), .A(_3103_), .B(_3102_), .Y(_3106_) );
INVX8 INVX8_94 ( .gnd(gnd), .vdd(vdd), .A(_3106__bF_buf5), .Y(_3107_) );
NOR2X1 NOR2X1_620 ( .gnd(gnd), .vdd(vdd), .A(_550_), .B(_3107__bF_buf3), .Y(_3108_) );
NOR2X1 NOR2X1_621 ( .gnd(gnd), .vdd(vdd), .A(_3105_), .B(_3108_), .Y(_3109_) );
XNOR2X1 XNOR2X1_98 ( .gnd(gnd), .vdd(vdd), .A(_3095_), .B(_3109_), .Y(_3110_) );
AOI21X1 AOI21X1_494 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_188_), .B(_3094__bF_buf2), .C(_3036_), .Y(_3111_) );
OAI21X1 OAI21X1_816 ( .gnd(gnd), .vdd(vdd), .A(_3102_), .B(_3103_), .C(_660_), .Y(_3112_) );
INVX1 INVX1_264 ( .gnd(gnd), .vdd(vdd), .A(_3112_), .Y(_3113_) );
NOR2X1 NOR2X1_622 ( .gnd(gnd), .vdd(vdd), .A(_660_), .B(_3107__bF_buf2), .Y(_3114_) );
NOR2X1 NOR2X1_623 ( .gnd(gnd), .vdd(vdd), .A(_3113_), .B(_3114_), .Y(_3115_) );
XNOR2X1 XNOR2X1_99 ( .gnd(gnd), .vdd(vdd), .A(_3115_), .B(_3111_), .Y(_3116_) );
OAI21X1 OAI21X1_817 ( .gnd(gnd), .vdd(vdd), .A(_574_), .B(_2857__bF_buf2), .C(_2974_), .Y(_3117_) );
XNOR2X1 XNOR2X1_100 ( .gnd(gnd), .vdd(vdd), .A(_3106__bF_buf4), .B(micro_hash_ucr_Wx_125_), .Y(_3118_) );
XNOR2X1 XNOR2X1_101 ( .gnd(gnd), .vdd(vdd), .A(_3117_), .B(_3118_), .Y(_3119_) );
AOI21X1 AOI21X1_495 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_4_), .B(_3094__bF_buf1), .C(_2861_), .Y(_3120_) );
INVX1 INVX1_265 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_5_), .Y(_3121_) );
OAI21X1 OAI21X1_818 ( .gnd(gnd), .vdd(vdd), .A(_3102_), .B(_3103_), .C(_3121_), .Y(_3122_) );
NAND2X1 NAND2X1_389 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_5_), .B(_3106__bF_buf3), .Y(_3123_) );
NAND2X1 NAND2X1_390 ( .gnd(gnd), .vdd(vdd), .A(_3122_), .B(_3123_), .Y(_3124_) );
XNOR2X1 XNOR2X1_102 ( .gnd(gnd), .vdd(vdd), .A(_3120_), .B(_3124_), .Y(_3125_) );
NOR2X1 NOR2X1_624 ( .gnd(gnd), .vdd(vdd), .A(_4459_), .B(_937_), .Y(_3126_) );
OAI21X1 OAI21X1_819 ( .gnd(gnd), .vdd(vdd), .A(_4460_), .B(micro_hash_ucr_pipe6), .C(_938_), .Y(_3127_) );
OAI21X1 OAI21X1_820 ( .gnd(gnd), .vdd(vdd), .A(_3127_), .B(_3126_), .C(_936_), .Y(_3128_) );
AOI21X1 AOI21X1_496 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe8), .B(_3125_), .C(_3128_), .Y(_3129_) );
NOR2X1 NOR2X1_625 ( .gnd(gnd), .vdd(vdd), .A(_2863_), .B(_2864_), .Y(_3130_) );
AOI21X1 AOI21X1_497 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_12_), .B(_3094__bF_buf0), .C(_3130_), .Y(_3131_) );
XNOR2X1 XNOR2X1_103 ( .gnd(gnd), .vdd(vdd), .A(_3106__bF_buf2), .B(micro_hash_ucr_Wx_13_), .Y(_3132_) );
XNOR2X1 XNOR2X1_104 ( .gnd(gnd), .vdd(vdd), .A(_3132_), .B(_3131_), .Y(_3133_) );
OAI21X1 OAI21X1_821 ( .gnd(gnd), .vdd(vdd), .A(_3133_), .B(_936_), .C(_931_), .Y(_3134_) );
AOI21X1 AOI21X1_498 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_20_), .B(_3094__bF_buf3), .C(_2874_), .Y(_3135_) );
INVX1 INVX1_266 ( .gnd(gnd), .vdd(vdd), .A(_3135_), .Y(_3136_) );
NOR2X1 NOR2X1_626 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_21_), .B(_3106__bF_buf1), .Y(_3137_) );
INVX1 INVX1_267 ( .gnd(gnd), .vdd(vdd), .A(_3137_), .Y(_3138_) );
NAND2X1 NAND2X1_391 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_21_), .B(_3106__bF_buf0), .Y(_3139_) );
NAND2X1 NAND2X1_392 ( .gnd(gnd), .vdd(vdd), .A(_3139_), .B(_3138_), .Y(_3140_) );
AOI21X1 AOI21X1_499 ( .gnd(gnd), .vdd(vdd), .A(_3136_), .B(_3140_), .C(_931_), .Y(_3141_) );
OAI21X1 OAI21X1_822 ( .gnd(gnd), .vdd(vdd), .A(_3136_), .B(_3140_), .C(_3141_), .Y(_3142_) );
OAI21X1 OAI21X1_823 ( .gnd(gnd), .vdd(vdd), .A(_3129_), .B(_3134_), .C(_3142_), .Y(_3143_) );
NAND2X1 NAND2X1_393 ( .gnd(gnd), .vdd(vdd), .A(_932_), .B(_3143_), .Y(_3144_) );
AOI21X1 AOI21X1_500 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_28_), .B(_3094__bF_buf2), .C(_2881_), .Y(_3145_) );
INVX2 INVX2_114 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_29_), .Y(_3146_) );
XNOR2X1 XNOR2X1_105 ( .gnd(gnd), .vdd(vdd), .A(_3106__bF_buf5), .B(_3146_), .Y(_3147_) );
XNOR2X1 XNOR2X1_106 ( .gnd(gnd), .vdd(vdd), .A(_3145_), .B(_3147_), .Y(_3148_) );
OAI21X1 OAI21X1_824 ( .gnd(gnd), .vdd(vdd), .A(_932_), .B(_3148_), .C(_3144_), .Y(_3149_) );
NAND2X1 NAND2X1_394 ( .gnd(gnd), .vdd(vdd), .A(_930__bF_buf0), .B(_3149_), .Y(_3150_) );
AOI21X1 AOI21X1_501 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_36_), .B(_3094__bF_buf1), .C(_2890_), .Y(_3151_) );
INVX2 INVX2_115 ( .gnd(gnd), .vdd(vdd), .A(_3151_), .Y(_3152_) );
INVX1 INVX1_268 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_37_), .Y(_3153_) );
OAI21X1 OAI21X1_825 ( .gnd(gnd), .vdd(vdd), .A(_3102_), .B(_3103_), .C(_3153_), .Y(_3154_) );
NOR2X1 NOR2X1_627 ( .gnd(gnd), .vdd(vdd), .A(_3153_), .B(_3107__bF_buf1), .Y(_3155_) );
INVX1 INVX1_269 ( .gnd(gnd), .vdd(vdd), .A(_3155_), .Y(_3156_) );
NAND2X1 NAND2X1_395 ( .gnd(gnd), .vdd(vdd), .A(_3154_), .B(_3156_), .Y(_3157_) );
AOI21X1 AOI21X1_502 ( .gnd(gnd), .vdd(vdd), .A(_3152_), .B(_3157_), .C(_930__bF_buf4), .Y(_3158_) );
OAI21X1 OAI21X1_826 ( .gnd(gnd), .vdd(vdd), .A(_3152_), .B(_3157_), .C(_3158_), .Y(_3159_) );
AND2X2 AND2X2_235 ( .gnd(gnd), .vdd(vdd), .A(_3159_), .B(_925__bF_buf2), .Y(_3160_) );
AOI21X1 AOI21X1_503 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_44_), .B(_3094__bF_buf0), .C(_2896_), .Y(_3161_) );
NOR2X1 NOR2X1_628 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_45_), .B(_3106__bF_buf4), .Y(_3162_) );
INVX1 INVX1_270 ( .gnd(gnd), .vdd(vdd), .A(_3162_), .Y(_3163_) );
NAND2X1 NAND2X1_396 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_45_), .B(_3106__bF_buf3), .Y(_3164_) );
NAND2X1 NAND2X1_397 ( .gnd(gnd), .vdd(vdd), .A(_3164_), .B(_3163_), .Y(_3165_) );
AND2X2 AND2X2_236 ( .gnd(gnd), .vdd(vdd), .A(_3165_), .B(_3161_), .Y(_3166_) );
OAI21X1 OAI21X1_827 ( .gnd(gnd), .vdd(vdd), .A(_3165_), .B(_3161_), .C(micro_hash_ucr_pipe18_bF_buf2), .Y(_3167_) );
OAI21X1 OAI21X1_828 ( .gnd(gnd), .vdd(vdd), .A(_3166_), .B(_3167_), .C(_926__bF_buf1), .Y(_3168_) );
AOI21X1 AOI21X1_504 ( .gnd(gnd), .vdd(vdd), .A(_3160_), .B(_3150_), .C(_3168_), .Y(_3169_) );
AOI21X1 AOI21X1_505 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_52_), .B(_3094__bF_buf3), .C(_2904_), .Y(_3170_) );
INVX1 INVX1_271 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_53_), .Y(_3171_) );
OAI21X1 OAI21X1_829 ( .gnd(gnd), .vdd(vdd), .A(_3102_), .B(_3103_), .C(_3171_), .Y(_3172_) );
INVX1 INVX1_272 ( .gnd(gnd), .vdd(vdd), .A(_3172_), .Y(_3173_) );
NOR2X1 NOR2X1_629 ( .gnd(gnd), .vdd(vdd), .A(_3171_), .B(_3107__bF_buf0), .Y(_3174_) );
NOR2X1 NOR2X1_630 ( .gnd(gnd), .vdd(vdd), .A(_3173_), .B(_3174_), .Y(_3175_) );
XNOR2X1 XNOR2X1_107 ( .gnd(gnd), .vdd(vdd), .A(_3170_), .B(_3175_), .Y(_3176_) );
OAI21X1 OAI21X1_830 ( .gnd(gnd), .vdd(vdd), .A(_3176_), .B(_926__bF_buf0), .C(_924__bF_buf4), .Y(_3177_) );
OAI21X1 OAI21X1_831 ( .gnd(gnd), .vdd(vdd), .A(_819_), .B(_2857__bF_buf1), .C(_2913_), .Y(_3178_) );
XNOR2X1 XNOR2X1_108 ( .gnd(gnd), .vdd(vdd), .A(_3106__bF_buf2), .B(micro_hash_ucr_Wx_61_), .Y(_3179_) );
XNOR2X1 XNOR2X1_109 ( .gnd(gnd), .vdd(vdd), .A(_3178_), .B(_3179_), .Y(_3180_) );
AOI21X1 AOI21X1_506 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe22_bF_buf0), .B(_3180_), .C(micro_hash_ucr_pipe24_bF_buf1), .Y(_3181_) );
OAI21X1 OAI21X1_832 ( .gnd(gnd), .vdd(vdd), .A(_3169_), .B(_3177_), .C(_3181_), .Y(_3182_) );
OAI21X1 OAI21X1_833 ( .gnd(gnd), .vdd(vdd), .A(_865_), .B(_2857__bF_buf0), .C(_2921_), .Y(_3183_) );
OAI21X1 OAI21X1_834 ( .gnd(gnd), .vdd(vdd), .A(_3102_), .B(_3103_), .C(_868_), .Y(_3184_) );
NOR2X1 NOR2X1_631 ( .gnd(gnd), .vdd(vdd), .A(_868_), .B(_3107__bF_buf3), .Y(_3185_) );
INVX1 INVX1_273 ( .gnd(gnd), .vdd(vdd), .A(_3185_), .Y(_3186_) );
NAND2X1 NAND2X1_398 ( .gnd(gnd), .vdd(vdd), .A(_3184_), .B(_3186_), .Y(_3187_) );
AOI21X1 AOI21X1_507 ( .gnd(gnd), .vdd(vdd), .A(_3183_), .B(_3187_), .C(_919__bF_buf3), .Y(_3188_) );
OAI21X1 OAI21X1_835 ( .gnd(gnd), .vdd(vdd), .A(_3183_), .B(_3187_), .C(_3188_), .Y(_3189_) );
AND2X2 AND2X2_237 ( .gnd(gnd), .vdd(vdd), .A(_3189_), .B(_920__bF_buf3), .Y(_3190_) );
OAI21X1 OAI21X1_836 ( .gnd(gnd), .vdd(vdd), .A(_841_), .B(_2857__bF_buf5), .C(_2930_), .Y(_3191_) );
INVX2 INVX2_116 ( .gnd(gnd), .vdd(vdd), .A(_3191_), .Y(_3192_) );
XNOR2X1 XNOR2X1_110 ( .gnd(gnd), .vdd(vdd), .A(_3106__bF_buf1), .B(micro_hash_ucr_Wx_77_), .Y(_3193_) );
AND2X2 AND2X2_238 ( .gnd(gnd), .vdd(vdd), .A(_3192_), .B(_3193_), .Y(_3194_) );
OAI21X1 OAI21X1_837 ( .gnd(gnd), .vdd(vdd), .A(_3192_), .B(_3193_), .C(micro_hash_ucr_pipe26_bF_buf3), .Y(_3195_) );
OAI21X1 OAI21X1_838 ( .gnd(gnd), .vdd(vdd), .A(_3194_), .B(_3195_), .C(_918__bF_buf3), .Y(_3196_) );
AOI21X1 AOI21X1_508 ( .gnd(gnd), .vdd(vdd), .A(_3190_), .B(_3182_), .C(_3196_), .Y(_3197_) );
OAI21X1 OAI21X1_839 ( .gnd(gnd), .vdd(vdd), .A(_752_), .B(_2857__bF_buf4), .C(_2938_), .Y(_3198_) );
XNOR2X1 XNOR2X1_111 ( .gnd(gnd), .vdd(vdd), .A(_3106__bF_buf0), .B(micro_hash_ucr_Wx_85_), .Y(_3199_) );
XNOR2X1 XNOR2X1_112 ( .gnd(gnd), .vdd(vdd), .A(_3198_), .B(_3199_), .Y(_3200_) );
OAI21X1 OAI21X1_840 ( .gnd(gnd), .vdd(vdd), .A(_3200_), .B(_918__bF_buf2), .C(_913__bF_buf0), .Y(_3201_) );
OAI21X1 OAI21X1_841 ( .gnd(gnd), .vdd(vdd), .A(_794_), .B(_2857__bF_buf3), .C(_2945_), .Y(_3202_) );
OAI21X1 OAI21X1_842 ( .gnd(gnd), .vdd(vdd), .A(_3102_), .B(_3103_), .C(_797_), .Y(_3203_) );
INVX1 INVX1_274 ( .gnd(gnd), .vdd(vdd), .A(_3203_), .Y(_3204_) );
NOR2X1 NOR2X1_632 ( .gnd(gnd), .vdd(vdd), .A(_797_), .B(_3107__bF_buf2), .Y(_3205_) );
NOR2X1 NOR2X1_633 ( .gnd(gnd), .vdd(vdd), .A(_3204_), .B(_3205_), .Y(_3206_) );
XOR2X1 XOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(_3202_), .B(_3206_), .Y(_3207_) );
AOI21X1 AOI21X1_509 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe30_bF_buf1), .B(_3207_), .C(micro_hash_ucr_pipe32_bF_buf1), .Y(_3208_) );
OAI21X1 OAI21X1_843 ( .gnd(gnd), .vdd(vdd), .A(_3197_), .B(_3201_), .C(_3208_), .Y(_3209_) );
AOI21X1 AOI21X1_510 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_100_), .B(_3094__bF_buf2), .C(_2953_), .Y(_3210_) );
XNOR2X1 XNOR2X1_113 ( .gnd(gnd), .vdd(vdd), .A(_3106__bF_buf5), .B(micro_hash_ucr_Wx_101_), .Y(_3211_) );
XNOR2X1 XNOR2X1_114 ( .gnd(gnd), .vdd(vdd), .A(_3210_), .B(_3211_), .Y(_3212_) );
AOI21X1 AOI21X1_511 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe32_bF_buf0), .B(_3212_), .C(micro_hash_ucr_pipe34_bF_buf0), .Y(_3213_) );
OAI21X1 OAI21X1_844 ( .gnd(gnd), .vdd(vdd), .A(_684_), .B(_2857__bF_buf2), .C(_2961_), .Y(_3214_) );
OAI21X1 OAI21X1_845 ( .gnd(gnd), .vdd(vdd), .A(_3102_), .B(_3103_), .C(_687_), .Y(_3215_) );
NOR2X1 NOR2X1_634 ( .gnd(gnd), .vdd(vdd), .A(_687_), .B(_3107__bF_buf1), .Y(_3216_) );
INVX1 INVX1_275 ( .gnd(gnd), .vdd(vdd), .A(_3216_), .Y(_3217_) );
NAND2X1 NAND2X1_399 ( .gnd(gnd), .vdd(vdd), .A(_3215_), .B(_3217_), .Y(_3218_) );
XOR2X1 XOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(_3214_), .B(_3218_), .Y(_3219_) );
OAI21X1 OAI21X1_846 ( .gnd(gnd), .vdd(vdd), .A(_3219_), .B(_912__bF_buf2), .C(_907__bF_buf1), .Y(_3220_) );
AOI21X1 AOI21X1_512 ( .gnd(gnd), .vdd(vdd), .A(_3213_), .B(_3209_), .C(_3220_), .Y(_3221_) );
AOI21X1 AOI21X1_513 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_116_), .B(_3094__bF_buf1), .C(_2967_), .Y(_3222_) );
NOR2X1 NOR2X1_635 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_117_), .B(_3106__bF_buf4), .Y(_3223_) );
NOR2X1 NOR2X1_636 ( .gnd(gnd), .vdd(vdd), .A(_521_), .B(_3107__bF_buf0), .Y(_3224_) );
NOR2X1 NOR2X1_637 ( .gnd(gnd), .vdd(vdd), .A(_3223_), .B(_3224_), .Y(_3225_) );
OAI21X1 OAI21X1_847 ( .gnd(gnd), .vdd(vdd), .A(_3225_), .B(_3222_), .C(micro_hash_ucr_pipe36_bF_buf0), .Y(_3226_) );
AOI21X1 AOI21X1_514 ( .gnd(gnd), .vdd(vdd), .A(_3222_), .B(_3225_), .C(_3226_), .Y(_3227_) );
OAI21X1 OAI21X1_848 ( .gnd(gnd), .vdd(vdd), .A(_3221_), .B(_3227_), .C(_908__bF_buf3), .Y(_3228_) );
OAI21X1 OAI21X1_849 ( .gnd(gnd), .vdd(vdd), .A(_908__bF_buf2), .B(_3119_), .C(_3228_), .Y(_3229_) );
NAND2X1 NAND2X1_400 ( .gnd(gnd), .vdd(vdd), .A(_906__bF_buf3), .B(_3229_), .Y(_3230_) );
OAI21X1 OAI21X1_850 ( .gnd(gnd), .vdd(vdd), .A(_546_), .B(_2857__bF_buf1), .C(_2984_), .Y(_3231_) );
OAI21X1 OAI21X1_851 ( .gnd(gnd), .vdd(vdd), .A(_3102_), .B(_3103_), .C(_549_), .Y(_3232_) );
NOR2X1 NOR2X1_638 ( .gnd(gnd), .vdd(vdd), .A(_549_), .B(_3107__bF_buf3), .Y(_3233_) );
INVX1 INVX1_276 ( .gnd(gnd), .vdd(vdd), .A(_3233_), .Y(_3234_) );
NAND2X1 NAND2X1_401 ( .gnd(gnd), .vdd(vdd), .A(_3232_), .B(_3234_), .Y(_3235_) );
AOI21X1 AOI21X1_515 ( .gnd(gnd), .vdd(vdd), .A(_3231_), .B(_3235_), .C(_906__bF_buf2), .Y(_3236_) );
OAI21X1 OAI21X1_852 ( .gnd(gnd), .vdd(vdd), .A(_3231_), .B(_3235_), .C(_3236_), .Y(_3237_) );
AND2X2 AND2X2_239 ( .gnd(gnd), .vdd(vdd), .A(_3237_), .B(_901__bF_buf4), .Y(_3238_) );
AOI21X1 AOI21X1_516 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_140_), .B(_3094__bF_buf0), .C(_2991_), .Y(_3239_) );
OAI21X1 OAI21X1_853 ( .gnd(gnd), .vdd(vdd), .A(_3102_), .B(_3103_), .C(_798_), .Y(_3240_) );
NAND2X1 NAND2X1_402 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_141_), .B(_3106__bF_buf3), .Y(_3241_) );
NAND2X1 NAND2X1_403 ( .gnd(gnd), .vdd(vdd), .A(_3240_), .B(_3241_), .Y(_3242_) );
AND2X2 AND2X2_240 ( .gnd(gnd), .vdd(vdd), .A(_3239_), .B(_3242_), .Y(_3243_) );
OAI21X1 OAI21X1_854 ( .gnd(gnd), .vdd(vdd), .A(_3239_), .B(_3242_), .C(micro_hash_ucr_pipe42_bF_buf2), .Y(_3244_) );
OAI21X1 OAI21X1_855 ( .gnd(gnd), .vdd(vdd), .A(_3243_), .B(_3244_), .C(_902__bF_buf0), .Y(_3245_) );
AOI21X1 AOI21X1_517 ( .gnd(gnd), .vdd(vdd), .A(_3238_), .B(_3230_), .C(_3245_), .Y(_3246_) );
OAI21X1 OAI21X1_856 ( .gnd(gnd), .vdd(vdd), .A(_627_), .B(_2857__bF_buf0), .C(_2998_), .Y(_3247_) );
OAI21X1 OAI21X1_857 ( .gnd(gnd), .vdd(vdd), .A(_3102_), .B(_3103_), .C(_630_), .Y(_3248_) );
NOR2X1 NOR2X1_639 ( .gnd(gnd), .vdd(vdd), .A(_630_), .B(_3107__bF_buf2), .Y(_3249_) );
INVX1 INVX1_277 ( .gnd(gnd), .vdd(vdd), .A(_3249_), .Y(_3250_) );
NAND2X1 NAND2X1_404 ( .gnd(gnd), .vdd(vdd), .A(_3248_), .B(_3250_), .Y(_3251_) );
XNOR2X1 XNOR2X1_115 ( .gnd(gnd), .vdd(vdd), .A(_3247_), .B(_3251_), .Y(_3252_) );
OAI21X1 OAI21X1_858 ( .gnd(gnd), .vdd(vdd), .A(_3252_), .B(_902__bF_buf4), .C(_900__bF_buf1), .Y(_3253_) );
AOI21X1 AOI21X1_518 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_156_), .B(_3094__bF_buf3), .C(_3007_), .Y(_3254_) );
NOR2X1 NOR2X1_640 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_157_), .B(_3106__bF_buf2), .Y(_3255_) );
INVX1 INVX1_278 ( .gnd(gnd), .vdd(vdd), .A(_3255_), .Y(_3256_) );
NAND2X1 NAND2X1_405 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_157_), .B(_3106__bF_buf1), .Y(_3257_) );
NAND2X1 NAND2X1_406 ( .gnd(gnd), .vdd(vdd), .A(_3257_), .B(_3256_), .Y(_3258_) );
XOR2X1 XOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(_3258_), .B(_3254_), .Y(_3259_) );
AOI21X1 AOI21X1_519 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe46_bF_buf0), .B(_3259_), .C(micro_hash_ucr_pipe48_bF_buf2), .Y(_3260_) );
OAI21X1 OAI21X1_859 ( .gnd(gnd), .vdd(vdd), .A(_3246_), .B(_3253_), .C(_3260_), .Y(_3261_) );
AOI21X1 AOI21X1_520 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_164_), .B(_3094__bF_buf2), .C(_3015_), .Y(_3262_) );
NOR2X1 NOR2X1_641 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_165_), .B(_3106__bF_buf0), .Y(_3263_) );
INVX1 INVX1_279 ( .gnd(gnd), .vdd(vdd), .A(_3263_), .Y(_3264_) );
NAND2X1 NAND2X1_407 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_165_), .B(_3106__bF_buf5), .Y(_3265_) );
NAND2X1 NAND2X1_408 ( .gnd(gnd), .vdd(vdd), .A(_3265_), .B(_3264_), .Y(_3266_) );
XNOR2X1 XNOR2X1_116 ( .gnd(gnd), .vdd(vdd), .A(_3262_), .B(_3266_), .Y(_3267_) );
AOI21X1 AOI21X1_521 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe48_bF_buf1), .B(_3267_), .C(micro_hash_ucr_pipe50_bF_buf0), .Y(_3268_) );
OAI21X1 OAI21X1_860 ( .gnd(gnd), .vdd(vdd), .A(_708_), .B(_2857__bF_buf5), .C(_3021_), .Y(_3269_) );
OAI21X1 OAI21X1_861 ( .gnd(gnd), .vdd(vdd), .A(_3102_), .B(_3103_), .C(_711_), .Y(_3270_) );
NOR2X1 NOR2X1_642 ( .gnd(gnd), .vdd(vdd), .A(_711_), .B(_3107__bF_buf1), .Y(_3271_) );
INVX1 INVX1_280 ( .gnd(gnd), .vdd(vdd), .A(_3271_), .Y(_3272_) );
NAND2X1 NAND2X1_409 ( .gnd(gnd), .vdd(vdd), .A(_3270_), .B(_3272_), .Y(_3273_) );
XOR2X1 XOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(_3273_), .B(_3269_), .Y(_3274_) );
OAI21X1 OAI21X1_862 ( .gnd(gnd), .vdd(vdd), .A(_3274_), .B(_896__bF_buf1), .C(_894__bF_buf3), .Y(_3275_) );
AOI21X1 AOI21X1_522 ( .gnd(gnd), .vdd(vdd), .A(_3268_), .B(_3261_), .C(_3275_), .Y(_3276_) );
AOI21X1 AOI21X1_523 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_180_), .B(_3094__bF_buf1), .C(_3028_), .Y(_3277_) );
NOR2X1 NOR2X1_643 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_181_), .B(_3106__bF_buf4), .Y(_3278_) );
NOR2X1 NOR2X1_644 ( .gnd(gnd), .vdd(vdd), .A(_602_), .B(_3107__bF_buf0), .Y(_3279_) );
NOR2X1 NOR2X1_645 ( .gnd(gnd), .vdd(vdd), .A(_3278_), .B(_3279_), .Y(_3280_) );
OAI21X1 OAI21X1_863 ( .gnd(gnd), .vdd(vdd), .A(_3277_), .B(_3280_), .C(micro_hash_ucr_pipe52_bF_buf3), .Y(_3281_) );
AOI21X1 AOI21X1_524 ( .gnd(gnd), .vdd(vdd), .A(_3277_), .B(_3280_), .C(_3281_), .Y(_3282_) );
OAI21X1 OAI21X1_864 ( .gnd(gnd), .vdd(vdd), .A(_3276_), .B(_3282_), .C(_889__bF_buf3), .Y(_3283_) );
OAI21X1 OAI21X1_865 ( .gnd(gnd), .vdd(vdd), .A(_889__bF_buf2), .B(_3116_), .C(_3283_), .Y(_3284_) );
NAND2X1 NAND2X1_410 ( .gnd(gnd), .vdd(vdd), .A(_890__bF_buf4), .B(_3284_), .Y(_3285_) );
AOI21X1 AOI21X1_525 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_196_), .B(_3094__bF_buf0), .C(_3042_), .Y(_3286_) );
NOR2X1 NOR2X1_646 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_197_), .B(_3106__bF_buf3), .Y(_3287_) );
INVX1 INVX1_281 ( .gnd(gnd), .vdd(vdd), .A(_3287_), .Y(_3288_) );
NAND2X1 NAND2X1_411 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_197_), .B(_3106__bF_buf2), .Y(_3289_) );
NAND2X1 NAND2X1_412 ( .gnd(gnd), .vdd(vdd), .A(_3289_), .B(_3288_), .Y(_3290_) );
XNOR2X1 XNOR2X1_117 ( .gnd(gnd), .vdd(vdd), .A(_3286_), .B(_3290_), .Y(_3291_) );
AOI21X1 AOI21X1_526 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe56_bF_buf2), .B(_3291_), .C(micro_hash_ucr_pipe58_bF_buf1), .Y(_3292_) );
AOI21X1 AOI21X1_527 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_204_), .B(_3094__bF_buf3), .C(_3050_), .Y(_3293_) );
NOR2X1 NOR2X1_647 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_205_), .B(_3106__bF_buf1), .Y(_3294_) );
INVX1 INVX1_282 ( .gnd(gnd), .vdd(vdd), .A(_3294_), .Y(_3295_) );
NAND2X1 NAND2X1_413 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_205_), .B(_3106__bF_buf0), .Y(_3296_) );
NAND2X1 NAND2X1_414 ( .gnd(gnd), .vdd(vdd), .A(_3296_), .B(_3295_), .Y(_3297_) );
AND2X2 AND2X2_241 ( .gnd(gnd), .vdd(vdd), .A(_3293_), .B(_3297_), .Y(_3298_) );
OAI21X1 OAI21X1_866 ( .gnd(gnd), .vdd(vdd), .A(_3293_), .B(_3297_), .C(micro_hash_ucr_pipe58_bF_buf0), .Y(_3299_) );
OAI21X1 OAI21X1_867 ( .gnd(gnd), .vdd(vdd), .A(_3298_), .B(_3299_), .C(_883__bF_buf0), .Y(_3300_) );
AOI21X1 AOI21X1_528 ( .gnd(gnd), .vdd(vdd), .A(_3292_), .B(_3285_), .C(_3300_), .Y(_3301_) );
AOI21X1 AOI21X1_529 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_212_), .B(_3094__bF_buf2), .C(_3057_), .Y(_3302_) );
NOR2X1 NOR2X1_648 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_213_), .B(_3106__bF_buf5), .Y(_3303_) );
NAND2X1 NAND2X1_415 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_213_), .B(_3106__bF_buf4), .Y(_3304_) );
INVX1 INVX1_283 ( .gnd(gnd), .vdd(vdd), .A(_3304_), .Y(_3305_) );
NOR2X1 NOR2X1_649 ( .gnd(gnd), .vdd(vdd), .A(_3303_), .B(_3305_), .Y(_3306_) );
OAI21X1 OAI21X1_868 ( .gnd(gnd), .vdd(vdd), .A(_3306_), .B(_3302_), .C(micro_hash_ucr_pipe60_bF_buf3), .Y(_3307_) );
AOI21X1 AOI21X1_530 ( .gnd(gnd), .vdd(vdd), .A(_3302_), .B(_3306_), .C(_3307_), .Y(_3308_) );
OAI21X1 OAI21X1_869 ( .gnd(gnd), .vdd(vdd), .A(_3301_), .B(_3308_), .C(_884__bF_buf1), .Y(_3309_) );
OAI21X1 OAI21X1_870 ( .gnd(gnd), .vdd(vdd), .A(_884__bF_buf0), .B(_3110_), .C(_3309_), .Y(_3310_) );
NAND2X1 NAND2X1_416 ( .gnd(gnd), .vdd(vdd), .A(_882__bF_buf1), .B(_3310_), .Y(_3311_) );
AOI21X1 AOI21X1_531 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_228_), .B(_3094__bF_buf1), .C(_3071_), .Y(_3312_) );
NOR2X1 NOR2X1_650 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_229_), .B(_3106__bF_buf3), .Y(_3313_) );
INVX1 INVX1_284 ( .gnd(gnd), .vdd(vdd), .A(_3313_), .Y(_3314_) );
NAND2X1 NAND2X1_417 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_229_), .B(_3106__bF_buf2), .Y(_3315_) );
NAND2X1 NAND2X1_418 ( .gnd(gnd), .vdd(vdd), .A(_3315_), .B(_3314_), .Y(_3316_) );
XNOR2X1 XNOR2X1_118 ( .gnd(gnd), .vdd(vdd), .A(_3316_), .B(_3312_), .Y(_3317_) );
AOI21X1 AOI21X1_532 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe64_bF_buf1), .B(_3317_), .C(micro_hash_ucr_pipe66_bF_buf4), .Y(_3318_) );
AOI21X1 AOI21X1_533 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_236_), .B(_3094__bF_buf0), .C(_3079_), .Y(_3319_) );
NOR2X1 NOR2X1_651 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_237_), .B(_3106__bF_buf1), .Y(_3320_) );
INVX1 INVX1_285 ( .gnd(gnd), .vdd(vdd), .A(_3320_), .Y(_3321_) );
NAND2X1 NAND2X1_419 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_237_), .B(_3106__bF_buf0), .Y(_3322_) );
NAND2X1 NAND2X1_420 ( .gnd(gnd), .vdd(vdd), .A(_3322_), .B(_3321_), .Y(_3323_) );
AND2X2 AND2X2_242 ( .gnd(gnd), .vdd(vdd), .A(_3323_), .B(_3319_), .Y(_3324_) );
OAI21X1 OAI21X1_871 ( .gnd(gnd), .vdd(vdd), .A(_3323_), .B(_3319_), .C(micro_hash_ucr_pipe66_bF_buf3), .Y(_3325_) );
OAI21X1 OAI21X1_872 ( .gnd(gnd), .vdd(vdd), .A(_3324_), .B(_3325_), .C(_878__bF_buf4), .Y(_3326_) );
AOI21X1 AOI21X1_534 ( .gnd(gnd), .vdd(vdd), .A(_3318_), .B(_3311_), .C(_3326_), .Y(_3327_) );
AOI21X1 AOI21X1_535 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_244_), .B(_3094__bF_buf3), .C(_3086_), .Y(_3328_) );
INVX1 INVX1_286 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_245_), .Y(_3329_) );
OAI21X1 OAI21X1_873 ( .gnd(gnd), .vdd(vdd), .A(_3102_), .B(_3103_), .C(_3329_), .Y(_3330_) );
INVX1 INVX1_287 ( .gnd(gnd), .vdd(vdd), .A(_3330_), .Y(_3331_) );
NOR2X1 NOR2X1_652 ( .gnd(gnd), .vdd(vdd), .A(_3329_), .B(_3107__bF_buf3), .Y(_3332_) );
NOR2X1 NOR2X1_653 ( .gnd(gnd), .vdd(vdd), .A(_3331_), .B(_3332_), .Y(_3333_) );
AND2X2 AND2X2_243 ( .gnd(gnd), .vdd(vdd), .A(_3333_), .B(_3328_), .Y(_3334_) );
OAI21X1 OAI21X1_874 ( .gnd(gnd), .vdd(vdd), .A(_3333_), .B(_3328_), .C(micro_hash_ucr_pipe68), .Y(_3335_) );
OAI21X1 OAI21X1_875 ( .gnd(gnd), .vdd(vdd), .A(_3334_), .B(_3335_), .C(_1949_), .Y(_3336_) );
NAND2X1 NAND2X1_421 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_252_), .B(_3094__bF_buf2), .Y(_3337_) );
INVX1 INVX1_288 ( .gnd(gnd), .vdd(vdd), .A(_3089_), .Y(_3338_) );
OAI21X1 OAI21X1_876 ( .gnd(gnd), .vdd(vdd), .A(_3090_), .B(_3338_), .C(_3337_), .Y(_3339_) );
INVX1 INVX1_289 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_253_), .Y(_3340_) );
OAI21X1 OAI21X1_877 ( .gnd(gnd), .vdd(vdd), .A(_3102_), .B(_3103_), .C(_3340_), .Y(_3341_) );
NOR2X1 NOR2X1_654 ( .gnd(gnd), .vdd(vdd), .A(_3340_), .B(_3107__bF_buf2), .Y(_3342_) );
INVX1 INVX1_290 ( .gnd(gnd), .vdd(vdd), .A(_3342_), .Y(_3343_) );
NAND2X1 NAND2X1_422 ( .gnd(gnd), .vdd(vdd), .A(_3341_), .B(_3343_), .Y(_3344_) );
XOR2X1 XOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(_3344_), .B(_3339_), .Y(_3345_) );
OAI22X1 OAI22X1_53 ( .gnd(gnd), .vdd(vdd), .A(_3093_), .B(_3345_), .C(_3327_), .D(_3336_), .Y(_299__5_) );
OAI21X1 OAI21X1_878 ( .gnd(gnd), .vdd(vdd), .A(_1834_), .B(_3098_), .C(_3101_), .Y(_3346_) );
XOR2X1 XOR2X1_61 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_k_6_), .B(micro_hash_ucr_x_6_), .Y(_3347_) );
NOR2X1 NOR2X1_655 ( .gnd(gnd), .vdd(vdd), .A(_3347_), .B(_3346_), .Y(_3348_) );
OAI21X1 OAI21X1_879 ( .gnd(gnd), .vdd(vdd), .A(_3102_), .B(_3099_), .C(_3347_), .Y(_3349_) );
INVX4 INVX4_56 ( .gnd(gnd), .vdd(vdd), .A(_3349_), .Y(_3350_) );
NOR2X1 NOR2X1_656 ( .gnd(gnd), .vdd(vdd), .A(_3348_), .B(_3350_), .Y(_3351_) );
INVX8 INVX8_95 ( .gnd(gnd), .vdd(vdd), .A(_3351__bF_buf4), .Y(_3352_) );
NOR2X1 NOR2X1_657 ( .gnd(gnd), .vdd(vdd), .A(_605_), .B(_3352__bF_buf4), .Y(_3353_) );
INVX1 INVX1_291 ( .gnd(gnd), .vdd(vdd), .A(_3353_), .Y(_3354_) );
OAI21X1 OAI21X1_880 ( .gnd(gnd), .vdd(vdd), .A(_3350_), .B(_3348_), .C(_605_), .Y(_3355_) );
NAND2X1 NAND2X1_423 ( .gnd(gnd), .vdd(vdd), .A(_3355_), .B(_3354_), .Y(_3356_) );
INVX1 INVX1_292 ( .gnd(gnd), .vdd(vdd), .A(_3279_), .Y(_3357_) );
OAI21X1 OAI21X1_881 ( .gnd(gnd), .vdd(vdd), .A(_3277_), .B(_3278_), .C(_3357_), .Y(_3358_) );
XOR2X1 XOR2X1_62 ( .gnd(gnd), .vdd(vdd), .A(_3356_), .B(_3358_), .Y(_3359_) );
NAND2X1 NAND2X1_424 ( .gnd(gnd), .vdd(vdd), .A(H_22_), .B(micro_hash_ucr_pipe6), .Y(_3360_) );
OAI21X1 OAI21X1_882 ( .gnd(gnd), .vdd(vdd), .A(_4472_), .B(micro_hash_ucr_pipe6), .C(_3360_), .Y(_3361_) );
XNOR2X1 XNOR2X1_119 ( .gnd(gnd), .vdd(vdd), .A(_3351__bF_buf3), .B(micro_hash_ucr_Wx_6_), .Y(_3362_) );
INVX1 INVX1_293 ( .gnd(gnd), .vdd(vdd), .A(_3362_), .Y(_3363_) );
INVX1 INVX1_294 ( .gnd(gnd), .vdd(vdd), .A(_3122_), .Y(_3364_) );
OAI21X1 OAI21X1_883 ( .gnd(gnd), .vdd(vdd), .A(_3120_), .B(_3364_), .C(_3123_), .Y(_3365_) );
NOR2X1 NOR2X1_658 ( .gnd(gnd), .vdd(vdd), .A(_3365_), .B(_3363_), .Y(_3366_) );
AND2X2 AND2X2_244 ( .gnd(gnd), .vdd(vdd), .A(_3363_), .B(_3365_), .Y(_3367_) );
OAI21X1 OAI21X1_884 ( .gnd(gnd), .vdd(vdd), .A(_3367_), .B(_3366_), .C(micro_hash_ucr_pipe8), .Y(_3368_) );
OAI21X1 OAI21X1_885 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe8), .B(_3361_), .C(_3368_), .Y(_3369_) );
INVX2 INVX2_117 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_14_), .Y(_3370_) );
XNOR2X1 XNOR2X1_120 ( .gnd(gnd), .vdd(vdd), .A(_3351__bF_buf2), .B(_3370_), .Y(_3371_) );
INVX1 INVX1_295 ( .gnd(gnd), .vdd(vdd), .A(_3371_), .Y(_3372_) );
INVX1 INVX1_296 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_13_), .Y(_3373_) );
OAI21X1 OAI21X1_886 ( .gnd(gnd), .vdd(vdd), .A(_3373_), .B(_3107__bF_buf1), .C(_3131_), .Y(_3374_) );
OAI21X1 OAI21X1_887 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_13_), .B(_3106__bF_buf5), .C(_3374_), .Y(_3375_) );
NAND2X1 NAND2X1_425 ( .gnd(gnd), .vdd(vdd), .A(_3375_), .B(_3372_), .Y(_3376_) );
OR2X2 OR2X2_34 ( .gnd(gnd), .vdd(vdd), .A(_3372_), .B(_3375_), .Y(_3377_) );
NAND3X1 NAND3X1_119 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe10), .B(_3376_), .C(_3377_), .Y(_3378_) );
OAI21X1 OAI21X1_888 ( .gnd(gnd), .vdd(vdd), .A(_3369_), .B(micro_hash_ucr_pipe10), .C(_3378_), .Y(_3379_) );
INVX2 INVX2_118 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_22_), .Y(_3380_) );
XNOR2X1 XNOR2X1_121 ( .gnd(gnd), .vdd(vdd), .A(_3351__bF_buf1), .B(_3380_), .Y(_3381_) );
OAI21X1 OAI21X1_889 ( .gnd(gnd), .vdd(vdd), .A(_3135_), .B(_3137_), .C(_3139_), .Y(_3382_) );
XOR2X1 XOR2X1_63 ( .gnd(gnd), .vdd(vdd), .A(_3381_), .B(_3382_), .Y(_3383_) );
MUX2X1 MUX2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_3379_), .B(_3383_), .S(_931_), .Y(_3384_) );
INVX2 INVX2_119 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_30_), .Y(_3385_) );
XNOR2X1 XNOR2X1_122 ( .gnd(gnd), .vdd(vdd), .A(_3351__bF_buf0), .B(_3385_), .Y(_3386_) );
INVX1 INVX1_297 ( .gnd(gnd), .vdd(vdd), .A(_3386_), .Y(_3387_) );
OAI21X1 OAI21X1_890 ( .gnd(gnd), .vdd(vdd), .A(_3146_), .B(_3107__bF_buf0), .C(_3145_), .Y(_3388_) );
OAI21X1 OAI21X1_891 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_29_), .B(_3106__bF_buf4), .C(_3388_), .Y(_3389_) );
NAND2X1 NAND2X1_426 ( .gnd(gnd), .vdd(vdd), .A(_3389_), .B(_3387_), .Y(_3390_) );
OR2X2 OR2X2_35 ( .gnd(gnd), .vdd(vdd), .A(_3387_), .B(_3389_), .Y(_3391_) );
NAND3X1 NAND3X1_120 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe14_bF_buf2), .B(_3390_), .C(_3391_), .Y(_3392_) );
OAI21X1 OAI21X1_892 ( .gnd(gnd), .vdd(vdd), .A(_3384_), .B(micro_hash_ucr_pipe14_bF_buf1), .C(_3392_), .Y(_3393_) );
NAND2X1 NAND2X1_427 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_38_), .B(_3351__bF_buf4), .Y(_3394_) );
INVX1 INVX1_298 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_38_), .Y(_3395_) );
OAI21X1 OAI21X1_893 ( .gnd(gnd), .vdd(vdd), .A(_3350_), .B(_3348_), .C(_3395_), .Y(_3396_) );
AND2X2 AND2X2_245 ( .gnd(gnd), .vdd(vdd), .A(_3394_), .B(_3396_), .Y(_3397_) );
AOI21X1 AOI21X1_536 ( .gnd(gnd), .vdd(vdd), .A(_3154_), .B(_3152_), .C(_3155_), .Y(_3398_) );
XNOR2X1 XNOR2X1_123 ( .gnd(gnd), .vdd(vdd), .A(_3398_), .B(_3397_), .Y(_3399_) );
MUX2X1 MUX2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_3393_), .B(_3399_), .S(_930__bF_buf3), .Y(_3400_) );
INVX2 INVX2_120 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_46_), .Y(_3401_) );
XNOR2X1 XNOR2X1_124 ( .gnd(gnd), .vdd(vdd), .A(_3351__bF_buf3), .B(_3401_), .Y(_3402_) );
OAI21X1 OAI21X1_894 ( .gnd(gnd), .vdd(vdd), .A(_3161_), .B(_3162_), .C(_3164_), .Y(_3403_) );
OR2X2 OR2X2_36 ( .gnd(gnd), .vdd(vdd), .A(_3402_), .B(_3403_), .Y(_3404_) );
NAND2X1 NAND2X1_428 ( .gnd(gnd), .vdd(vdd), .A(_3403_), .B(_3402_), .Y(_3405_) );
NAND3X1 NAND3X1_121 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe18_bF_buf1), .B(_3405_), .C(_3404_), .Y(_3406_) );
OAI21X1 OAI21X1_895 ( .gnd(gnd), .vdd(vdd), .A(_3400_), .B(micro_hash_ucr_pipe18_bF_buf0), .C(_3406_), .Y(_3407_) );
INVX2 INVX2_121 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_54_), .Y(_3408_) );
XNOR2X1 XNOR2X1_125 ( .gnd(gnd), .vdd(vdd), .A(_3351__bF_buf2), .B(_3408_), .Y(_3409_) );
INVX1 INVX1_299 ( .gnd(gnd), .vdd(vdd), .A(_3174_), .Y(_3410_) );
OAI21X1 OAI21X1_896 ( .gnd(gnd), .vdd(vdd), .A(_3170_), .B(_3173_), .C(_3410_), .Y(_3411_) );
NAND2X1 NAND2X1_429 ( .gnd(gnd), .vdd(vdd), .A(_3409_), .B(_3411_), .Y(_3412_) );
INVX1 INVX1_300 ( .gnd(gnd), .vdd(vdd), .A(_3412_), .Y(_3413_) );
OAI21X1 OAI21X1_897 ( .gnd(gnd), .vdd(vdd), .A(_3411_), .B(_3409_), .C(micro_hash_ucr_pipe20_bF_buf3), .Y(_3414_) );
OAI21X1 OAI21X1_898 ( .gnd(gnd), .vdd(vdd), .A(_3413_), .B(_3414_), .C(_924__bF_buf3), .Y(_3415_) );
AOI21X1 AOI21X1_537 ( .gnd(gnd), .vdd(vdd), .A(_926__bF_buf4), .B(_3407_), .C(_3415_), .Y(_3416_) );
NOR2X1 NOR2X1_659 ( .gnd(gnd), .vdd(vdd), .A(_825_), .B(_3352__bF_buf3), .Y(_3417_) );
INVX1 INVX1_301 ( .gnd(gnd), .vdd(vdd), .A(_3417_), .Y(_3418_) );
OAI21X1 OAI21X1_899 ( .gnd(gnd), .vdd(vdd), .A(_3350_), .B(_3348_), .C(_825_), .Y(_3419_) );
NAND2X1 NAND2X1_430 ( .gnd(gnd), .vdd(vdd), .A(_3419_), .B(_3418_), .Y(_3420_) );
OAI21X1 OAI21X1_900 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_61_), .B(_3106__bF_buf3), .C(_3178_), .Y(_3421_) );
OAI21X1 OAI21X1_901 ( .gnd(gnd), .vdd(vdd), .A(_822_), .B(_3107__bF_buf3), .C(_3421_), .Y(_3422_) );
XNOR2X1 XNOR2X1_126 ( .gnd(gnd), .vdd(vdd), .A(_3420_), .B(_3422_), .Y(_3423_) );
OAI21X1 OAI21X1_902 ( .gnd(gnd), .vdd(vdd), .A(_3423_), .B(_924__bF_buf2), .C(_919__bF_buf2), .Y(_3424_) );
XNOR2X1 XNOR2X1_127 ( .gnd(gnd), .vdd(vdd), .A(_3351__bF_buf1), .B(_690_), .Y(_3425_) );
INVX1 INVX1_302 ( .gnd(gnd), .vdd(vdd), .A(_3425_), .Y(_3426_) );
AOI21X1 AOI21X1_538 ( .gnd(gnd), .vdd(vdd), .A(_3184_), .B(_3183_), .C(_3185_), .Y(_3427_) );
NOR2X1 NOR2X1_660 ( .gnd(gnd), .vdd(vdd), .A(_3426_), .B(_3427_), .Y(_3428_) );
INVX1 INVX1_303 ( .gnd(gnd), .vdd(vdd), .A(_3427_), .Y(_3429_) );
OAI21X1 OAI21X1_903 ( .gnd(gnd), .vdd(vdd), .A(_3429_), .B(_3425_), .C(micro_hash_ucr_pipe24_bF_buf0), .Y(_3430_) );
OAI22X1 OAI22X1_54 ( .gnd(gnd), .vdd(vdd), .A(_3428_), .B(_3430_), .C(_3416_), .D(_3424_), .Y(_3431_) );
XNOR2X1 XNOR2X1_128 ( .gnd(gnd), .vdd(vdd), .A(_3351__bF_buf0), .B(micro_hash_ucr_Wx_78_), .Y(_3432_) );
OAI21X1 OAI21X1_904 ( .gnd(gnd), .vdd(vdd), .A(_844_), .B(_3107__bF_buf2), .C(_3192_), .Y(_3433_) );
OAI21X1 OAI21X1_905 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_77_), .B(_3106__bF_buf2), .C(_3433_), .Y(_3434_) );
NAND2X1 NAND2X1_431 ( .gnd(gnd), .vdd(vdd), .A(_3432_), .B(_3434_), .Y(_3435_) );
OR2X2 OR2X2_37 ( .gnd(gnd), .vdd(vdd), .A(_3434_), .B(_3432_), .Y(_3436_) );
NAND2X1 NAND2X1_432 ( .gnd(gnd), .vdd(vdd), .A(_3435_), .B(_3436_), .Y(_3437_) );
OAI21X1 OAI21X1_906 ( .gnd(gnd), .vdd(vdd), .A(_3437_), .B(_920__bF_buf2), .C(_918__bF_buf1), .Y(_3438_) );
AOI21X1 AOI21X1_539 ( .gnd(gnd), .vdd(vdd), .A(_920__bF_buf1), .B(_3431_), .C(_3438_), .Y(_3439_) );
XNOR2X1 XNOR2X1_129 ( .gnd(gnd), .vdd(vdd), .A(_3351__bF_buf4), .B(_758_), .Y(_3440_) );
OAI21X1 OAI21X1_907 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_85_), .B(_3106__bF_buf1), .C(_3198_), .Y(_3441_) );
OAI21X1 OAI21X1_908 ( .gnd(gnd), .vdd(vdd), .A(_755_), .B(_3107__bF_buf1), .C(_3441_), .Y(_3442_) );
XOR2X1 XOR2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_3442_), .B(_3440_), .Y(_3443_) );
OAI21X1 OAI21X1_909 ( .gnd(gnd), .vdd(vdd), .A(_3443_), .B(_918__bF_buf0), .C(_913__bF_buf4), .Y(_3444_) );
XNOR2X1 XNOR2X1_130 ( .gnd(gnd), .vdd(vdd), .A(_3351__bF_buf3), .B(_801_), .Y(_3445_) );
INVX1 INVX1_304 ( .gnd(gnd), .vdd(vdd), .A(_3445_), .Y(_3446_) );
AOI21X1 AOI21X1_540 ( .gnd(gnd), .vdd(vdd), .A(_3203_), .B(_3202_), .C(_3205_), .Y(_3447_) );
OR2X2 OR2X2_38 ( .gnd(gnd), .vdd(vdd), .A(_3447_), .B(_3446_), .Y(_3448_) );
NAND2X1 NAND2X1_433 ( .gnd(gnd), .vdd(vdd), .A(_3446_), .B(_3447_), .Y(_3449_) );
NAND2X1 NAND2X1_434 ( .gnd(gnd), .vdd(vdd), .A(_3449_), .B(_3448_), .Y(_3450_) );
OAI22X1 OAI22X1_55 ( .gnd(gnd), .vdd(vdd), .A(_913__bF_buf3), .B(_3450_), .C(_3439_), .D(_3444_), .Y(_3451_) );
XNOR2X1 XNOR2X1_131 ( .gnd(gnd), .vdd(vdd), .A(_3351__bF_buf2), .B(micro_hash_ucr_Wx_102_), .Y(_3452_) );
OAI21X1 OAI21X1_910 ( .gnd(gnd), .vdd(vdd), .A(_659_), .B(_3107__bF_buf0), .C(_3210_), .Y(_3453_) );
OAI21X1 OAI21X1_911 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_101_), .B(_3106__bF_buf0), .C(_3453_), .Y(_3454_) );
NAND2X1 NAND2X1_435 ( .gnd(gnd), .vdd(vdd), .A(_3452_), .B(_3454_), .Y(_3455_) );
OR2X2 OR2X2_39 ( .gnd(gnd), .vdd(vdd), .A(_3454_), .B(_3452_), .Y(_3456_) );
NAND2X1 NAND2X1_436 ( .gnd(gnd), .vdd(vdd), .A(_3455_), .B(_3456_), .Y(_3457_) );
OAI21X1 OAI21X1_912 ( .gnd(gnd), .vdd(vdd), .A(_3457_), .B(_914__bF_buf2), .C(_912__bF_buf1), .Y(_3458_) );
AOI21X1 AOI21X1_541 ( .gnd(gnd), .vdd(vdd), .A(_914__bF_buf1), .B(_3451_), .C(_3458_), .Y(_3459_) );
XNOR2X1 XNOR2X1_132 ( .gnd(gnd), .vdd(vdd), .A(_3351__bF_buf1), .B(micro_hash_ucr_Wx_110_), .Y(_3460_) );
AOI21X1 AOI21X1_542 ( .gnd(gnd), .vdd(vdd), .A(_3215_), .B(_3214_), .C(_3216_), .Y(_3461_) );
XOR2X1 XOR2X1_65 ( .gnd(gnd), .vdd(vdd), .A(_3461_), .B(_3460_), .Y(_3462_) );
OAI21X1 OAI21X1_913 ( .gnd(gnd), .vdd(vdd), .A(_3462_), .B(_912__bF_buf0), .C(_907__bF_buf0), .Y(_3463_) );
NOR2X1 NOR2X1_661 ( .gnd(gnd), .vdd(vdd), .A(_3463_), .B(_3459_), .Y(_3464_) );
XNOR2X1 XNOR2X1_133 ( .gnd(gnd), .vdd(vdd), .A(_3351__bF_buf0), .B(_524_), .Y(_3465_) );
INVX1 INVX1_305 ( .gnd(gnd), .vdd(vdd), .A(_3224_), .Y(_3466_) );
OAI21X1 OAI21X1_914 ( .gnd(gnd), .vdd(vdd), .A(_3222_), .B(_3223_), .C(_3466_), .Y(_3467_) );
OAI21X1 OAI21X1_915 ( .gnd(gnd), .vdd(vdd), .A(_3465_), .B(_3467_), .C(micro_hash_ucr_pipe36_bF_buf3), .Y(_3468_) );
AOI21X1 AOI21X1_543 ( .gnd(gnd), .vdd(vdd), .A(_3465_), .B(_3467_), .C(_3468_), .Y(_3469_) );
OAI21X1 OAI21X1_916 ( .gnd(gnd), .vdd(vdd), .A(_3464_), .B(_3469_), .C(_908__bF_buf1), .Y(_3470_) );
XNOR2X1 XNOR2X1_134 ( .gnd(gnd), .vdd(vdd), .A(_3351__bF_buf4), .B(_580_), .Y(_3471_) );
OAI21X1 OAI21X1_917 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_125_), .B(_3106__bF_buf5), .C(_3117_), .Y(_3472_) );
OAI21X1 OAI21X1_918 ( .gnd(gnd), .vdd(vdd), .A(_577_), .B(_3107__bF_buf3), .C(_3472_), .Y(_3473_) );
OR2X2 OR2X2_40 ( .gnd(gnd), .vdd(vdd), .A(_3473_), .B(_3471_), .Y(_3474_) );
NAND2X1 NAND2X1_437 ( .gnd(gnd), .vdd(vdd), .A(_3471_), .B(_3473_), .Y(_3475_) );
NAND3X1 NAND3X1_122 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe38_bF_buf3), .B(_3475_), .C(_3474_), .Y(_3476_) );
AOI21X1 AOI21X1_544 ( .gnd(gnd), .vdd(vdd), .A(_3476_), .B(_3470_), .C(micro_hash_ucr_pipe40_bF_buf3), .Y(_3477_) );
XNOR2X1 XNOR2X1_135 ( .gnd(gnd), .vdd(vdd), .A(_3351__bF_buf3), .B(_553_), .Y(_3478_) );
AOI21X1 AOI21X1_545 ( .gnd(gnd), .vdd(vdd), .A(_3232_), .B(_3231_), .C(_3233_), .Y(_3479_) );
INVX1 INVX1_306 ( .gnd(gnd), .vdd(vdd), .A(_3479_), .Y(_3480_) );
NOR2X1 NOR2X1_662 ( .gnd(gnd), .vdd(vdd), .A(_3478_), .B(_3480_), .Y(_3481_) );
NAND2X1 NAND2X1_438 ( .gnd(gnd), .vdd(vdd), .A(_3478_), .B(_3480_), .Y(_3482_) );
NAND2X1 NAND2X1_439 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe40_bF_buf2), .B(_3482_), .Y(_3483_) );
OAI21X1 OAI21X1_919 ( .gnd(gnd), .vdd(vdd), .A(_3483_), .B(_3481_), .C(_901__bF_buf3), .Y(_3484_) );
XNOR2X1 XNOR2X1_136 ( .gnd(gnd), .vdd(vdd), .A(_3351__bF_buf2), .B(_802_), .Y(_3485_) );
INVX1 INVX1_307 ( .gnd(gnd), .vdd(vdd), .A(_3240_), .Y(_3486_) );
OAI21X1 OAI21X1_920 ( .gnd(gnd), .vdd(vdd), .A(_3239_), .B(_3486_), .C(_3241_), .Y(_3487_) );
XOR2X1 XOR2X1_66 ( .gnd(gnd), .vdd(vdd), .A(_3487_), .B(_3485_), .Y(_3488_) );
OAI22X1 OAI22X1_56 ( .gnd(gnd), .vdd(vdd), .A(_901__bF_buf2), .B(_3488_), .C(_3477_), .D(_3484_), .Y(_3489_) );
XNOR2X1 XNOR2X1_137 ( .gnd(gnd), .vdd(vdd), .A(_3351__bF_buf1), .B(_633_), .Y(_3490_) );
INVX1 INVX1_308 ( .gnd(gnd), .vdd(vdd), .A(_3490_), .Y(_3491_) );
AOI21X1 AOI21X1_546 ( .gnd(gnd), .vdd(vdd), .A(_3248_), .B(_3247_), .C(_3249_), .Y(_3492_) );
OR2X2 OR2X2_41 ( .gnd(gnd), .vdd(vdd), .A(_3492_), .B(_3491_), .Y(_3493_) );
NAND2X1 NAND2X1_440 ( .gnd(gnd), .vdd(vdd), .A(_3491_), .B(_3492_), .Y(_3494_) );
AOI21X1 AOI21X1_547 ( .gnd(gnd), .vdd(vdd), .A(_3494_), .B(_3493_), .C(_902__bF_buf3), .Y(_3495_) );
AOI21X1 AOI21X1_548 ( .gnd(gnd), .vdd(vdd), .A(_902__bF_buf2), .B(_3489_), .C(_3495_), .Y(_3496_) );
XNOR2X1 XNOR2X1_138 ( .gnd(gnd), .vdd(vdd), .A(_3351__bF_buf0), .B(_691_), .Y(_3497_) );
OAI21X1 OAI21X1_921 ( .gnd(gnd), .vdd(vdd), .A(_3254_), .B(_3255_), .C(_3257_), .Y(_3498_) );
NOR2X1 NOR2X1_663 ( .gnd(gnd), .vdd(vdd), .A(_3498_), .B(_3497_), .Y(_3499_) );
NAND2X1 NAND2X1_441 ( .gnd(gnd), .vdd(vdd), .A(_3498_), .B(_3497_), .Y(_3500_) );
NAND2X1 NAND2X1_442 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe46_bF_buf4), .B(_3500_), .Y(_3501_) );
OAI21X1 OAI21X1_922 ( .gnd(gnd), .vdd(vdd), .A(_3501_), .B(_3499_), .C(_895__bF_buf4), .Y(_3502_) );
AOI21X1 AOI21X1_549 ( .gnd(gnd), .vdd(vdd), .A(_900__bF_buf0), .B(_3496_), .C(_3502_), .Y(_3503_) );
XNOR2X1 XNOR2X1_139 ( .gnd(gnd), .vdd(vdd), .A(_3351__bF_buf4), .B(_735_), .Y(_3504_) );
OAI21X1 OAI21X1_923 ( .gnd(gnd), .vdd(vdd), .A(_3262_), .B(_3263_), .C(_3265_), .Y(_3505_) );
XOR2X1 XOR2X1_67 ( .gnd(gnd), .vdd(vdd), .A(_3505_), .B(_3504_), .Y(_3506_) );
OAI21X1 OAI21X1_924 ( .gnd(gnd), .vdd(vdd), .A(_3506_), .B(_895__bF_buf3), .C(_896__bF_buf0), .Y(_3507_) );
NOR2X1 NOR2X1_664 ( .gnd(gnd), .vdd(vdd), .A(_3507_), .B(_3503_), .Y(_3508_) );
XNOR2X1 XNOR2X1_140 ( .gnd(gnd), .vdd(vdd), .A(_3351__bF_buf3), .B(micro_hash_ucr_Wx_174_), .Y(_3509_) );
AOI21X1 AOI21X1_550 ( .gnd(gnd), .vdd(vdd), .A(_3270_), .B(_3269_), .C(_3271_), .Y(_3510_) );
OR2X2 OR2X2_42 ( .gnd(gnd), .vdd(vdd), .A(_3510_), .B(_3509_), .Y(_3511_) );
AOI21X1 AOI21X1_551 ( .gnd(gnd), .vdd(vdd), .A(_3509_), .B(_3510_), .C(_896__bF_buf4), .Y(_3512_) );
AND2X2 AND2X2_246 ( .gnd(gnd), .vdd(vdd), .A(_3511_), .B(_3512_), .Y(_3513_) );
OAI21X1 OAI21X1_925 ( .gnd(gnd), .vdd(vdd), .A(_3508_), .B(_3513_), .C(_894__bF_buf2), .Y(_3514_) );
OAI21X1 OAI21X1_926 ( .gnd(gnd), .vdd(vdd), .A(_894__bF_buf1), .B(_3359_), .C(_3514_), .Y(_3515_) );
XNOR2X1 XNOR2X1_141 ( .gnd(gnd), .vdd(vdd), .A(_3351__bF_buf2), .B(_664_), .Y(_3516_) );
INVX1 INVX1_309 ( .gnd(gnd), .vdd(vdd), .A(_3114_), .Y(_3517_) );
OAI21X1 OAI21X1_927 ( .gnd(gnd), .vdd(vdd), .A(_3111_), .B(_3113_), .C(_3517_), .Y(_3518_) );
NAND2X1 NAND2X1_443 ( .gnd(gnd), .vdd(vdd), .A(_3518_), .B(_3516_), .Y(_3519_) );
INVX1 INVX1_310 ( .gnd(gnd), .vdd(vdd), .A(_3519_), .Y(_3520_) );
OAI21X1 OAI21X1_928 ( .gnd(gnd), .vdd(vdd), .A(_3516_), .B(_3518_), .C(micro_hash_ucr_pipe54_bF_buf2), .Y(_3521_) );
OAI21X1 OAI21X1_929 ( .gnd(gnd), .vdd(vdd), .A(_3520_), .B(_3521_), .C(_890__bF_buf3), .Y(_3522_) );
AOI21X1 AOI21X1_552 ( .gnd(gnd), .vdd(vdd), .A(_889__bF_buf1), .B(_3515_), .C(_3522_), .Y(_3523_) );
NOR2X1 NOR2X1_665 ( .gnd(gnd), .vdd(vdd), .A(_634_), .B(_3352__bF_buf2), .Y(_3524_) );
INVX1 INVX1_311 ( .gnd(gnd), .vdd(vdd), .A(_3524_), .Y(_3525_) );
OAI21X1 OAI21X1_930 ( .gnd(gnd), .vdd(vdd), .A(_3350_), .B(_3348_), .C(_634_), .Y(_3526_) );
NAND2X1 NAND2X1_444 ( .gnd(gnd), .vdd(vdd), .A(_3526_), .B(_3525_), .Y(_3527_) );
OAI21X1 OAI21X1_931 ( .gnd(gnd), .vdd(vdd), .A(_3286_), .B(_3287_), .C(_3289_), .Y(_3528_) );
XNOR2X1 XNOR2X1_142 ( .gnd(gnd), .vdd(vdd), .A(_3527_), .B(_3528_), .Y(_3529_) );
OAI21X1 OAI21X1_932 ( .gnd(gnd), .vdd(vdd), .A(_3529_), .B(_890__bF_buf2), .C(_888__bF_buf1), .Y(_3530_) );
XNOR2X1 XNOR2X1_143 ( .gnd(gnd), .vdd(vdd), .A(_3351__bF_buf1), .B(_525_), .Y(_3531_) );
OAI21X1 OAI21X1_933 ( .gnd(gnd), .vdd(vdd), .A(_3293_), .B(_3294_), .C(_3296_), .Y(_3532_) );
XOR2X1 XOR2X1_68 ( .gnd(gnd), .vdd(vdd), .A(_3532_), .B(_3531_), .Y(_3533_) );
AOI21X1 AOI21X1_553 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe58_bF_buf4), .B(_3533_), .C(micro_hash_ucr_pipe60_bF_buf2), .Y(_3534_) );
OAI21X1 OAI21X1_934 ( .gnd(gnd), .vdd(vdd), .A(_3523_), .B(_3530_), .C(_3534_), .Y(_3535_) );
XNOR2X1 XNOR2X1_144 ( .gnd(gnd), .vdd(vdd), .A(_3351__bF_buf0), .B(_581_), .Y(_3536_) );
OAI21X1 OAI21X1_935 ( .gnd(gnd), .vdd(vdd), .A(_3302_), .B(_3303_), .C(_3304_), .Y(_3537_) );
XNOR2X1 XNOR2X1_145 ( .gnd(gnd), .vdd(vdd), .A(_3536_), .B(_3537_), .Y(_3538_) );
AOI21X1 AOI21X1_554 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe60_bF_buf1), .B(_3538_), .C(micro_hash_ucr_pipe62_bF_buf4), .Y(_3539_) );
XNOR2X1 XNOR2X1_146 ( .gnd(gnd), .vdd(vdd), .A(_3351__bF_buf4), .B(_554_), .Y(_3540_) );
INVX1 INVX1_312 ( .gnd(gnd), .vdd(vdd), .A(_3108_), .Y(_3541_) );
OAI21X1 OAI21X1_936 ( .gnd(gnd), .vdd(vdd), .A(_3095_), .B(_3105_), .C(_3541_), .Y(_3542_) );
NAND2X1 NAND2X1_445 ( .gnd(gnd), .vdd(vdd), .A(_3540_), .B(_3542_), .Y(_3543_) );
NOR2X1 NOR2X1_666 ( .gnd(gnd), .vdd(vdd), .A(_3540_), .B(_3542_), .Y(_3544_) );
NOR2X1 NOR2X1_667 ( .gnd(gnd), .vdd(vdd), .A(_884__bF_buf4), .B(_3544_), .Y(_3545_) );
AOI22X1 AOI22X1_33 ( .gnd(gnd), .vdd(vdd), .A(_3543_), .B(_3545_), .C(_3535_), .D(_3539_), .Y(_3546_) );
INVX2 INVX2_122 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_230_), .Y(_3547_) );
XNOR2X1 XNOR2X1_147 ( .gnd(gnd), .vdd(vdd), .A(_3351__bF_buf3), .B(_3547_), .Y(_3548_) );
OAI21X1 OAI21X1_937 ( .gnd(gnd), .vdd(vdd), .A(_3312_), .B(_3313_), .C(_3315_), .Y(_3549_) );
XOR2X1 XOR2X1_69 ( .gnd(gnd), .vdd(vdd), .A(_3548_), .B(_3549_), .Y(_3550_) );
AOI21X1 AOI21X1_555 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe64_bF_buf0), .B(_3550_), .C(micro_hash_ucr_pipe66_bF_buf2), .Y(_3551_) );
OAI21X1 OAI21X1_938 ( .gnd(gnd), .vdd(vdd), .A(_3546_), .B(micro_hash_ucr_pipe64_bF_buf4), .C(_3551_), .Y(_3552_) );
INVX2 INVX2_123 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_238_), .Y(_3553_) );
XNOR2X1 XNOR2X1_148 ( .gnd(gnd), .vdd(vdd), .A(_3351__bF_buf2), .B(_3553_), .Y(_3554_) );
OAI21X1 OAI21X1_939 ( .gnd(gnd), .vdd(vdd), .A(_3319_), .B(_3320_), .C(_3322_), .Y(_3555_) );
NOR2X1 NOR2X1_668 ( .gnd(gnd), .vdd(vdd), .A(_3555_), .B(_3554_), .Y(_3556_) );
NAND2X1 NAND2X1_446 ( .gnd(gnd), .vdd(vdd), .A(_3555_), .B(_3554_), .Y(_3557_) );
INVX1 INVX1_313 ( .gnd(gnd), .vdd(vdd), .A(_3557_), .Y(_3558_) );
OAI21X1 OAI21X1_940 ( .gnd(gnd), .vdd(vdd), .A(_3558_), .B(_3556_), .C(micro_hash_ucr_pipe66_bF_buf1), .Y(_3559_) );
NAND3X1 NAND3X1_123 ( .gnd(gnd), .vdd(vdd), .A(_878__bF_buf3), .B(_3559_), .C(_3552_), .Y(_3560_) );
INVX2 INVX2_124 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_246_), .Y(_3561_) );
XNOR2X1 XNOR2X1_149 ( .gnd(gnd), .vdd(vdd), .A(_3351__bF_buf1), .B(_3561_), .Y(_3562_) );
INVX1 INVX1_314 ( .gnd(gnd), .vdd(vdd), .A(_3332_), .Y(_3563_) );
OAI21X1 OAI21X1_941 ( .gnd(gnd), .vdd(vdd), .A(_3328_), .B(_3331_), .C(_3563_), .Y(_3564_) );
XOR2X1 XOR2X1_70 ( .gnd(gnd), .vdd(vdd), .A(_3562_), .B(_3564_), .Y(_3565_) );
AOI21X1 AOI21X1_556 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe68), .B(_3565_), .C(micro_hash_ucr_pipe69), .Y(_3566_) );
XNOR2X1 XNOR2X1_150 ( .gnd(gnd), .vdd(vdd), .A(_3351__bF_buf0), .B(micro_hash_ucr_Wx_254_), .Y(_3567_) );
AOI21X1 AOI21X1_557 ( .gnd(gnd), .vdd(vdd), .A(_3341_), .B(_3339_), .C(_3342_), .Y(_3568_) );
AND2X2 AND2X2_247 ( .gnd(gnd), .vdd(vdd), .A(_3568_), .B(_3567_), .Y(_3569_) );
NOR2X1 NOR2X1_669 ( .gnd(gnd), .vdd(vdd), .A(_400__bF_buf4), .B(_3569_), .Y(_3570_) );
OAI21X1 OAI21X1_942 ( .gnd(gnd), .vdd(vdd), .A(_3567_), .B(_3568_), .C(_3570_), .Y(_3571_) );
AOI22X1 AOI22X1_34 ( .gnd(gnd), .vdd(vdd), .A(_1950_), .B(_3571_), .C(_3560_), .D(_3566_), .Y(_299__6_) );
NAND2X1 NAND2X1_447 ( .gnd(gnd), .vdd(vdd), .A(_3537_), .B(_3536_), .Y(_3572_) );
OAI21X1 OAI21X1_943 ( .gnd(gnd), .vdd(vdd), .A(_581_), .B(_3352__bF_buf1), .C(_3572_), .Y(_3573_) );
AOI21X1 AOI21X1_558 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_k_6_), .B(micro_hash_ucr_x_6_), .C(_3350_), .Y(_3574_) );
XOR2X1 XOR2X1_71 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_k_7_), .B(micro_hash_ucr_x_7_), .Y(_3575_) );
XNOR2X1 XNOR2X1_151 ( .gnd(gnd), .vdd(vdd), .A(_3574_), .B(_3575_), .Y(_3576_) );
XNOR2X1 XNOR2X1_152 ( .gnd(gnd), .vdd(vdd), .A(_3576__bF_buf4), .B(micro_hash_ucr_Wx_215_), .Y(_3577_) );
XNOR2X1 XNOR2X1_153 ( .gnd(gnd), .vdd(vdd), .A(_3573_), .B(_3577_), .Y(_3578_) );
NAND2X1 NAND2X1_448 ( .gnd(gnd), .vdd(vdd), .A(_3504_), .B(_3505_), .Y(_3579_) );
OAI21X1 OAI21X1_944 ( .gnd(gnd), .vdd(vdd), .A(_735_), .B(_3352__bF_buf0), .C(_3579_), .Y(_3580_) );
XNOR2X1 XNOR2X1_154 ( .gnd(gnd), .vdd(vdd), .A(_3576__bF_buf3), .B(micro_hash_ucr_Wx_167_), .Y(_3581_) );
XNOR2X1 XNOR2X1_155 ( .gnd(gnd), .vdd(vdd), .A(_3580_), .B(_3581_), .Y(_3582_) );
NAND2X1 NAND2X1_449 ( .gnd(gnd), .vdd(vdd), .A(_3485_), .B(_3487_), .Y(_3583_) );
OAI21X1 OAI21X1_945 ( .gnd(gnd), .vdd(vdd), .A(_802_), .B(_3352__bF_buf4), .C(_3583_), .Y(_3584_) );
XNOR2X1 XNOR2X1_156 ( .gnd(gnd), .vdd(vdd), .A(_3576__bF_buf2), .B(micro_hash_ucr_Wx_143_), .Y(_3585_) );
XNOR2X1 XNOR2X1_157 ( .gnd(gnd), .vdd(vdd), .A(_3584_), .B(_3585_), .Y(_3586_) );
NAND2X1 NAND2X1_450 ( .gnd(gnd), .vdd(vdd), .A(_3467_), .B(_3465_), .Y(_3587_) );
OAI21X1 OAI21X1_946 ( .gnd(gnd), .vdd(vdd), .A(_524_), .B(_3352__bF_buf3), .C(_3587_), .Y(_3588_) );
XNOR2X1 XNOR2X1_158 ( .gnd(gnd), .vdd(vdd), .A(_3576__bF_buf1), .B(micro_hash_ucr_Wx_119_), .Y(_3589_) );
AND2X2 AND2X2_248 ( .gnd(gnd), .vdd(vdd), .A(_3588_), .B(_3589_), .Y(_3590_) );
OAI21X1 OAI21X1_947 ( .gnd(gnd), .vdd(vdd), .A(_801_), .B(_3352__bF_buf2), .C(_3448_), .Y(_3591_) );
XNOR2X1 XNOR2X1_159 ( .gnd(gnd), .vdd(vdd), .A(_3576__bF_buf0), .B(micro_hash_ucr_Wx_95_), .Y(_3592_) );
XNOR2X1 XNOR2X1_160 ( .gnd(gnd), .vdd(vdd), .A(_3591_), .B(_3592_), .Y(_3593_) );
OAI21X1 OAI21X1_948 ( .gnd(gnd), .vdd(vdd), .A(_3401_), .B(_3352__bF_buf1), .C(_3405_), .Y(_3594_) );
XNOR2X1 XNOR2X1_161 ( .gnd(gnd), .vdd(vdd), .A(_3576__bF_buf4), .B(micro_hash_ucr_Wx_47_), .Y(_3595_) );
XNOR2X1 XNOR2X1_162 ( .gnd(gnd), .vdd(vdd), .A(_3594_), .B(_3595_), .Y(_3596_) );
INVX1 INVX1_315 ( .gnd(gnd), .vdd(vdd), .A(_3397_), .Y(_3597_) );
OAI21X1 OAI21X1_949 ( .gnd(gnd), .vdd(vdd), .A(_3597_), .B(_3398_), .C(_3394_), .Y(_3598_) );
XNOR2X1 XNOR2X1_163 ( .gnd(gnd), .vdd(vdd), .A(_3576__bF_buf3), .B(micro_hash_ucr_Wx_39_), .Y(_3599_) );
XNOR2X1 XNOR2X1_164 ( .gnd(gnd), .vdd(vdd), .A(_3598_), .B(_3599_), .Y(_3600_) );
AOI21X1 AOI21X1_559 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_6_), .B(_3351__bF_buf4), .C(_3367_), .Y(_3601_) );
XNOR2X1 XNOR2X1_165 ( .gnd(gnd), .vdd(vdd), .A(_3576__bF_buf2), .B(micro_hash_ucr_Wx_7_), .Y(_3602_) );
XNOR2X1 XNOR2X1_166 ( .gnd(gnd), .vdd(vdd), .A(_3601_), .B(_3602_), .Y(_3603_) );
OAI21X1 OAI21X1_950 ( .gnd(gnd), .vdd(vdd), .A(_1720_), .B(micro_hash_ucr_pipe6), .C(_938_), .Y(_3604_) );
AOI21X1 AOI21X1_560 ( .gnd(gnd), .vdd(vdd), .A(H_23_), .B(micro_hash_ucr_pipe6), .C(_3604_), .Y(_3605_) );
AOI21X1 AOI21X1_561 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe8), .B(_3603_), .C(_3605_), .Y(_3606_) );
OAI21X1 OAI21X1_951 ( .gnd(gnd), .vdd(vdd), .A(_3370_), .B(_3352__bF_buf0), .C(_3377_), .Y(_3607_) );
XOR2X1 XOR2X1_72 ( .gnd(gnd), .vdd(vdd), .A(_3576__bF_buf1), .B(micro_hash_ucr_Wx_15_), .Y(_3608_) );
XNOR2X1 XNOR2X1_167 ( .gnd(gnd), .vdd(vdd), .A(_3607_), .B(_3608_), .Y(_3609_) );
NAND2X1 NAND2X1_451 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe10), .B(_3609_), .Y(_3610_) );
OAI21X1 OAI21X1_952 ( .gnd(gnd), .vdd(vdd), .A(_3606_), .B(micro_hash_ucr_pipe10), .C(_3610_), .Y(_3611_) );
NAND2X1 NAND2X1_452 ( .gnd(gnd), .vdd(vdd), .A(_3382_), .B(_3381_), .Y(_3612_) );
OAI21X1 OAI21X1_953 ( .gnd(gnd), .vdd(vdd), .A(_3380_), .B(_3352__bF_buf4), .C(_3612_), .Y(_3613_) );
XNOR2X1 XNOR2X1_168 ( .gnd(gnd), .vdd(vdd), .A(_3576__bF_buf0), .B(micro_hash_ucr_Wx_23_), .Y(_3614_) );
XOR2X1 XOR2X1_73 ( .gnd(gnd), .vdd(vdd), .A(_3613_), .B(_3614_), .Y(_3615_) );
MUX2X1 MUX2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_3611_), .B(_3615_), .S(_931_), .Y(_3616_) );
OAI21X1 OAI21X1_954 ( .gnd(gnd), .vdd(vdd), .A(_3385_), .B(_3352__bF_buf3), .C(_3391_), .Y(_3617_) );
XNOR2X1 XNOR2X1_169 ( .gnd(gnd), .vdd(vdd), .A(_3576__bF_buf4), .B(micro_hash_ucr_Wx_31_), .Y(_3618_) );
AND2X2 AND2X2_249 ( .gnd(gnd), .vdd(vdd), .A(_3617_), .B(_3618_), .Y(_3619_) );
OAI21X1 OAI21X1_955 ( .gnd(gnd), .vdd(vdd), .A(_3617_), .B(_3618_), .C(micro_hash_ucr_pipe14_bF_buf0), .Y(_3620_) );
OAI22X1 OAI22X1_57 ( .gnd(gnd), .vdd(vdd), .A(_3619_), .B(_3620_), .C(_3616_), .D(micro_hash_ucr_pipe14_bF_buf4), .Y(_3621_) );
NAND2X1 NAND2X1_453 ( .gnd(gnd), .vdd(vdd), .A(_930__bF_buf2), .B(_3621_), .Y(_3622_) );
OAI21X1 OAI21X1_956 ( .gnd(gnd), .vdd(vdd), .A(_930__bF_buf1), .B(_3600_), .C(_3622_), .Y(_3623_) );
NAND2X1 NAND2X1_454 ( .gnd(gnd), .vdd(vdd), .A(_925__bF_buf1), .B(_3623_), .Y(_3624_) );
OAI21X1 OAI21X1_957 ( .gnd(gnd), .vdd(vdd), .A(_925__bF_buf0), .B(_3596_), .C(_3624_), .Y(_3625_) );
OAI21X1 OAI21X1_958 ( .gnd(gnd), .vdd(vdd), .A(_3408_), .B(_3352__bF_buf2), .C(_3412_), .Y(_3626_) );
XNOR2X1 XNOR2X1_170 ( .gnd(gnd), .vdd(vdd), .A(_3576__bF_buf3), .B(micro_hash_ucr_Wx_55_), .Y(_3627_) );
XNOR2X1 XNOR2X1_171 ( .gnd(gnd), .vdd(vdd), .A(_3626_), .B(_3627_), .Y(_3628_) );
OAI21X1 OAI21X1_959 ( .gnd(gnd), .vdd(vdd), .A(_3628_), .B(_926__bF_buf3), .C(_924__bF_buf1), .Y(_3629_) );
AOI21X1 AOI21X1_562 ( .gnd(gnd), .vdd(vdd), .A(_926__bF_buf2), .B(_3625_), .C(_3629_), .Y(_3630_) );
AOI21X1 AOI21X1_563 ( .gnd(gnd), .vdd(vdd), .A(_3419_), .B(_3422_), .C(_3417_), .Y(_3631_) );
XNOR2X1 XNOR2X1_172 ( .gnd(gnd), .vdd(vdd), .A(_3576__bF_buf2), .B(micro_hash_ucr_Wx_63_), .Y(_3632_) );
AND2X2 AND2X2_250 ( .gnd(gnd), .vdd(vdd), .A(_3631_), .B(_3632_), .Y(_3633_) );
OAI21X1 OAI21X1_960 ( .gnd(gnd), .vdd(vdd), .A(_3631_), .B(_3632_), .C(micro_hash_ucr_pipe22_bF_buf4), .Y(_3634_) );
OAI21X1 OAI21X1_961 ( .gnd(gnd), .vdd(vdd), .A(_3633_), .B(_3634_), .C(_919__bF_buf1), .Y(_3635_) );
AOI21X1 AOI21X1_564 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_70_), .B(_3351__bF_buf3), .C(_3428_), .Y(_3636_) );
XNOR2X1 XNOR2X1_173 ( .gnd(gnd), .vdd(vdd), .A(_3576__bF_buf1), .B(_873_), .Y(_3637_) );
AOI21X1 AOI21X1_565 ( .gnd(gnd), .vdd(vdd), .A(_3637_), .B(_3636_), .C(_919__bF_buf0), .Y(_3638_) );
OAI21X1 OAI21X1_962 ( .gnd(gnd), .vdd(vdd), .A(_3636_), .B(_3637_), .C(_3638_), .Y(_3639_) );
OAI21X1 OAI21X1_963 ( .gnd(gnd), .vdd(vdd), .A(_3630_), .B(_3635_), .C(_3639_), .Y(_3640_) );
OAI21X1 OAI21X1_964 ( .gnd(gnd), .vdd(vdd), .A(_847_), .B(_3352__bF_buf1), .C(_3436_), .Y(_3641_) );
XNOR2X1 XNOR2X1_174 ( .gnd(gnd), .vdd(vdd), .A(_3576__bF_buf0), .B(_850_), .Y(_3642_) );
XNOR2X1 XNOR2X1_175 ( .gnd(gnd), .vdd(vdd), .A(_3641_), .B(_3642_), .Y(_3643_) );
MUX2X1 MUX2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_3640_), .B(_3643_), .S(_920__bF_buf0), .Y(_3644_) );
NOR2X1 NOR2X1_670 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe28_bF_buf3), .B(_3644_), .Y(_3645_) );
NAND2X1 NAND2X1_455 ( .gnd(gnd), .vdd(vdd), .A(_3440_), .B(_3442_), .Y(_3646_) );
OAI21X1 OAI21X1_965 ( .gnd(gnd), .vdd(vdd), .A(_758_), .B(_3352__bF_buf0), .C(_3646_), .Y(_3647_) );
XNOR2X1 XNOR2X1_176 ( .gnd(gnd), .vdd(vdd), .A(_3576__bF_buf4), .B(micro_hash_ucr_Wx_87_), .Y(_3648_) );
OAI21X1 OAI21X1_966 ( .gnd(gnd), .vdd(vdd), .A(_3647_), .B(_3648_), .C(micro_hash_ucr_pipe28_bF_buf2), .Y(_3649_) );
AOI21X1 AOI21X1_566 ( .gnd(gnd), .vdd(vdd), .A(_3647_), .B(_3648_), .C(_3649_), .Y(_3650_) );
OAI21X1 OAI21X1_967 ( .gnd(gnd), .vdd(vdd), .A(_3645_), .B(_3650_), .C(_913__bF_buf2), .Y(_3651_) );
OAI21X1 OAI21X1_968 ( .gnd(gnd), .vdd(vdd), .A(_913__bF_buf1), .B(_3593_), .C(_3651_), .Y(_3652_) );
OAI21X1 OAI21X1_969 ( .gnd(gnd), .vdd(vdd), .A(_663_), .B(_3352__bF_buf4), .C(_3456_), .Y(_3653_) );
XNOR2X1 XNOR2X1_177 ( .gnd(gnd), .vdd(vdd), .A(_3576__bF_buf3), .B(_667_), .Y(_3654_) );
XNOR2X1 XNOR2X1_178 ( .gnd(gnd), .vdd(vdd), .A(_3653_), .B(_3654_), .Y(_3655_) );
MUX2X1 MUX2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_3652_), .B(_3655_), .S(_914__bF_buf0), .Y(_3656_) );
NOR2X1 NOR2X1_671 ( .gnd(gnd), .vdd(vdd), .A(_3460_), .B(_3461_), .Y(_3657_) );
AOI21X1 AOI21X1_567 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_110_), .B(_3351__bF_buf2), .C(_3657_), .Y(_3658_) );
XNOR2X1 XNOR2X1_179 ( .gnd(gnd), .vdd(vdd), .A(_3576__bF_buf2), .B(_694_), .Y(_3659_) );
AOI21X1 AOI21X1_568 ( .gnd(gnd), .vdd(vdd), .A(_3659_), .B(_3658_), .C(_912__bF_buf4), .Y(_3660_) );
OAI21X1 OAI21X1_970 ( .gnd(gnd), .vdd(vdd), .A(_3658_), .B(_3659_), .C(_3660_), .Y(_3661_) );
OAI21X1 OAI21X1_971 ( .gnd(gnd), .vdd(vdd), .A(_3656_), .B(micro_hash_ucr_pipe34_bF_buf3), .C(_3661_), .Y(_3662_) );
NAND2X1 NAND2X1_456 ( .gnd(gnd), .vdd(vdd), .A(_907__bF_buf4), .B(_3662_), .Y(_3663_) );
OAI21X1 OAI21X1_972 ( .gnd(gnd), .vdd(vdd), .A(_3588_), .B(_3589_), .C(micro_hash_ucr_pipe36_bF_buf2), .Y(_3664_) );
OAI21X1 OAI21X1_973 ( .gnd(gnd), .vdd(vdd), .A(_3590_), .B(_3664_), .C(_3663_), .Y(_3665_) );
OAI21X1 OAI21X1_974 ( .gnd(gnd), .vdd(vdd), .A(_580_), .B(_3352__bF_buf3), .C(_3475_), .Y(_3666_) );
XNOR2X1 XNOR2X1_180 ( .gnd(gnd), .vdd(vdd), .A(_3576__bF_buf1), .B(_584_), .Y(_3667_) );
XNOR2X1 XNOR2X1_181 ( .gnd(gnd), .vdd(vdd), .A(_3666_), .B(_3667_), .Y(_3668_) );
MUX2X1 MUX2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_3665_), .B(_3668_), .S(_908__bF_buf0), .Y(_3669_) );
NOR2X1 NOR2X1_672 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe40_bF_buf1), .B(_3669_), .Y(_3670_) );
OAI21X1 OAI21X1_975 ( .gnd(gnd), .vdd(vdd), .A(_553_), .B(_3352__bF_buf2), .C(_3482_), .Y(_3671_) );
XNOR2X1 XNOR2X1_182 ( .gnd(gnd), .vdd(vdd), .A(_3576__bF_buf0), .B(micro_hash_ucr_Wx_135_), .Y(_3672_) );
OAI21X1 OAI21X1_976 ( .gnd(gnd), .vdd(vdd), .A(_3671_), .B(_3672_), .C(micro_hash_ucr_pipe40_bF_buf0), .Y(_3673_) );
AOI21X1 AOI21X1_569 ( .gnd(gnd), .vdd(vdd), .A(_3671_), .B(_3672_), .C(_3673_), .Y(_3674_) );
OAI21X1 OAI21X1_977 ( .gnd(gnd), .vdd(vdd), .A(_3670_), .B(_3674_), .C(_901__bF_buf1), .Y(_3675_) );
OAI21X1 OAI21X1_978 ( .gnd(gnd), .vdd(vdd), .A(_901__bF_buf0), .B(_3586_), .C(_3675_), .Y(_3676_) );
OAI21X1 OAI21X1_979 ( .gnd(gnd), .vdd(vdd), .A(_633_), .B(_3352__bF_buf1), .C(_3493_), .Y(_3677_) );
XNOR2X1 XNOR2X1_183 ( .gnd(gnd), .vdd(vdd), .A(_3576__bF_buf4), .B(_637_), .Y(_3678_) );
XNOR2X1 XNOR2X1_184 ( .gnd(gnd), .vdd(vdd), .A(_3677_), .B(_3678_), .Y(_3679_) );
MUX2X1 MUX2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_3676_), .B(_3679_), .S(_902__bF_buf1), .Y(_3680_) );
NOR2X1 NOR2X1_673 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe46_bF_buf3), .B(_3680_), .Y(_3681_) );
OAI21X1 OAI21X1_980 ( .gnd(gnd), .vdd(vdd), .A(_691_), .B(_3352__bF_buf0), .C(_3500_), .Y(_3682_) );
XNOR2X1 XNOR2X1_185 ( .gnd(gnd), .vdd(vdd), .A(_3576__bF_buf3), .B(micro_hash_ucr_Wx_159_), .Y(_3683_) );
OAI21X1 OAI21X1_981 ( .gnd(gnd), .vdd(vdd), .A(_3682_), .B(_3683_), .C(micro_hash_ucr_pipe46_bF_buf2), .Y(_3684_) );
AOI21X1 AOI21X1_570 ( .gnd(gnd), .vdd(vdd), .A(_3682_), .B(_3683_), .C(_3684_), .Y(_3685_) );
OAI21X1 OAI21X1_982 ( .gnd(gnd), .vdd(vdd), .A(_3681_), .B(_3685_), .C(_895__bF_buf2), .Y(_3686_) );
OAI21X1 OAI21X1_983 ( .gnd(gnd), .vdd(vdd), .A(_895__bF_buf1), .B(_3582_), .C(_3686_), .Y(_3687_) );
OAI21X1 OAI21X1_984 ( .gnd(gnd), .vdd(vdd), .A(_714_), .B(_3352__bF_buf4), .C(_3511_), .Y(_3688_) );
XOR2X1 XOR2X1_74 ( .gnd(gnd), .vdd(vdd), .A(_3576__bF_buf2), .B(micro_hash_ucr_Wx_175_), .Y(_3689_) );
XNOR2X1 XNOR2X1_186 ( .gnd(gnd), .vdd(vdd), .A(_3688_), .B(_3689_), .Y(_3690_) );
MUX2X1 MUX2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_3687_), .B(_3690_), .S(_896__bF_buf3), .Y(_3691_) );
AOI21X1 AOI21X1_571 ( .gnd(gnd), .vdd(vdd), .A(_3355_), .B(_3358_), .C(_3353_), .Y(_3692_) );
XNOR2X1 XNOR2X1_187 ( .gnd(gnd), .vdd(vdd), .A(_3576__bF_buf1), .B(_608_), .Y(_3693_) );
AOI21X1 AOI21X1_572 ( .gnd(gnd), .vdd(vdd), .A(_3692_), .B(_3693_), .C(_894__bF_buf0), .Y(_3694_) );
OAI21X1 OAI21X1_985 ( .gnd(gnd), .vdd(vdd), .A(_3692_), .B(_3693_), .C(_3694_), .Y(_3695_) );
OAI21X1 OAI21X1_986 ( .gnd(gnd), .vdd(vdd), .A(_3691_), .B(micro_hash_ucr_pipe52_bF_buf2), .C(_3695_), .Y(_3696_) );
OAI21X1 OAI21X1_987 ( .gnd(gnd), .vdd(vdd), .A(_664_), .B(_3352__bF_buf3), .C(_3519_), .Y(_3697_) );
XNOR2X1 XNOR2X1_188 ( .gnd(gnd), .vdd(vdd), .A(_3576__bF_buf0), .B(micro_hash_ucr_Wx_191_), .Y(_3698_) );
OAI21X1 OAI21X1_988 ( .gnd(gnd), .vdd(vdd), .A(_3697_), .B(_3698_), .C(micro_hash_ucr_pipe54_bF_buf1), .Y(_3699_) );
AOI21X1 AOI21X1_573 ( .gnd(gnd), .vdd(vdd), .A(_3697_), .B(_3698_), .C(_3699_), .Y(_3700_) );
AOI21X1 AOI21X1_574 ( .gnd(gnd), .vdd(vdd), .A(_889__bF_buf0), .B(_3696_), .C(_3700_), .Y(_3701_) );
AOI21X1 AOI21X1_575 ( .gnd(gnd), .vdd(vdd), .A(_3526_), .B(_3528_), .C(_3524_), .Y(_3702_) );
XNOR2X1 XNOR2X1_189 ( .gnd(gnd), .vdd(vdd), .A(_3576__bF_buf4), .B(micro_hash_ucr_Wx_199_), .Y(_3703_) );
AND2X2 AND2X2_251 ( .gnd(gnd), .vdd(vdd), .A(_3703_), .B(_3702_), .Y(_3704_) );
OAI21X1 OAI21X1_989 ( .gnd(gnd), .vdd(vdd), .A(_3703_), .B(_3702_), .C(micro_hash_ucr_pipe56_bF_buf1), .Y(_3705_) );
OAI21X1 OAI21X1_990 ( .gnd(gnd), .vdd(vdd), .A(_3704_), .B(_3705_), .C(_888__bF_buf0), .Y(_3706_) );
AOI21X1 AOI21X1_576 ( .gnd(gnd), .vdd(vdd), .A(_890__bF_buf1), .B(_3701_), .C(_3706_), .Y(_3707_) );
NAND2X1 NAND2X1_457 ( .gnd(gnd), .vdd(vdd), .A(_3531_), .B(_3532_), .Y(_3708_) );
OAI21X1 OAI21X1_991 ( .gnd(gnd), .vdd(vdd), .A(_525_), .B(_3352__bF_buf2), .C(_3708_), .Y(_3709_) );
XNOR2X1 XNOR2X1_190 ( .gnd(gnd), .vdd(vdd), .A(_3576__bF_buf3), .B(micro_hash_ucr_Wx_207_), .Y(_3710_) );
OAI21X1 OAI21X1_992 ( .gnd(gnd), .vdd(vdd), .A(_3709_), .B(_3710_), .C(micro_hash_ucr_pipe58_bF_buf3), .Y(_3711_) );
AOI21X1 AOI21X1_577 ( .gnd(gnd), .vdd(vdd), .A(_3709_), .B(_3710_), .C(_3711_), .Y(_3712_) );
OAI21X1 OAI21X1_993 ( .gnd(gnd), .vdd(vdd), .A(_3707_), .B(_3712_), .C(_883__bF_buf3), .Y(_3713_) );
OAI21X1 OAI21X1_994 ( .gnd(gnd), .vdd(vdd), .A(_883__bF_buf2), .B(_3578_), .C(_3713_), .Y(_3714_) );
OAI21X1 OAI21X1_995 ( .gnd(gnd), .vdd(vdd), .A(_554_), .B(_3352__bF_buf1), .C(_3543_), .Y(_3715_) );
XNOR2X1 XNOR2X1_191 ( .gnd(gnd), .vdd(vdd), .A(_3576__bF_buf2), .B(micro_hash_ucr_Wx_223_), .Y(_3716_) );
OAI21X1 OAI21X1_996 ( .gnd(gnd), .vdd(vdd), .A(_3715_), .B(_3716_), .C(micro_hash_ucr_pipe62_bF_buf3), .Y(_3717_) );
AOI21X1 AOI21X1_578 ( .gnd(gnd), .vdd(vdd), .A(_3715_), .B(_3716_), .C(_3717_), .Y(_3718_) );
AOI21X1 AOI21X1_579 ( .gnd(gnd), .vdd(vdd), .A(_884__bF_buf3), .B(_3714_), .C(_3718_), .Y(_3719_) );
NAND2X1 NAND2X1_458 ( .gnd(gnd), .vdd(vdd), .A(_3549_), .B(_3548_), .Y(_3720_) );
OAI21X1 OAI21X1_997 ( .gnd(gnd), .vdd(vdd), .A(_3547_), .B(_3352__bF_buf0), .C(_3720_), .Y(_3721_) );
XOR2X1 XOR2X1_75 ( .gnd(gnd), .vdd(vdd), .A(_3576__bF_buf1), .B(micro_hash_ucr_Wx_231_), .Y(_3722_) );
NOR2X1 NOR2X1_674 ( .gnd(gnd), .vdd(vdd), .A(_3722_), .B(_3721_), .Y(_3723_) );
AND2X2 AND2X2_252 ( .gnd(gnd), .vdd(vdd), .A(_3721_), .B(_3722_), .Y(_3724_) );
OAI21X1 OAI21X1_998 ( .gnd(gnd), .vdd(vdd), .A(_3723_), .B(_3724_), .C(micro_hash_ucr_pipe64_bF_buf3), .Y(_3725_) );
OAI21X1 OAI21X1_999 ( .gnd(gnd), .vdd(vdd), .A(_3719_), .B(micro_hash_ucr_pipe64_bF_buf2), .C(_3725_), .Y(_3726_) );
OAI21X1 OAI21X1_1000 ( .gnd(gnd), .vdd(vdd), .A(_3553_), .B(_3352__bF_buf4), .C(_3557_), .Y(_3727_) );
XNOR2X1 XNOR2X1_192 ( .gnd(gnd), .vdd(vdd), .A(_3576__bF_buf0), .B(micro_hash_ucr_Wx_239_), .Y(_3728_) );
OAI21X1 OAI21X1_1001 ( .gnd(gnd), .vdd(vdd), .A(_3727_), .B(_3728_), .C(micro_hash_ucr_pipe66_bF_buf0), .Y(_3729_) );
AOI21X1 AOI21X1_580 ( .gnd(gnd), .vdd(vdd), .A(_3727_), .B(_3728_), .C(_3729_), .Y(_3730_) );
AOI21X1 AOI21X1_581 ( .gnd(gnd), .vdd(vdd), .A(_877__bF_buf2), .B(_3726_), .C(_3730_), .Y(_3731_) );
NAND2X1 NAND2X1_459 ( .gnd(gnd), .vdd(vdd), .A(_3564_), .B(_3562_), .Y(_3732_) );
OAI21X1 OAI21X1_1002 ( .gnd(gnd), .vdd(vdd), .A(_3561_), .B(_3352__bF_buf3), .C(_3732_), .Y(_3733_) );
XNOR2X1 XNOR2X1_193 ( .gnd(gnd), .vdd(vdd), .A(_3576__bF_buf4), .B(micro_hash_ucr_Wx_247_), .Y(_3734_) );
XOR2X1 XOR2X1_76 ( .gnd(gnd), .vdd(vdd), .A(_3733_), .B(_3734_), .Y(_3735_) );
OAI21X1 OAI21X1_1003 ( .gnd(gnd), .vdd(vdd), .A(_3735_), .B(_878__bF_buf2), .C(_876__bF_buf2), .Y(_3736_) );
AOI21X1 AOI21X1_582 ( .gnd(gnd), .vdd(vdd), .A(_878__bF_buf1), .B(_3731_), .C(_3736_), .Y(_3737_) );
NAND2X1 NAND2X1_460 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_254_), .B(_3351__bF_buf1), .Y(_3738_) );
OAI21X1 OAI21X1_1004 ( .gnd(gnd), .vdd(vdd), .A(_3568_), .B(_3567_), .C(_3738_), .Y(_3739_) );
XNOR2X1 XNOR2X1_194 ( .gnd(gnd), .vdd(vdd), .A(_3576__bF_buf3), .B(micro_hash_ucr_Wx_255_), .Y(_3740_) );
AND2X2 AND2X2_253 ( .gnd(gnd), .vdd(vdd), .A(_3739_), .B(_3740_), .Y(_3741_) );
OAI21X1 OAI21X1_1005 ( .gnd(gnd), .vdd(vdd), .A(_3739_), .B(_3740_), .C(micro_hash_ucr_pipe69), .Y(_3742_) );
OAI21X1 OAI21X1_1006 ( .gnd(gnd), .vdd(vdd), .A(_3741_), .B(_3742_), .C(_302__bF_buf0), .Y(_3743_) );
NOR2X1 NOR2X1_675 ( .gnd(gnd), .vdd(vdd), .A(_3743_), .B(_3737_), .Y(_299__7_) );
NOR2X1 NOR2X1_676 ( .gnd(gnd), .vdd(vdd), .A(_1403_), .B(_956_), .Y(_3744_) );
OAI21X1 OAI21X1_1007 ( .gnd(gnd), .vdd(vdd), .A(_1849_), .B(_4478_), .C(_947_), .Y(_3745_) );
NOR2X1 NOR2X1_677 ( .gnd(gnd), .vdd(vdd), .A(_3745_), .B(_3744_), .Y(_3746_) );
NAND2X1 NAND2X1_461 ( .gnd(gnd), .vdd(vdd), .A(_936_), .B(_1073_), .Y(_3747_) );
NOR2X1 NOR2X1_678 ( .gnd(gnd), .vdd(vdd), .A(_1295_), .B(_3747_), .Y(_3748_) );
OAI21X1 OAI21X1_1008 ( .gnd(gnd), .vdd(vdd), .A(_3748_), .B(micro_hash_ucr_b_0_bF_buf3_), .C(_928_), .Y(_3749_) );
OAI21X1 OAI21X1_1009 ( .gnd(gnd), .vdd(vdd), .A(_3746_), .B(_3749_), .C(_930__bF_buf0), .Y(_3750_) );
AOI21X1 AOI21X1_583 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe16_bF_buf1), .B(_4481_), .C(micro_hash_ucr_pipe17_bF_buf3), .Y(_3751_) );
AOI21X1 AOI21X1_584 ( .gnd(gnd), .vdd(vdd), .A(_3751_), .B(_3750_), .C(micro_hash_ucr_pipe18_bF_buf4), .Y(_3752_) );
OAI21X1 OAI21X1_1010 ( .gnd(gnd), .vdd(vdd), .A(_925__bF_buf4), .B(micro_hash_ucr_b_0_bF_buf2_), .C(_927__bF_buf1), .Y(_3753_) );
OAI21X1 OAI21X1_1011 ( .gnd(gnd), .vdd(vdd), .A(_3752_), .B(_3753_), .C(_926__bF_buf1), .Y(_3754_) );
AOI21X1 AOI21X1_585 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe20_bF_buf2), .B(_4481_), .C(micro_hash_ucr_pipe21_bF_buf1), .Y(_3755_) );
AOI21X1 AOI21X1_586 ( .gnd(gnd), .vdd(vdd), .A(_3755_), .B(_3754_), .C(micro_hash_ucr_pipe22_bF_buf3), .Y(_3756_) );
OAI21X1 OAI21X1_1012 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf0), .B(micro_hash_ucr_b_0_bF_buf1_), .C(_923_), .Y(_3757_) );
OAI21X1 OAI21X1_1013 ( .gnd(gnd), .vdd(vdd), .A(_3756_), .B(_3757_), .C(_919__bF_buf4), .Y(_3758_) );
AOI21X1 AOI21X1_587 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe24_bF_buf4), .B(_4481_), .C(micro_hash_ucr_pipe25), .Y(_3759_) );
AOI21X1 AOI21X1_588 ( .gnd(gnd), .vdd(vdd), .A(_3759_), .B(_3758_), .C(micro_hash_ucr_pipe26_bF_buf2), .Y(_3760_) );
OAI21X1 OAI21X1_1014 ( .gnd(gnd), .vdd(vdd), .A(_920__bF_buf4), .B(micro_hash_ucr_b_0_bF_buf0_), .C(_916_), .Y(_3761_) );
OAI21X1 OAI21X1_1015 ( .gnd(gnd), .vdd(vdd), .A(_3760_), .B(_3761_), .C(_918__bF_buf4), .Y(_3762_) );
AOI21X1 AOI21X1_589 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe28_bF_buf1), .B(_4481_), .C(micro_hash_ucr_pipe29_bF_buf3), .Y(_3763_) );
AOI21X1 AOI21X1_590 ( .gnd(gnd), .vdd(vdd), .A(_3763_), .B(_3762_), .C(micro_hash_ucr_pipe30_bF_buf0), .Y(_3764_) );
OAI21X1 OAI21X1_1016 ( .gnd(gnd), .vdd(vdd), .A(_913__bF_buf0), .B(micro_hash_ucr_b_0_bF_buf3_), .C(_915__bF_buf2), .Y(_3765_) );
OAI21X1 OAI21X1_1017 ( .gnd(gnd), .vdd(vdd), .A(_3764_), .B(_3765_), .C(_914__bF_buf4), .Y(_3766_) );
AOI21X1 AOI21X1_591 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe32_bF_buf3), .B(_4481_), .C(micro_hash_ucr_pipe33_bF_buf0), .Y(_3767_) );
AOI21X1 AOI21X1_592 ( .gnd(gnd), .vdd(vdd), .A(_3767_), .B(_3766_), .C(micro_hash_ucr_pipe34_bF_buf2), .Y(_3768_) );
OAI21X1 OAI21X1_1018 ( .gnd(gnd), .vdd(vdd), .A(_912__bF_buf3), .B(micro_hash_ucr_b_0_bF_buf2_), .C(_911__bF_buf3), .Y(_3769_) );
OAI21X1 OAI21X1_1019 ( .gnd(gnd), .vdd(vdd), .A(_3768_), .B(_3769_), .C(_907__bF_buf3), .Y(_3770_) );
AOI21X1 AOI21X1_593 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe36_bF_buf1), .B(_4481_), .C(micro_hash_ucr_pipe37), .Y(_3771_) );
AOI21X1 AOI21X1_594 ( .gnd(gnd), .vdd(vdd), .A(_3771_), .B(_3770_), .C(micro_hash_ucr_pipe38_bF_buf2), .Y(_3772_) );
OAI21X1 OAI21X1_1020 ( .gnd(gnd), .vdd(vdd), .A(_908__bF_buf4), .B(micro_hash_ucr_b_0_bF_buf1_), .C(_904__bF_buf3), .Y(_3773_) );
OAI21X1 OAI21X1_1021 ( .gnd(gnd), .vdd(vdd), .A(_3772_), .B(_3773_), .C(_906__bF_buf1), .Y(_3774_) );
AOI21X1 AOI21X1_595 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe40_bF_buf4), .B(_4481_), .C(micro_hash_ucr_pipe41), .Y(_3775_) );
AOI21X1 AOI21X1_596 ( .gnd(gnd), .vdd(vdd), .A(_3775_), .B(_3774_), .C(micro_hash_ucr_pipe42_bF_buf1), .Y(_3776_) );
OAI21X1 OAI21X1_1022 ( .gnd(gnd), .vdd(vdd), .A(_901__bF_buf4), .B(micro_hash_ucr_b_0_bF_buf0_), .C(_903__bF_buf2), .Y(_3777_) );
OAI21X1 OAI21X1_1023 ( .gnd(gnd), .vdd(vdd), .A(_3776_), .B(_3777_), .C(_902__bF_buf0), .Y(_3778_) );
AOI21X1 AOI21X1_597 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe44), .B(_4481_), .C(micro_hash_ucr_pipe45_bF_buf1), .Y(_3779_) );
AOI21X1 AOI21X1_598 ( .gnd(gnd), .vdd(vdd), .A(_3779_), .B(_3778_), .C(micro_hash_ucr_pipe46_bF_buf1), .Y(_3780_) );
OAI21X1 OAI21X1_1024 ( .gnd(gnd), .vdd(vdd), .A(_900__bF_buf3), .B(micro_hash_ucr_b_0_bF_buf3_), .C(_899__bF_buf1), .Y(_3781_) );
OAI21X1 OAI21X1_1025 ( .gnd(gnd), .vdd(vdd), .A(_3780_), .B(_3781_), .C(_895__bF_buf0), .Y(_3782_) );
AOI21X1 AOI21X1_599 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe48_bF_buf0), .B(_4481_), .C(micro_hash_ucr_pipe49), .Y(_3783_) );
AOI21X1 AOI21X1_600 ( .gnd(gnd), .vdd(vdd), .A(_3783_), .B(_3782_), .C(micro_hash_ucr_pipe50_bF_buf3), .Y(_3784_) );
OAI21X1 OAI21X1_1026 ( .gnd(gnd), .vdd(vdd), .A(_896__bF_buf2), .B(micro_hash_ucr_b_0_bF_buf2_), .C(_892_), .Y(_3785_) );
OAI21X1 OAI21X1_1027 ( .gnd(gnd), .vdd(vdd), .A(_3784_), .B(_3785_), .C(_894__bF_buf3), .Y(_3786_) );
AOI21X1 AOI21X1_601 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe52_bF_buf1), .B(_4481_), .C(micro_hash_ucr_pipe53_bF_buf1), .Y(_3787_) );
AOI21X1 AOI21X1_602 ( .gnd(gnd), .vdd(vdd), .A(_3787_), .B(_3786_), .C(micro_hash_ucr_pipe54_bF_buf0), .Y(_3788_) );
OAI21X1 OAI21X1_1028 ( .gnd(gnd), .vdd(vdd), .A(_889__bF_buf4), .B(micro_hash_ucr_b_0_bF_buf1_), .C(_891_), .Y(_3789_) );
OAI21X1 OAI21X1_1029 ( .gnd(gnd), .vdd(vdd), .A(_3788_), .B(_3789_), .C(_890__bF_buf0), .Y(_3790_) );
AOI21X1 AOI21X1_603 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe56_bF_buf0), .B(_4481_), .C(micro_hash_ucr_pipe57_bF_buf3), .Y(_3791_) );
AOI21X1 AOI21X1_604 ( .gnd(gnd), .vdd(vdd), .A(_3791_), .B(_3790_), .C(micro_hash_ucr_pipe58_bF_buf2), .Y(_3792_) );
OAI21X1 OAI21X1_1030 ( .gnd(gnd), .vdd(vdd), .A(_888__bF_buf3), .B(micro_hash_ucr_b_0_bF_buf0_), .C(_887__bF_buf1), .Y(_3793_) );
OAI21X1 OAI21X1_1031 ( .gnd(gnd), .vdd(vdd), .A(_3792_), .B(_3793_), .C(_883__bF_buf1), .Y(_3794_) );
AOI21X1 AOI21X1_605 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe60_bF_buf0), .B(_4481_), .C(micro_hash_ucr_pipe61_bF_buf1), .Y(_3795_) );
AOI21X1 AOI21X1_606 ( .gnd(gnd), .vdd(vdd), .A(_3795_), .B(_3794_), .C(micro_hash_ucr_pipe62_bF_buf2), .Y(_3796_) );
OAI21X1 OAI21X1_1032 ( .gnd(gnd), .vdd(vdd), .A(_884__bF_buf2), .B(micro_hash_ucr_b_0_bF_buf3_), .C(_880__bF_buf0), .Y(_3797_) );
OAI21X1 OAI21X1_1033 ( .gnd(gnd), .vdd(vdd), .A(_3796_), .B(_3797_), .C(_882__bF_buf0), .Y(_3798_) );
AOI21X1 AOI21X1_607 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe64_bF_buf1), .B(_4481_), .C(micro_hash_ucr_pipe65_bF_buf3), .Y(_3799_) );
AOI21X1 AOI21X1_608 ( .gnd(gnd), .vdd(vdd), .A(_3799_), .B(_3798_), .C(micro_hash_ucr_pipe66_bF_buf4), .Y(_3800_) );
OAI21X1 OAI21X1_1034 ( .gnd(gnd), .vdd(vdd), .A(_877__bF_buf1), .B(micro_hash_ucr_b_0_bF_buf2_), .C(_879__bF_buf0), .Y(_3801_) );
OAI21X1 OAI21X1_1035 ( .gnd(gnd), .vdd(vdd), .A(_3800_), .B(_3801_), .C(_878__bF_buf0), .Y(_3802_) );
OAI21X1 OAI21X1_1036 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_0_bF_buf1_), .B(_878__bF_buf4), .C(_3802_), .Y(_3803_) );
NOR2X1 NOR2X1_679 ( .gnd(gnd), .vdd(vdd), .A(_1950_), .B(_3803_), .Y(_298__0_) );
OAI21X1 OAI21X1_1037 ( .gnd(gnd), .vdd(vdd), .A(_1849_), .B(_4485_), .C(_947_), .Y(_3804_) );
NOR2X1 NOR2X1_680 ( .gnd(gnd), .vdd(vdd), .A(_3804_), .B(_3744_), .Y(_3805_) );
OAI21X1 OAI21X1_1038 ( .gnd(gnd), .vdd(vdd), .A(_3748_), .B(micro_hash_ucr_b_1_bF_buf3_), .C(_928_), .Y(_3806_) );
OAI21X1 OAI21X1_1039 ( .gnd(gnd), .vdd(vdd), .A(_3805_), .B(_3806_), .C(_930__bF_buf4), .Y(_3807_) );
AOI21X1 AOI21X1_609 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe16_bF_buf0), .B(_4487_), .C(micro_hash_ucr_pipe17_bF_buf2), .Y(_3808_) );
AOI21X1 AOI21X1_610 ( .gnd(gnd), .vdd(vdd), .A(_3808_), .B(_3807_), .C(micro_hash_ucr_pipe18_bF_buf3), .Y(_3809_) );
OAI21X1 OAI21X1_1040 ( .gnd(gnd), .vdd(vdd), .A(_925__bF_buf3), .B(micro_hash_ucr_b_1_bF_buf2_), .C(_927__bF_buf0), .Y(_3810_) );
OAI21X1 OAI21X1_1041 ( .gnd(gnd), .vdd(vdd), .A(_3809_), .B(_3810_), .C(_926__bF_buf0), .Y(_3811_) );
AOI21X1 AOI21X1_611 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe20_bF_buf1), .B(_4487_), .C(micro_hash_ucr_pipe21_bF_buf0), .Y(_3812_) );
AOI21X1 AOI21X1_612 ( .gnd(gnd), .vdd(vdd), .A(_3812_), .B(_3811_), .C(micro_hash_ucr_pipe22_bF_buf2), .Y(_3813_) );
OAI21X1 OAI21X1_1042 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf4), .B(micro_hash_ucr_b_1_bF_buf1_), .C(_923_), .Y(_3814_) );
OAI21X1 OAI21X1_1043 ( .gnd(gnd), .vdd(vdd), .A(_3813_), .B(_3814_), .C(_919__bF_buf3), .Y(_3815_) );
AOI21X1 AOI21X1_613 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe24_bF_buf3), .B(_4487_), .C(micro_hash_ucr_pipe25), .Y(_3816_) );
AOI21X1 AOI21X1_614 ( .gnd(gnd), .vdd(vdd), .A(_3816_), .B(_3815_), .C(micro_hash_ucr_pipe26_bF_buf1), .Y(_3817_) );
OAI21X1 OAI21X1_1044 ( .gnd(gnd), .vdd(vdd), .A(_920__bF_buf3), .B(micro_hash_ucr_b_1_bF_buf0_), .C(_916_), .Y(_3818_) );
OAI21X1 OAI21X1_1045 ( .gnd(gnd), .vdd(vdd), .A(_3817_), .B(_3818_), .C(_918__bF_buf3), .Y(_3819_) );
AOI21X1 AOI21X1_615 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe28_bF_buf0), .B(_4487_), .C(micro_hash_ucr_pipe29_bF_buf2), .Y(_3820_) );
AOI21X1 AOI21X1_616 ( .gnd(gnd), .vdd(vdd), .A(_3820_), .B(_3819_), .C(micro_hash_ucr_pipe30_bF_buf3), .Y(_3821_) );
OAI21X1 OAI21X1_1046 ( .gnd(gnd), .vdd(vdd), .A(_913__bF_buf4), .B(micro_hash_ucr_b_1_bF_buf3_), .C(_915__bF_buf1), .Y(_3822_) );
OAI21X1 OAI21X1_1047 ( .gnd(gnd), .vdd(vdd), .A(_3821_), .B(_3822_), .C(_914__bF_buf3), .Y(_3823_) );
AOI21X1 AOI21X1_617 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe32_bF_buf2), .B(_4487_), .C(micro_hash_ucr_pipe33_bF_buf3), .Y(_3824_) );
AOI21X1 AOI21X1_618 ( .gnd(gnd), .vdd(vdd), .A(_3824_), .B(_3823_), .C(micro_hash_ucr_pipe34_bF_buf1), .Y(_3825_) );
OAI21X1 OAI21X1_1048 ( .gnd(gnd), .vdd(vdd), .A(_912__bF_buf2), .B(micro_hash_ucr_b_1_bF_buf2_), .C(_911__bF_buf2), .Y(_3826_) );
OAI21X1 OAI21X1_1049 ( .gnd(gnd), .vdd(vdd), .A(_3825_), .B(_3826_), .C(_907__bF_buf2), .Y(_3827_) );
AOI21X1 AOI21X1_619 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe36_bF_buf0), .B(_4487_), .C(micro_hash_ucr_pipe37), .Y(_3828_) );
AOI21X1 AOI21X1_620 ( .gnd(gnd), .vdd(vdd), .A(_3828_), .B(_3827_), .C(micro_hash_ucr_pipe38_bF_buf1), .Y(_3829_) );
OAI21X1 OAI21X1_1050 ( .gnd(gnd), .vdd(vdd), .A(_908__bF_buf3), .B(micro_hash_ucr_b_1_bF_buf1_), .C(_904__bF_buf2), .Y(_3830_) );
OAI21X1 OAI21X1_1051 ( .gnd(gnd), .vdd(vdd), .A(_3829_), .B(_3830_), .C(_906__bF_buf0), .Y(_3831_) );
AOI21X1 AOI21X1_621 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe40_bF_buf3), .B(_4487_), .C(micro_hash_ucr_pipe41), .Y(_3832_) );
AOI21X1 AOI21X1_622 ( .gnd(gnd), .vdd(vdd), .A(_3832_), .B(_3831_), .C(micro_hash_ucr_pipe42_bF_buf0), .Y(_3833_) );
OAI21X1 OAI21X1_1052 ( .gnd(gnd), .vdd(vdd), .A(_901__bF_buf3), .B(micro_hash_ucr_b_1_bF_buf0_), .C(_903__bF_buf1), .Y(_3834_) );
OAI21X1 OAI21X1_1053 ( .gnd(gnd), .vdd(vdd), .A(_3833_), .B(_3834_), .C(_902__bF_buf4), .Y(_3835_) );
AOI21X1 AOI21X1_623 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe44), .B(_4487_), .C(micro_hash_ucr_pipe45_bF_buf0), .Y(_3836_) );
AOI21X1 AOI21X1_624 ( .gnd(gnd), .vdd(vdd), .A(_3836_), .B(_3835_), .C(micro_hash_ucr_pipe46_bF_buf0), .Y(_3837_) );
OAI21X1 OAI21X1_1054 ( .gnd(gnd), .vdd(vdd), .A(_900__bF_buf2), .B(micro_hash_ucr_b_1_bF_buf3_), .C(_899__bF_buf0), .Y(_3838_) );
OAI21X1 OAI21X1_1055 ( .gnd(gnd), .vdd(vdd), .A(_3837_), .B(_3838_), .C(_895__bF_buf4), .Y(_3839_) );
AOI21X1 AOI21X1_625 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe48_bF_buf3), .B(_4487_), .C(micro_hash_ucr_pipe49), .Y(_3840_) );
AOI21X1 AOI21X1_626 ( .gnd(gnd), .vdd(vdd), .A(_3840_), .B(_3839_), .C(micro_hash_ucr_pipe50_bF_buf2), .Y(_3841_) );
OAI21X1 OAI21X1_1056 ( .gnd(gnd), .vdd(vdd), .A(_896__bF_buf1), .B(micro_hash_ucr_b_1_bF_buf2_), .C(_892_), .Y(_3842_) );
OAI21X1 OAI21X1_1057 ( .gnd(gnd), .vdd(vdd), .A(_3841_), .B(_3842_), .C(_894__bF_buf2), .Y(_3843_) );
AOI21X1 AOI21X1_627 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe52_bF_buf0), .B(_4487_), .C(micro_hash_ucr_pipe53_bF_buf0), .Y(_3844_) );
AOI21X1 AOI21X1_628 ( .gnd(gnd), .vdd(vdd), .A(_3844_), .B(_3843_), .C(micro_hash_ucr_pipe54_bF_buf3), .Y(_3845_) );
OAI21X1 OAI21X1_1058 ( .gnd(gnd), .vdd(vdd), .A(_889__bF_buf3), .B(micro_hash_ucr_b_1_bF_buf1_), .C(_891_), .Y(_3846_) );
OAI21X1 OAI21X1_1059 ( .gnd(gnd), .vdd(vdd), .A(_3845_), .B(_3846_), .C(_890__bF_buf4), .Y(_3847_) );
AOI21X1 AOI21X1_629 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe56_bF_buf3), .B(_4487_), .C(micro_hash_ucr_pipe57_bF_buf2), .Y(_3848_) );
AOI21X1 AOI21X1_630 ( .gnd(gnd), .vdd(vdd), .A(_3848_), .B(_3847_), .C(micro_hash_ucr_pipe58_bF_buf1), .Y(_3849_) );
OAI21X1 OAI21X1_1060 ( .gnd(gnd), .vdd(vdd), .A(_888__bF_buf2), .B(micro_hash_ucr_b_1_bF_buf0_), .C(_887__bF_buf0), .Y(_3850_) );
OAI21X1 OAI21X1_1061 ( .gnd(gnd), .vdd(vdd), .A(_3849_), .B(_3850_), .C(_883__bF_buf0), .Y(_3851_) );
AOI21X1 AOI21X1_631 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe60_bF_buf4), .B(_4487_), .C(micro_hash_ucr_pipe61_bF_buf0), .Y(_3852_) );
AOI21X1 AOI21X1_632 ( .gnd(gnd), .vdd(vdd), .A(_3852_), .B(_3851_), .C(micro_hash_ucr_pipe62_bF_buf1), .Y(_3853_) );
OAI21X1 OAI21X1_1062 ( .gnd(gnd), .vdd(vdd), .A(_884__bF_buf1), .B(micro_hash_ucr_b_1_bF_buf3_), .C(_880__bF_buf3), .Y(_3854_) );
OAI21X1 OAI21X1_1063 ( .gnd(gnd), .vdd(vdd), .A(_3853_), .B(_3854_), .C(_882__bF_buf3), .Y(_3855_) );
AOI21X1 AOI21X1_633 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe64_bF_buf0), .B(_4487_), .C(micro_hash_ucr_pipe65_bF_buf2), .Y(_3856_) );
AOI21X1 AOI21X1_634 ( .gnd(gnd), .vdd(vdd), .A(_3856_), .B(_3855_), .C(micro_hash_ucr_pipe66_bF_buf3), .Y(_3857_) );
OAI21X1 OAI21X1_1064 ( .gnd(gnd), .vdd(vdd), .A(_877__bF_buf0), .B(micro_hash_ucr_b_1_bF_buf2_), .C(_879__bF_buf3), .Y(_3858_) );
OAI21X1 OAI21X1_1065 ( .gnd(gnd), .vdd(vdd), .A(_3857_), .B(_3858_), .C(_878__bF_buf3), .Y(_3859_) );
OAI21X1 OAI21X1_1066 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_1_bF_buf1_), .B(_878__bF_buf2), .C(_3859_), .Y(_3860_) );
NOR2X1 NOR2X1_681 ( .gnd(gnd), .vdd(vdd), .A(_1950_), .B(_3860_), .Y(_298__1_) );
OAI21X1 OAI21X1_1067 ( .gnd(gnd), .vdd(vdd), .A(_1849_), .B(_379_), .C(_947_), .Y(_3861_) );
NOR2X1 NOR2X1_682 ( .gnd(gnd), .vdd(vdd), .A(_3861_), .B(_3744_), .Y(_3862_) );
OAI21X1 OAI21X1_1068 ( .gnd(gnd), .vdd(vdd), .A(_3748_), .B(micro_hash_ucr_b_2_bF_buf2_), .C(_928_), .Y(_3863_) );
OAI21X1 OAI21X1_1069 ( .gnd(gnd), .vdd(vdd), .A(_3862_), .B(_3863_), .C(_930__bF_buf3), .Y(_3864_) );
AOI21X1 AOI21X1_635 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe16_bF_buf3), .B(_389_), .C(micro_hash_ucr_pipe17_bF_buf1), .Y(_3865_) );
AOI21X1 AOI21X1_636 ( .gnd(gnd), .vdd(vdd), .A(_3865_), .B(_3864_), .C(micro_hash_ucr_pipe18_bF_buf2), .Y(_3866_) );
OAI21X1 OAI21X1_1070 ( .gnd(gnd), .vdd(vdd), .A(_925__bF_buf2), .B(micro_hash_ucr_b_2_bF_buf1_), .C(_927__bF_buf3), .Y(_3867_) );
OAI21X1 OAI21X1_1071 ( .gnd(gnd), .vdd(vdd), .A(_3866_), .B(_3867_), .C(_926__bF_buf4), .Y(_3868_) );
AOI21X1 AOI21X1_637 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe20_bF_buf0), .B(_389_), .C(micro_hash_ucr_pipe21_bF_buf3), .Y(_3869_) );
AOI21X1 AOI21X1_638 ( .gnd(gnd), .vdd(vdd), .A(_3869_), .B(_3868_), .C(micro_hash_ucr_pipe22_bF_buf1), .Y(_3870_) );
OAI21X1 OAI21X1_1072 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf3), .B(micro_hash_ucr_b_2_bF_buf0_), .C(_923_), .Y(_3871_) );
OAI21X1 OAI21X1_1073 ( .gnd(gnd), .vdd(vdd), .A(_3870_), .B(_3871_), .C(_919__bF_buf2), .Y(_3872_) );
AOI21X1 AOI21X1_639 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe24_bF_buf2), .B(_389_), .C(micro_hash_ucr_pipe25), .Y(_3873_) );
AOI21X1 AOI21X1_640 ( .gnd(gnd), .vdd(vdd), .A(_3873_), .B(_3872_), .C(micro_hash_ucr_pipe26_bF_buf0), .Y(_3874_) );
OAI21X1 OAI21X1_1074 ( .gnd(gnd), .vdd(vdd), .A(_920__bF_buf2), .B(micro_hash_ucr_b_2_bF_buf3_), .C(_916_), .Y(_3875_) );
OAI21X1 OAI21X1_1075 ( .gnd(gnd), .vdd(vdd), .A(_3874_), .B(_3875_), .C(_918__bF_buf2), .Y(_3876_) );
AOI21X1 AOI21X1_641 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe28_bF_buf3), .B(_389_), .C(micro_hash_ucr_pipe29_bF_buf1), .Y(_3877_) );
AOI21X1 AOI21X1_642 ( .gnd(gnd), .vdd(vdd), .A(_3877_), .B(_3876_), .C(micro_hash_ucr_pipe30_bF_buf2), .Y(_3878_) );
OAI21X1 OAI21X1_1076 ( .gnd(gnd), .vdd(vdd), .A(_913__bF_buf3), .B(micro_hash_ucr_b_2_bF_buf2_), .C(_915__bF_buf0), .Y(_3879_) );
OAI21X1 OAI21X1_1077 ( .gnd(gnd), .vdd(vdd), .A(_3878_), .B(_3879_), .C(_914__bF_buf2), .Y(_3880_) );
AOI21X1 AOI21X1_643 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe32_bF_buf1), .B(_389_), .C(micro_hash_ucr_pipe33_bF_buf2), .Y(_3881_) );
AOI21X1 AOI21X1_644 ( .gnd(gnd), .vdd(vdd), .A(_3881_), .B(_3880_), .C(micro_hash_ucr_pipe34_bF_buf0), .Y(_3882_) );
OAI21X1 OAI21X1_1078 ( .gnd(gnd), .vdd(vdd), .A(_912__bF_buf1), .B(micro_hash_ucr_b_2_bF_buf1_), .C(_911__bF_buf1), .Y(_3883_) );
OAI21X1 OAI21X1_1079 ( .gnd(gnd), .vdd(vdd), .A(_3882_), .B(_3883_), .C(_907__bF_buf1), .Y(_3884_) );
AOI21X1 AOI21X1_645 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe36_bF_buf3), .B(_389_), .C(micro_hash_ucr_pipe37), .Y(_3885_) );
AOI21X1 AOI21X1_646 ( .gnd(gnd), .vdd(vdd), .A(_3885_), .B(_3884_), .C(micro_hash_ucr_pipe38_bF_buf0), .Y(_3886_) );
OAI21X1 OAI21X1_1080 ( .gnd(gnd), .vdd(vdd), .A(_908__bF_buf2), .B(micro_hash_ucr_b_2_bF_buf0_), .C(_904__bF_buf1), .Y(_3887_) );
OAI21X1 OAI21X1_1081 ( .gnd(gnd), .vdd(vdd), .A(_3886_), .B(_3887_), .C(_906__bF_buf4), .Y(_3888_) );
AOI21X1 AOI21X1_647 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe40_bF_buf2), .B(_389_), .C(micro_hash_ucr_pipe41), .Y(_3889_) );
AOI21X1 AOI21X1_648 ( .gnd(gnd), .vdd(vdd), .A(_3889_), .B(_3888_), .C(micro_hash_ucr_pipe42_bF_buf3), .Y(_3890_) );
OAI21X1 OAI21X1_1082 ( .gnd(gnd), .vdd(vdd), .A(_901__bF_buf2), .B(micro_hash_ucr_b_2_bF_buf3_), .C(_903__bF_buf0), .Y(_3891_) );
OAI21X1 OAI21X1_1083 ( .gnd(gnd), .vdd(vdd), .A(_3890_), .B(_3891_), .C(_902__bF_buf3), .Y(_3892_) );
AOI21X1 AOI21X1_649 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe44), .B(_389_), .C(micro_hash_ucr_pipe45_bF_buf3), .Y(_3893_) );
AOI21X1 AOI21X1_650 ( .gnd(gnd), .vdd(vdd), .A(_3893_), .B(_3892_), .C(micro_hash_ucr_pipe46_bF_buf4), .Y(_3894_) );
OAI21X1 OAI21X1_1084 ( .gnd(gnd), .vdd(vdd), .A(_900__bF_buf1), .B(micro_hash_ucr_b_2_bF_buf2_), .C(_899__bF_buf3), .Y(_3895_) );
OAI21X1 OAI21X1_1085 ( .gnd(gnd), .vdd(vdd), .A(_3894_), .B(_3895_), .C(_895__bF_buf3), .Y(_3896_) );
AOI21X1 AOI21X1_651 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe48_bF_buf2), .B(_389_), .C(micro_hash_ucr_pipe49), .Y(_3897_) );
AOI21X1 AOI21X1_652 ( .gnd(gnd), .vdd(vdd), .A(_3897_), .B(_3896_), .C(micro_hash_ucr_pipe50_bF_buf1), .Y(_3898_) );
OAI21X1 OAI21X1_1086 ( .gnd(gnd), .vdd(vdd), .A(_896__bF_buf0), .B(micro_hash_ucr_b_2_bF_buf1_), .C(_892_), .Y(_3899_) );
OAI21X1 OAI21X1_1087 ( .gnd(gnd), .vdd(vdd), .A(_3898_), .B(_3899_), .C(_894__bF_buf1), .Y(_3900_) );
AOI21X1 AOI21X1_653 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe52_bF_buf4), .B(_389_), .C(micro_hash_ucr_pipe53_bF_buf3), .Y(_3901_) );
AOI21X1 AOI21X1_654 ( .gnd(gnd), .vdd(vdd), .A(_3901_), .B(_3900_), .C(micro_hash_ucr_pipe54_bF_buf2), .Y(_3902_) );
OAI21X1 OAI21X1_1088 ( .gnd(gnd), .vdd(vdd), .A(_889__bF_buf2), .B(micro_hash_ucr_b_2_bF_buf0_), .C(_891_), .Y(_3903_) );
OAI21X1 OAI21X1_1089 ( .gnd(gnd), .vdd(vdd), .A(_3902_), .B(_3903_), .C(_890__bF_buf3), .Y(_3904_) );
AOI21X1 AOI21X1_655 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe56_bF_buf2), .B(_389_), .C(micro_hash_ucr_pipe57_bF_buf1), .Y(_3905_) );
AOI21X1 AOI21X1_656 ( .gnd(gnd), .vdd(vdd), .A(_3905_), .B(_3904_), .C(micro_hash_ucr_pipe58_bF_buf0), .Y(_3906_) );
OAI21X1 OAI21X1_1090 ( .gnd(gnd), .vdd(vdd), .A(_888__bF_buf1), .B(micro_hash_ucr_b_2_bF_buf3_), .C(_887__bF_buf3), .Y(_3907_) );
OAI21X1 OAI21X1_1091 ( .gnd(gnd), .vdd(vdd), .A(_3906_), .B(_3907_), .C(_883__bF_buf3), .Y(_3908_) );
AOI21X1 AOI21X1_657 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe60_bF_buf3), .B(_389_), .C(micro_hash_ucr_pipe61_bF_buf3), .Y(_3909_) );
AOI21X1 AOI21X1_658 ( .gnd(gnd), .vdd(vdd), .A(_3909_), .B(_3908_), .C(micro_hash_ucr_pipe62_bF_buf0), .Y(_3910_) );
OAI21X1 OAI21X1_1092 ( .gnd(gnd), .vdd(vdd), .A(_884__bF_buf0), .B(micro_hash_ucr_b_2_bF_buf2_), .C(_880__bF_buf2), .Y(_3911_) );
OAI21X1 OAI21X1_1093 ( .gnd(gnd), .vdd(vdd), .A(_3910_), .B(_3911_), .C(_882__bF_buf2), .Y(_3912_) );
AOI21X1 AOI21X1_659 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe64_bF_buf4), .B(_389_), .C(micro_hash_ucr_pipe65_bF_buf1), .Y(_3913_) );
AOI21X1 AOI21X1_660 ( .gnd(gnd), .vdd(vdd), .A(_3913_), .B(_3912_), .C(micro_hash_ucr_pipe66_bF_buf2), .Y(_3914_) );
OAI21X1 OAI21X1_1094 ( .gnd(gnd), .vdd(vdd), .A(_877__bF_buf3), .B(micro_hash_ucr_b_2_bF_buf1_), .C(_879__bF_buf2), .Y(_3915_) );
OAI21X1 OAI21X1_1095 ( .gnd(gnd), .vdd(vdd), .A(_3914_), .B(_3915_), .C(_878__bF_buf1), .Y(_3916_) );
OAI21X1 OAI21X1_1096 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_2_bF_buf0_), .B(_878__bF_buf0), .C(_3916_), .Y(_3917_) );
NOR2X1 NOR2X1_683 ( .gnd(gnd), .vdd(vdd), .A(_1950_), .B(_3917_), .Y(_298__2_) );
OAI21X1 OAI21X1_1097 ( .gnd(gnd), .vdd(vdd), .A(_1849_), .B(_393_), .C(_947_), .Y(_3918_) );
NOR2X1 NOR2X1_684 ( .gnd(gnd), .vdd(vdd), .A(_3918_), .B(_3744_), .Y(_3919_) );
OAI21X1 OAI21X1_1098 ( .gnd(gnd), .vdd(vdd), .A(_3748_), .B(micro_hash_ucr_b_3_bF_buf2_), .C(_928_), .Y(_3920_) );
OAI21X1 OAI21X1_1099 ( .gnd(gnd), .vdd(vdd), .A(_3919_), .B(_3920_), .C(_930__bF_buf2), .Y(_3921_) );
AOI21X1 AOI21X1_661 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe16_bF_buf2), .B(_394_), .C(micro_hash_ucr_pipe17_bF_buf0), .Y(_3922_) );
AOI21X1 AOI21X1_662 ( .gnd(gnd), .vdd(vdd), .A(_3922_), .B(_3921_), .C(micro_hash_ucr_pipe18_bF_buf1), .Y(_3923_) );
OAI21X1 OAI21X1_1100 ( .gnd(gnd), .vdd(vdd), .A(_925__bF_buf1), .B(micro_hash_ucr_b_3_bF_buf1_), .C(_927__bF_buf2), .Y(_3924_) );
OAI21X1 OAI21X1_1101 ( .gnd(gnd), .vdd(vdd), .A(_3923_), .B(_3924_), .C(_926__bF_buf3), .Y(_3925_) );
AOI21X1 AOI21X1_663 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe20_bF_buf4), .B(_394_), .C(micro_hash_ucr_pipe21_bF_buf2), .Y(_3926_) );
AOI21X1 AOI21X1_664 ( .gnd(gnd), .vdd(vdd), .A(_3926_), .B(_3925_), .C(micro_hash_ucr_pipe22_bF_buf0), .Y(_3927_) );
OAI21X1 OAI21X1_1102 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf2), .B(micro_hash_ucr_b_3_bF_buf0_), .C(_923_), .Y(_3928_) );
OAI21X1 OAI21X1_1103 ( .gnd(gnd), .vdd(vdd), .A(_3927_), .B(_3928_), .C(_919__bF_buf1), .Y(_3929_) );
AOI21X1 AOI21X1_665 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe24_bF_buf1), .B(_394_), .C(micro_hash_ucr_pipe25), .Y(_3930_) );
AOI21X1 AOI21X1_666 ( .gnd(gnd), .vdd(vdd), .A(_3930_), .B(_3929_), .C(micro_hash_ucr_pipe26_bF_buf3), .Y(_3931_) );
OAI21X1 OAI21X1_1104 ( .gnd(gnd), .vdd(vdd), .A(_920__bF_buf1), .B(micro_hash_ucr_b_3_bF_buf3_), .C(_916_), .Y(_3932_) );
OAI21X1 OAI21X1_1105 ( .gnd(gnd), .vdd(vdd), .A(_3931_), .B(_3932_), .C(_918__bF_buf1), .Y(_3933_) );
AOI21X1 AOI21X1_667 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe28_bF_buf2), .B(_394_), .C(micro_hash_ucr_pipe29_bF_buf0), .Y(_3934_) );
AOI21X1 AOI21X1_668 ( .gnd(gnd), .vdd(vdd), .A(_3934_), .B(_3933_), .C(micro_hash_ucr_pipe30_bF_buf1), .Y(_3935_) );
OAI21X1 OAI21X1_1106 ( .gnd(gnd), .vdd(vdd), .A(_913__bF_buf2), .B(micro_hash_ucr_b_3_bF_buf2_), .C(_915__bF_buf3), .Y(_3936_) );
OAI21X1 OAI21X1_1107 ( .gnd(gnd), .vdd(vdd), .A(_3935_), .B(_3936_), .C(_914__bF_buf1), .Y(_3937_) );
AOI21X1 AOI21X1_669 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe32_bF_buf0), .B(_394_), .C(micro_hash_ucr_pipe33_bF_buf1), .Y(_3938_) );
AOI21X1 AOI21X1_670 ( .gnd(gnd), .vdd(vdd), .A(_3938_), .B(_3937_), .C(micro_hash_ucr_pipe34_bF_buf3), .Y(_3939_) );
OAI21X1 OAI21X1_1108 ( .gnd(gnd), .vdd(vdd), .A(_912__bF_buf0), .B(micro_hash_ucr_b_3_bF_buf1_), .C(_911__bF_buf0), .Y(_3940_) );
OAI21X1 OAI21X1_1109 ( .gnd(gnd), .vdd(vdd), .A(_3939_), .B(_3940_), .C(_907__bF_buf0), .Y(_3941_) );
AOI21X1 AOI21X1_671 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe36_bF_buf2), .B(_394_), .C(micro_hash_ucr_pipe37), .Y(_3942_) );
AOI21X1 AOI21X1_672 ( .gnd(gnd), .vdd(vdd), .A(_3942_), .B(_3941_), .C(micro_hash_ucr_pipe38_bF_buf3), .Y(_3943_) );
OAI21X1 OAI21X1_1110 ( .gnd(gnd), .vdd(vdd), .A(_908__bF_buf1), .B(micro_hash_ucr_b_3_bF_buf0_), .C(_904__bF_buf0), .Y(_3944_) );
OAI21X1 OAI21X1_1111 ( .gnd(gnd), .vdd(vdd), .A(_3943_), .B(_3944_), .C(_906__bF_buf3), .Y(_3945_) );
AOI21X1 AOI21X1_673 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe40_bF_buf1), .B(_394_), .C(micro_hash_ucr_pipe41), .Y(_3946_) );
AOI21X1 AOI21X1_674 ( .gnd(gnd), .vdd(vdd), .A(_3946_), .B(_3945_), .C(micro_hash_ucr_pipe42_bF_buf2), .Y(_3947_) );
OAI21X1 OAI21X1_1112 ( .gnd(gnd), .vdd(vdd), .A(_901__bF_buf1), .B(micro_hash_ucr_b_3_bF_buf3_), .C(_903__bF_buf3), .Y(_3948_) );
OAI21X1 OAI21X1_1113 ( .gnd(gnd), .vdd(vdd), .A(_3947_), .B(_3948_), .C(_902__bF_buf2), .Y(_3949_) );
AOI21X1 AOI21X1_675 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe44), .B(_394_), .C(micro_hash_ucr_pipe45_bF_buf2), .Y(_3950_) );
AOI21X1 AOI21X1_676 ( .gnd(gnd), .vdd(vdd), .A(_3950_), .B(_3949_), .C(micro_hash_ucr_pipe46_bF_buf3), .Y(_3951_) );
OAI21X1 OAI21X1_1114 ( .gnd(gnd), .vdd(vdd), .A(_900__bF_buf0), .B(micro_hash_ucr_b_3_bF_buf2_), .C(_899__bF_buf2), .Y(_3952_) );
OAI21X1 OAI21X1_1115 ( .gnd(gnd), .vdd(vdd), .A(_3951_), .B(_3952_), .C(_895__bF_buf2), .Y(_3953_) );
AOI21X1 AOI21X1_677 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe48_bF_buf1), .B(_394_), .C(micro_hash_ucr_pipe49), .Y(_3954_) );
AOI21X1 AOI21X1_678 ( .gnd(gnd), .vdd(vdd), .A(_3954_), .B(_3953_), .C(micro_hash_ucr_pipe50_bF_buf0), .Y(_3955_) );
OAI21X1 OAI21X1_1116 ( .gnd(gnd), .vdd(vdd), .A(_896__bF_buf4), .B(micro_hash_ucr_b_3_bF_buf1_), .C(_892_), .Y(_3956_) );
OAI21X1 OAI21X1_1117 ( .gnd(gnd), .vdd(vdd), .A(_3955_), .B(_3956_), .C(_894__bF_buf0), .Y(_3957_) );
AOI21X1 AOI21X1_679 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe52_bF_buf3), .B(_394_), .C(micro_hash_ucr_pipe53_bF_buf2), .Y(_3958_) );
AOI21X1 AOI21X1_680 ( .gnd(gnd), .vdd(vdd), .A(_3958_), .B(_3957_), .C(micro_hash_ucr_pipe54_bF_buf1), .Y(_3959_) );
OAI21X1 OAI21X1_1118 ( .gnd(gnd), .vdd(vdd), .A(_889__bF_buf1), .B(micro_hash_ucr_b_3_bF_buf0_), .C(_891_), .Y(_3960_) );
OAI21X1 OAI21X1_1119 ( .gnd(gnd), .vdd(vdd), .A(_3959_), .B(_3960_), .C(_890__bF_buf2), .Y(_3961_) );
AOI21X1 AOI21X1_681 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe56_bF_buf1), .B(_394_), .C(micro_hash_ucr_pipe57_bF_buf0), .Y(_3962_) );
AOI21X1 AOI21X1_682 ( .gnd(gnd), .vdd(vdd), .A(_3962_), .B(_3961_), .C(micro_hash_ucr_pipe58_bF_buf4), .Y(_3963_) );
OAI21X1 OAI21X1_1120 ( .gnd(gnd), .vdd(vdd), .A(_888__bF_buf0), .B(micro_hash_ucr_b_3_bF_buf3_), .C(_887__bF_buf2), .Y(_3964_) );
OAI21X1 OAI21X1_1121 ( .gnd(gnd), .vdd(vdd), .A(_3963_), .B(_3964_), .C(_883__bF_buf2), .Y(_3965_) );
AOI21X1 AOI21X1_683 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe60_bF_buf2), .B(_394_), .C(micro_hash_ucr_pipe61_bF_buf2), .Y(_3966_) );
AOI21X1 AOI21X1_684 ( .gnd(gnd), .vdd(vdd), .A(_3966_), .B(_3965_), .C(micro_hash_ucr_pipe62_bF_buf4), .Y(_3967_) );
OAI21X1 OAI21X1_1122 ( .gnd(gnd), .vdd(vdd), .A(_884__bF_buf4), .B(micro_hash_ucr_b_3_bF_buf2_), .C(_880__bF_buf1), .Y(_3968_) );
OAI21X1 OAI21X1_1123 ( .gnd(gnd), .vdd(vdd), .A(_3967_), .B(_3968_), .C(_882__bF_buf1), .Y(_3969_) );
AOI21X1 AOI21X1_685 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe64_bF_buf3), .B(_394_), .C(micro_hash_ucr_pipe65_bF_buf0), .Y(_3970_) );
AOI21X1 AOI21X1_686 ( .gnd(gnd), .vdd(vdd), .A(_3970_), .B(_3969_), .C(micro_hash_ucr_pipe66_bF_buf1), .Y(_3971_) );
OAI21X1 OAI21X1_1124 ( .gnd(gnd), .vdd(vdd), .A(_877__bF_buf2), .B(micro_hash_ucr_b_3_bF_buf1_), .C(_879__bF_buf1), .Y(_3972_) );
OAI21X1 OAI21X1_1125 ( .gnd(gnd), .vdd(vdd), .A(_3971_), .B(_3972_), .C(_878__bF_buf4), .Y(_3973_) );
OAI21X1 OAI21X1_1126 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_3_bF_buf0_), .B(_878__bF_buf3), .C(_3973_), .Y(_3974_) );
NOR2X1 NOR2X1_685 ( .gnd(gnd), .vdd(vdd), .A(_1950_), .B(_3974_), .Y(_298__3_) );
NAND2X1 NAND2X1_462 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_4_bF_buf2_), .B(micro_hash_ucr_pipe66_bF_buf0), .Y(_3975_) );
NOR2X1 NOR2X1_686 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_4_bF_buf1_), .B(_882__bF_buf0), .Y(_3976_) );
NAND2X1 NAND2X1_463 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe63), .B(_4423__bF_buf0), .Y(_3977_) );
NOR2X1 NOR2X1_687 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_4_bF_buf0_), .B(_884__bF_buf3), .Y(_3978_) );
NAND2X1 NAND2X1_464 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe61_bF_buf1), .B(_4423__bF_buf3), .Y(_3979_) );
NOR2X1 NOR2X1_688 ( .gnd(gnd), .vdd(vdd), .A(_1395_), .B(_894__bF_buf3), .Y(_3980_) );
NAND2X1 NAND2X1_465 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_0_bF_buf3_), .B(micro_hash_ucr_pipe51), .Y(_3981_) );
NOR2X1 NOR2X1_689 ( .gnd(gnd), .vdd(vdd), .A(_1395_), .B(_896__bF_buf3), .Y(_3982_) );
NAND2X1 NAND2X1_466 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_0_bF_buf2_), .B(micro_hash_ucr_pipe49), .Y(_3983_) );
NOR2X1 NOR2X1_690 ( .gnd(gnd), .vdd(vdd), .A(_1395_), .B(_895__bF_buf1), .Y(_3984_) );
NAND2X1 NAND2X1_467 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_0_bF_buf1_), .B(micro_hash_ucr_pipe47), .Y(_3985_) );
NOR2X1 NOR2X1_691 ( .gnd(gnd), .vdd(vdd), .A(_1395_), .B(_900__bF_buf3), .Y(_3986_) );
NAND2X1 NAND2X1_468 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_0_bF_buf0_), .B(micro_hash_ucr_pipe45_bF_buf1), .Y(_3987_) );
NAND2X1 NAND2X1_469 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_4_bF_buf3_), .B(micro_hash_ucr_pipe32_bF_buf3), .Y(_3988_) );
NAND2X1 NAND2X1_470 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_4_bF_buf2_), .B(micro_hash_ucr_pipe30_bF_buf0), .Y(_3989_) );
NAND2X1 NAND2X1_471 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_0_bF_buf3_), .B(micro_hash_ucr_pipe23_bF_buf0), .Y(_3990_) );
NAND2X1 NAND2X1_472 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_0_bF_buf2_), .B(micro_hash_ucr_pipe21_bF_buf1), .Y(_3991_) );
NAND2X1 NAND2X1_473 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_0_bF_buf1_), .B(micro_hash_ucr_pipe19_bF_buf3), .Y(_3992_) );
NAND2X1 NAND2X1_474 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_0_bF_buf0_), .B(micro_hash_ucr_pipe17_bF_buf3), .Y(_3993_) );
NAND2X1 NAND2X1_475 ( .gnd(gnd), .vdd(vdd), .A(_4423__bF_buf2), .B(_1071_), .Y(_3994_) );
NOR2X1 NOR2X1_692 ( .gnd(gnd), .vdd(vdd), .A(H_12_), .B(micro_hash_ucr_pipe12), .Y(_3995_) );
NAND3X1 NAND3X1_124 ( .gnd(gnd), .vdd(vdd), .A(_935_), .B(_936_), .C(_3995_), .Y(_3996_) );
NAND3X1 NAND3X1_125 ( .gnd(gnd), .vdd(vdd), .A(_932_), .B(_933_), .C(_965_), .Y(_3997_) );
OR2X2 OR2X2_43 ( .gnd(gnd), .vdd(vdd), .A(_3996_), .B(_3997_), .Y(_3998_) );
OAI22X1 OAI22X1_58 ( .gnd(gnd), .vdd(vdd), .A(_955_), .B(_3998_), .C(_1079_), .D(micro_hash_ucr_b_4_bF_buf1_), .Y(_3999_) );
AOI21X1 AOI21X1_687 ( .gnd(gnd), .vdd(vdd), .A(_928_), .B(_3999_), .C(micro_hash_ucr_pipe16_bF_buf1), .Y(_4000_) );
AOI22X1 AOI22X1_35 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_4_bF_buf0_), .B(micro_hash_ucr_pipe16_bF_buf0), .C(_4000_), .D(_3994_), .Y(_4001_) );
OAI21X1 OAI21X1_1127 ( .gnd(gnd), .vdd(vdd), .A(_4001_), .B(micro_hash_ucr_pipe17_bF_buf2), .C(_3993_), .Y(_4002_) );
NAND2X1 NAND2X1_476 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe18_bF_buf0), .B(_1395_), .Y(_4003_) );
OAI21X1 OAI21X1_1128 ( .gnd(gnd), .vdd(vdd), .A(_4002_), .B(micro_hash_ucr_pipe18_bF_buf4), .C(_4003_), .Y(_4004_) );
OAI21X1 OAI21X1_1129 ( .gnd(gnd), .vdd(vdd), .A(_4004_), .B(micro_hash_ucr_pipe19_bF_buf2), .C(_3992_), .Y(_4005_) );
NAND2X1 NAND2X1_477 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe20_bF_buf3), .B(_1395_), .Y(_4006_) );
OAI21X1 OAI21X1_1130 ( .gnd(gnd), .vdd(vdd), .A(_4005_), .B(micro_hash_ucr_pipe20_bF_buf2), .C(_4006_), .Y(_4007_) );
OAI21X1 OAI21X1_1131 ( .gnd(gnd), .vdd(vdd), .A(_4007_), .B(micro_hash_ucr_pipe21_bF_buf0), .C(_3991_), .Y(_4008_) );
NAND2X1 NAND2X1_478 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe22_bF_buf4), .B(_1395_), .Y(_4009_) );
OAI21X1 OAI21X1_1132 ( .gnd(gnd), .vdd(vdd), .A(_4008_), .B(micro_hash_ucr_pipe22_bF_buf3), .C(_4009_), .Y(_4010_) );
OAI21X1 OAI21X1_1133 ( .gnd(gnd), .vdd(vdd), .A(_4010_), .B(micro_hash_ucr_pipe23_bF_buf3), .C(_3990_), .Y(_4011_) );
NAND2X1 NAND2X1_479 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe24_bF_buf0), .B(_1395_), .Y(_4012_) );
OAI21X1 OAI21X1_1134 ( .gnd(gnd), .vdd(vdd), .A(_4011_), .B(micro_hash_ucr_pipe24_bF_buf4), .C(_4012_), .Y(_4013_) );
NOR2X1 NOR2X1_693 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe25), .B(_4013_), .Y(_4014_) );
OAI21X1 OAI21X1_1135 ( .gnd(gnd), .vdd(vdd), .A(_4423__bF_buf1), .B(_921__bF_buf1), .C(_920__bF_buf0), .Y(_4015_) );
AOI21X1 AOI21X1_688 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe26_bF_buf2), .B(_1395_), .C(micro_hash_ucr_pipe27), .Y(_4016_) );
OAI21X1 OAI21X1_1136 ( .gnd(gnd), .vdd(vdd), .A(_4014_), .B(_4015_), .C(_4016_), .Y(_4017_) );
OAI21X1 OAI21X1_1137 ( .gnd(gnd), .vdd(vdd), .A(_4423__bF_buf0), .B(_916_), .C(_4017_), .Y(_4018_) );
NAND2X1 NAND2X1_480 ( .gnd(gnd), .vdd(vdd), .A(_918__bF_buf0), .B(_4018_), .Y(_4019_) );
OAI21X1 OAI21X1_1138 ( .gnd(gnd), .vdd(vdd), .A(_1395_), .B(_918__bF_buf4), .C(_4019_), .Y(_4020_) );
NAND2X1 NAND2X1_481 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe29_bF_buf3), .B(_4423__bF_buf3), .Y(_4021_) );
OAI21X1 OAI21X1_1139 ( .gnd(gnd), .vdd(vdd), .A(_4020_), .B(micro_hash_ucr_pipe29_bF_buf2), .C(_4021_), .Y(_4022_) );
OAI21X1 OAI21X1_1140 ( .gnd(gnd), .vdd(vdd), .A(_4022_), .B(micro_hash_ucr_pipe30_bF_buf3), .C(_3989_), .Y(_4023_) );
NAND2X1 NAND2X1_482 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe31), .B(_4423__bF_buf2), .Y(_4024_) );
OAI21X1 OAI21X1_1141 ( .gnd(gnd), .vdd(vdd), .A(_4023_), .B(micro_hash_ucr_pipe31), .C(_4024_), .Y(_4025_) );
OAI21X1 OAI21X1_1142 ( .gnd(gnd), .vdd(vdd), .A(_4025_), .B(micro_hash_ucr_pipe32_bF_buf2), .C(_3988_), .Y(_4026_) );
NAND2X1 NAND2X1_483 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe33_bF_buf0), .B(_4423__bF_buf1), .Y(_4027_) );
OAI21X1 OAI21X1_1143 ( .gnd(gnd), .vdd(vdd), .A(_4026_), .B(micro_hash_ucr_pipe33_bF_buf3), .C(_4027_), .Y(_4028_) );
OAI21X1 OAI21X1_1144 ( .gnd(gnd), .vdd(vdd), .A(_912__bF_buf4), .B(micro_hash_ucr_b_4_bF_buf3_), .C(_911__bF_buf4), .Y(_4029_) );
AOI21X1 AOI21X1_689 ( .gnd(gnd), .vdd(vdd), .A(_912__bF_buf3), .B(_4028_), .C(_4029_), .Y(_4030_) );
OAI21X1 OAI21X1_1145 ( .gnd(gnd), .vdd(vdd), .A(_4423__bF_buf0), .B(_911__bF_buf3), .C(_907__bF_buf4), .Y(_4031_) );
OAI22X1 OAI22X1_59 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_4_bF_buf2_), .B(_907__bF_buf3), .C(_4030_), .D(_4031_), .Y(_4032_) );
OAI21X1 OAI21X1_1146 ( .gnd(gnd), .vdd(vdd), .A(_909__bF_buf0), .B(micro_hash_ucr_c_0_bF_buf3_), .C(_908__bF_buf0), .Y(_4033_) );
AOI21X1 AOI21X1_690 ( .gnd(gnd), .vdd(vdd), .A(_909__bF_buf3), .B(_4032_), .C(_4033_), .Y(_4034_) );
NOR2X1 NOR2X1_694 ( .gnd(gnd), .vdd(vdd), .A(_1395_), .B(_908__bF_buf4), .Y(_4035_) );
OAI21X1 OAI21X1_1147 ( .gnd(gnd), .vdd(vdd), .A(_4034_), .B(_4035_), .C(_904__bF_buf3), .Y(_4036_) );
AOI21X1 AOI21X1_691 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_0_bF_buf2_), .B(micro_hash_ucr_pipe39), .C(micro_hash_ucr_pipe40_bF_buf0), .Y(_4037_) );
OAI21X1 OAI21X1_1148 ( .gnd(gnd), .vdd(vdd), .A(_906__bF_buf2), .B(micro_hash_ucr_b_4_bF_buf1_), .C(_905__bF_buf0), .Y(_4038_) );
AOI21X1 AOI21X1_692 ( .gnd(gnd), .vdd(vdd), .A(_4037_), .B(_4036_), .C(_4038_), .Y(_4039_) );
OAI21X1 OAI21X1_1149 ( .gnd(gnd), .vdd(vdd), .A(_4423__bF_buf3), .B(_905__bF_buf3), .C(_901__bF_buf0), .Y(_4040_) );
OAI22X1 OAI22X1_60 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_4_bF_buf0_), .B(_901__bF_buf4), .C(_4039_), .D(_4040_), .Y(_4041_) );
OAI21X1 OAI21X1_1150 ( .gnd(gnd), .vdd(vdd), .A(_903__bF_buf2), .B(micro_hash_ucr_c_0_bF_buf1_), .C(_902__bF_buf1), .Y(_4042_) );
AOI21X1 AOI21X1_693 ( .gnd(gnd), .vdd(vdd), .A(_903__bF_buf1), .B(_4041_), .C(_4042_), .Y(_4043_) );
NOR2X1 NOR2X1_695 ( .gnd(gnd), .vdd(vdd), .A(_1395_), .B(_902__bF_buf0), .Y(_4044_) );
OAI21X1 OAI21X1_1151 ( .gnd(gnd), .vdd(vdd), .A(_4043_), .B(_4044_), .C(_898_), .Y(_4045_) );
AOI21X1 AOI21X1_694 ( .gnd(gnd), .vdd(vdd), .A(_3987_), .B(_4045_), .C(micro_hash_ucr_pipe46_bF_buf2), .Y(_4046_) );
OAI21X1 OAI21X1_1152 ( .gnd(gnd), .vdd(vdd), .A(_4046_), .B(_3986_), .C(_899__bF_buf1), .Y(_4047_) );
AOI21X1 AOI21X1_695 ( .gnd(gnd), .vdd(vdd), .A(_3985_), .B(_4047_), .C(micro_hash_ucr_pipe48_bF_buf0), .Y(_4048_) );
OAI21X1 OAI21X1_1153 ( .gnd(gnd), .vdd(vdd), .A(_4048_), .B(_3984_), .C(_897__bF_buf1), .Y(_4049_) );
AOI21X1 AOI21X1_696 ( .gnd(gnd), .vdd(vdd), .A(_3983_), .B(_4049_), .C(micro_hash_ucr_pipe50_bF_buf3), .Y(_4050_) );
OAI21X1 OAI21X1_1154 ( .gnd(gnd), .vdd(vdd), .A(_4050_), .B(_3982_), .C(_892_), .Y(_4051_) );
AOI21X1 AOI21X1_697 ( .gnd(gnd), .vdd(vdd), .A(_3981_), .B(_4051_), .C(micro_hash_ucr_pipe52_bF_buf2), .Y(_4052_) );
OAI21X1 OAI21X1_1155 ( .gnd(gnd), .vdd(vdd), .A(_4052_), .B(_3980_), .C(_893_), .Y(_4053_) );
AOI21X1 AOI21X1_698 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_0_bF_buf0_), .B(micro_hash_ucr_pipe53_bF_buf1), .C(micro_hash_ucr_pipe54_bF_buf0), .Y(_4054_) );
OAI21X1 OAI21X1_1156 ( .gnd(gnd), .vdd(vdd), .A(_889__bF_buf0), .B(micro_hash_ucr_b_4_bF_buf3_), .C(_891_), .Y(_4055_) );
AOI21X1 AOI21X1_699 ( .gnd(gnd), .vdd(vdd), .A(_4054_), .B(_4053_), .C(_4055_), .Y(_4056_) );
OAI21X1 OAI21X1_1157 ( .gnd(gnd), .vdd(vdd), .A(_4423__bF_buf2), .B(_891_), .C(_890__bF_buf1), .Y(_4057_) );
OAI22X1 OAI22X1_61 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_4_bF_buf2_), .B(_890__bF_buf0), .C(_4056_), .D(_4057_), .Y(_4058_) );
AOI21X1 AOI21X1_700 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_0_bF_buf3_), .B(micro_hash_ucr_pipe57_bF_buf3), .C(micro_hash_ucr_pipe58_bF_buf3), .Y(_4059_) );
OAI21X1 OAI21X1_1158 ( .gnd(gnd), .vdd(vdd), .A(_4058_), .B(micro_hash_ucr_pipe57_bF_buf2), .C(_4059_), .Y(_4060_) );
AOI21X1 AOI21X1_701 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe58_bF_buf2), .B(_1395_), .C(micro_hash_ucr_pipe59), .Y(_4061_) );
OAI21X1 OAI21X1_1159 ( .gnd(gnd), .vdd(vdd), .A(_4423__bF_buf1), .B(_887__bF_buf1), .C(_883__bF_buf1), .Y(_4062_) );
AOI21X1 AOI21X1_702 ( .gnd(gnd), .vdd(vdd), .A(_4061_), .B(_4060_), .C(_4062_), .Y(_4063_) );
NOR2X1 NOR2X1_696 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_4_bF_buf1_), .B(_883__bF_buf0), .Y(_4064_) );
OAI21X1 OAI21X1_1160 ( .gnd(gnd), .vdd(vdd), .A(_4063_), .B(_4064_), .C(_885_), .Y(_4065_) );
AOI21X1 AOI21X1_703 ( .gnd(gnd), .vdd(vdd), .A(_3979_), .B(_4065_), .C(micro_hash_ucr_pipe62_bF_buf3), .Y(_4066_) );
OAI21X1 OAI21X1_1161 ( .gnd(gnd), .vdd(vdd), .A(_4066_), .B(_3978_), .C(_880__bF_buf0), .Y(_4067_) );
AOI21X1 AOI21X1_704 ( .gnd(gnd), .vdd(vdd), .A(_3977_), .B(_4067_), .C(micro_hash_ucr_pipe64_bF_buf2), .Y(_4068_) );
OAI21X1 OAI21X1_1162 ( .gnd(gnd), .vdd(vdd), .A(_4068_), .B(_3976_), .C(_881_), .Y(_4069_) );
OAI21X1 OAI21X1_1163 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_0_bF_buf2_), .B(_881_), .C(_4069_), .Y(_4070_) );
OAI21X1 OAI21X1_1164 ( .gnd(gnd), .vdd(vdd), .A(_4070_), .B(micro_hash_ucr_pipe66_bF_buf4), .C(_3975_), .Y(_4071_) );
OAI21X1 OAI21X1_1165 ( .gnd(gnd), .vdd(vdd), .A(_4423__bF_buf0), .B(_879__bF_buf0), .C(_878__bF_buf2), .Y(_4072_) );
AOI21X1 AOI21X1_705 ( .gnd(gnd), .vdd(vdd), .A(_879__bF_buf3), .B(_4071_), .C(_4072_), .Y(_4073_) );
OAI21X1 OAI21X1_1166 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_4_bF_buf0_), .B(_878__bF_buf1), .C(_1949_), .Y(_4074_) );
OAI22X1 OAI22X1_62 ( .gnd(gnd), .vdd(vdd), .A(_4423__bF_buf3), .B(_3093_), .C(_4073_), .D(_4074_), .Y(_298__4_) );
NAND2X1 NAND2X1_484 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe64_bF_buf1), .B(_414__bF_buf1), .Y(_4075_) );
NAND2X1 NAND2X1_485 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_1_bF_buf3_), .B(micro_hash_ucr_pipe63), .Y(_4076_) );
NAND2X1 NAND2X1_486 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe62_bF_buf2), .B(_414__bF_buf0), .Y(_4077_) );
NAND2X1 NAND2X1_487 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_1_bF_buf2_), .B(micro_hash_ucr_pipe61_bF_buf0), .Y(_4078_) );
NAND2X1 NAND2X1_488 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe60_bF_buf1), .B(_414__bF_buf3), .Y(_4079_) );
NAND2X1 NAND2X1_489 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_1_bF_buf1_), .B(micro_hash_ucr_pipe59), .Y(_4080_) );
NAND2X1 NAND2X1_490 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe58_bF_buf1), .B(_414__bF_buf2), .Y(_4081_) );
NAND2X1 NAND2X1_491 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_1_bF_buf0_), .B(micro_hash_ucr_pipe57_bF_buf1), .Y(_4082_) );
NAND2X1 NAND2X1_492 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe56_bF_buf0), .B(_414__bF_buf1), .Y(_4083_) );
NAND2X1 NAND2X1_493 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_1_bF_buf3_), .B(micro_hash_ucr_pipe55), .Y(_4084_) );
NAND2X1 NAND2X1_494 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_1_bF_buf2_), .B(micro_hash_ucr_pipe51), .Y(_4085_) );
NAND2X1 NAND2X1_495 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe46_bF_buf1), .B(_414__bF_buf0), .Y(_4086_) );
NOR2X1 NOR2X1_697 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_1_bF_buf1_), .B(_898_), .Y(_4087_) );
NAND2X1 NAND2X1_496 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_5_bF_buf2_), .B(micro_hash_ucr_pipe36_bF_buf1), .Y(_4088_) );
NOR2X1 NOR2X1_698 ( .gnd(gnd), .vdd(vdd), .A(_1058__bF_buf1), .B(_911__bF_buf2), .Y(_4089_) );
NAND2X1 NAND2X1_497 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_5_bF_buf1_), .B(micro_hash_ucr_pipe34_bF_buf2), .Y(_4090_) );
NOR2X1 NOR2X1_699 ( .gnd(gnd), .vdd(vdd), .A(_1058__bF_buf0), .B(_910_), .Y(_4091_) );
NAND2X1 NAND2X1_498 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_5_bF_buf0_), .B(micro_hash_ucr_pipe28_bF_buf1), .Y(_4092_) );
NAND2X1 NAND2X1_499 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_5_bF_buf3_), .B(micro_hash_ucr_pipe26_bF_buf1), .Y(_4093_) );
NAND2X1 NAND2X1_500 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_5_bF_buf2_), .B(micro_hash_ucr_pipe16_bF_buf3), .Y(_4094_) );
NOR2X1 NOR2X1_700 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe6), .B(micro_hash_ucr_pipe7), .Y(_4095_) );
NOR3X1 NOR3X1_4 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe9), .B(micro_hash_ucr_pipe8), .C(_4095_), .Y(_4096_) );
NOR2X1 NOR2X1_701 ( .gnd(gnd), .vdd(vdd), .A(H_13_), .B(micro_hash_ucr_pipe11), .Y(_4097_) );
NOR2X1 NOR2X1_702 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe10), .B(micro_hash_ucr_pipe7), .Y(_4098_) );
NAND3X1 NAND3X1_126 ( .gnd(gnd), .vdd(vdd), .A(_4097_), .B(_4098_), .C(_4096_), .Y(_4099_) );
OAI21X1 OAI21X1_1167 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_1_bF_buf0_), .B(_968_), .C(_4099_), .Y(_4100_) );
AOI22X1 AOI22X1_36 ( .gnd(gnd), .vdd(vdd), .A(_414__bF_buf3), .B(_957_), .C(_4100_), .D(_931_), .Y(_4101_) );
NAND2X1 NAND2X1_501 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe13), .B(_1058__bF_buf3), .Y(_4102_) );
OAI21X1 OAI21X1_1168 ( .gnd(gnd), .vdd(vdd), .A(_4101_), .B(micro_hash_ucr_pipe13), .C(_4102_), .Y(_4103_) );
NAND2X1 NAND2X1_502 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_5_bF_buf1_), .B(micro_hash_ucr_pipe14_bF_buf3), .Y(_4104_) );
OAI21X1 OAI21X1_1169 ( .gnd(gnd), .vdd(vdd), .A(_4103_), .B(micro_hash_ucr_pipe14_bF_buf2), .C(_4104_), .Y(_4105_) );
NAND2X1 NAND2X1_503 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe15_bF_buf0), .B(_1058__bF_buf2), .Y(_4106_) );
OAI21X1 OAI21X1_1170 ( .gnd(gnd), .vdd(vdd), .A(_4105_), .B(micro_hash_ucr_pipe15_bF_buf3), .C(_4106_), .Y(_4107_) );
OAI21X1 OAI21X1_1171 ( .gnd(gnd), .vdd(vdd), .A(_4107_), .B(micro_hash_ucr_pipe16_bF_buf2), .C(_4094_), .Y(_4108_) );
NAND2X1 NAND2X1_504 ( .gnd(gnd), .vdd(vdd), .A(_929_), .B(_4108_), .Y(_4109_) );
OAI21X1 OAI21X1_1172 ( .gnd(gnd), .vdd(vdd), .A(_1058__bF_buf1), .B(_929_), .C(_4109_), .Y(_4110_) );
AOI21X1 AOI21X1_706 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe18_bF_buf3), .B(_414__bF_buf2), .C(micro_hash_ucr_pipe19_bF_buf1), .Y(_4111_) );
OAI21X1 OAI21X1_1173 ( .gnd(gnd), .vdd(vdd), .A(_4110_), .B(micro_hash_ucr_pipe18_bF_buf2), .C(_4111_), .Y(_4112_) );
OAI21X1 OAI21X1_1174 ( .gnd(gnd), .vdd(vdd), .A(_1058__bF_buf0), .B(_927__bF_buf1), .C(_4112_), .Y(_4113_) );
NAND2X1 NAND2X1_505 ( .gnd(gnd), .vdd(vdd), .A(_926__bF_buf2), .B(_4113_), .Y(_4114_) );
OAI21X1 OAI21X1_1175 ( .gnd(gnd), .vdd(vdd), .A(_414__bF_buf1), .B(_926__bF_buf1), .C(_4114_), .Y(_4115_) );
NAND2X1 NAND2X1_506 ( .gnd(gnd), .vdd(vdd), .A(_922_), .B(_4115_), .Y(_4116_) );
OAI21X1 OAI21X1_1176 ( .gnd(gnd), .vdd(vdd), .A(_1058__bF_buf3), .B(_922_), .C(_4116_), .Y(_4117_) );
AOI21X1 AOI21X1_707 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe22_bF_buf2), .B(_414__bF_buf0), .C(micro_hash_ucr_pipe23_bF_buf2), .Y(_4118_) );
OAI21X1 OAI21X1_1177 ( .gnd(gnd), .vdd(vdd), .A(_4117_), .B(micro_hash_ucr_pipe22_bF_buf1), .C(_4118_), .Y(_4119_) );
AOI21X1 AOI21X1_708 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_1_bF_buf3_), .B(micro_hash_ucr_pipe23_bF_buf1), .C(micro_hash_ucr_pipe24_bF_buf3), .Y(_4120_) );
AOI22X1 AOI22X1_37 ( .gnd(gnd), .vdd(vdd), .A(_414__bF_buf3), .B(micro_hash_ucr_pipe24_bF_buf2), .C(_4119_), .D(_4120_), .Y(_4121_) );
NAND2X1 NAND2X1_507 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe25), .B(_1058__bF_buf2), .Y(_4122_) );
OAI21X1 OAI21X1_1178 ( .gnd(gnd), .vdd(vdd), .A(_4121_), .B(micro_hash_ucr_pipe25), .C(_4122_), .Y(_4123_) );
OAI21X1 OAI21X1_1179 ( .gnd(gnd), .vdd(vdd), .A(_4123_), .B(micro_hash_ucr_pipe26_bF_buf0), .C(_4093_), .Y(_4124_) );
NAND2X1 NAND2X1_508 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe27), .B(_1058__bF_buf1), .Y(_4125_) );
OAI21X1 OAI21X1_1180 ( .gnd(gnd), .vdd(vdd), .A(_4124_), .B(micro_hash_ucr_pipe27), .C(_4125_), .Y(_4126_) );
OAI21X1 OAI21X1_1181 ( .gnd(gnd), .vdd(vdd), .A(_4126_), .B(micro_hash_ucr_pipe28_bF_buf0), .C(_4092_), .Y(_4127_) );
NAND2X1 NAND2X1_509 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe29_bF_buf1), .B(_1058__bF_buf0), .Y(_4128_) );
OAI21X1 OAI21X1_1182 ( .gnd(gnd), .vdd(vdd), .A(_4127_), .B(micro_hash_ucr_pipe29_bF_buf0), .C(_4128_), .Y(_4129_) );
NOR2X1 NOR2X1_703 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe30_bF_buf2), .B(_4129_), .Y(_4130_) );
OAI21X1 OAI21X1_1183 ( .gnd(gnd), .vdd(vdd), .A(_414__bF_buf2), .B(_913__bF_buf1), .C(_915__bF_buf2), .Y(_4131_) );
AOI21X1 AOI21X1_709 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe31), .B(_1058__bF_buf3), .C(micro_hash_ucr_pipe32_bF_buf1), .Y(_4132_) );
OAI21X1 OAI21X1_1184 ( .gnd(gnd), .vdd(vdd), .A(_4130_), .B(_4131_), .C(_4132_), .Y(_4133_) );
NAND2X1 NAND2X1_510 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_5_bF_buf0_), .B(micro_hash_ucr_pipe32_bF_buf0), .Y(_4134_) );
AOI21X1 AOI21X1_710 ( .gnd(gnd), .vdd(vdd), .A(_4134_), .B(_4133_), .C(micro_hash_ucr_pipe33_bF_buf2), .Y(_4135_) );
OAI21X1 OAI21X1_1185 ( .gnd(gnd), .vdd(vdd), .A(_4135_), .B(_4091_), .C(_912__bF_buf2), .Y(_4136_) );
AOI21X1 AOI21X1_711 ( .gnd(gnd), .vdd(vdd), .A(_4090_), .B(_4136_), .C(micro_hash_ucr_pipe35), .Y(_4137_) );
OAI21X1 OAI21X1_1186 ( .gnd(gnd), .vdd(vdd), .A(_4137_), .B(_4089_), .C(_907__bF_buf2), .Y(_4138_) );
AOI21X1 AOI21X1_712 ( .gnd(gnd), .vdd(vdd), .A(_4088_), .B(_4138_), .C(micro_hash_ucr_pipe37), .Y(_4139_) );
OAI21X1 OAI21X1_1187 ( .gnd(gnd), .vdd(vdd), .A(_1058__bF_buf2), .B(_909__bF_buf2), .C(_908__bF_buf3), .Y(_4140_) );
AOI21X1 AOI21X1_713 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe38_bF_buf2), .B(_414__bF_buf1), .C(micro_hash_ucr_pipe39), .Y(_4141_) );
OAI21X1 OAI21X1_1188 ( .gnd(gnd), .vdd(vdd), .A(_4139_), .B(_4140_), .C(_4141_), .Y(_4142_) );
AOI21X1 AOI21X1_714 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_1_bF_buf2_), .B(micro_hash_ucr_pipe39), .C(micro_hash_ucr_pipe40_bF_buf4), .Y(_4143_) );
AOI22X1 AOI22X1_38 ( .gnd(gnd), .vdd(vdd), .A(_414__bF_buf0), .B(micro_hash_ucr_pipe40_bF_buf3), .C(_4142_), .D(_4143_), .Y(_4144_) );
OAI21X1 OAI21X1_1189 ( .gnd(gnd), .vdd(vdd), .A(_1058__bF_buf1), .B(_905__bF_buf2), .C(_901__bF_buf3), .Y(_4145_) );
AOI21X1 AOI21X1_715 ( .gnd(gnd), .vdd(vdd), .A(_905__bF_buf1), .B(_4144_), .C(_4145_), .Y(_4146_) );
OAI21X1 OAI21X1_1190 ( .gnd(gnd), .vdd(vdd), .A(_901__bF_buf2), .B(micro_hash_ucr_b_5_bF_buf3_), .C(_903__bF_buf0), .Y(_4147_) );
AOI21X1 AOI21X1_716 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_1_bF_buf1_), .B(micro_hash_ucr_pipe43), .C(micro_hash_ucr_pipe44), .Y(_4148_) );
OAI21X1 OAI21X1_1191 ( .gnd(gnd), .vdd(vdd), .A(_4146_), .B(_4147_), .C(_4148_), .Y(_4149_) );
NAND2X1 NAND2X1_511 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe44), .B(_414__bF_buf3), .Y(_4150_) );
AOI21X1 AOI21X1_717 ( .gnd(gnd), .vdd(vdd), .A(_4150_), .B(_4149_), .C(micro_hash_ucr_pipe45_bF_buf0), .Y(_4151_) );
OAI21X1 OAI21X1_1192 ( .gnd(gnd), .vdd(vdd), .A(_4151_), .B(_4087_), .C(_900__bF_buf2), .Y(_4152_) );
NAND3X1 NAND3X1_127 ( .gnd(gnd), .vdd(vdd), .A(_899__bF_buf0), .B(_4086_), .C(_4152_), .Y(_4153_) );
AOI21X1 AOI21X1_718 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_1_bF_buf0_), .B(micro_hash_ucr_pipe47), .C(micro_hash_ucr_pipe48_bF_buf3), .Y(_4154_) );
OAI21X1 OAI21X1_1193 ( .gnd(gnd), .vdd(vdd), .A(_895__bF_buf0), .B(micro_hash_ucr_b_5_bF_buf2_), .C(_897__bF_buf0), .Y(_4155_) );
AOI21X1 AOI21X1_719 ( .gnd(gnd), .vdd(vdd), .A(_4154_), .B(_4153_), .C(_4155_), .Y(_4156_) );
OAI21X1 OAI21X1_1194 ( .gnd(gnd), .vdd(vdd), .A(_1058__bF_buf0), .B(_897__bF_buf3), .C(_896__bF_buf2), .Y(_4157_) );
OAI22X1 OAI22X1_63 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_5_bF_buf1_), .B(_896__bF_buf1), .C(_4156_), .D(_4157_), .Y(_4158_) );
OAI21X1 OAI21X1_1195 ( .gnd(gnd), .vdd(vdd), .A(_4158_), .B(micro_hash_ucr_pipe51), .C(_4085_), .Y(_4159_) );
NAND2X1 NAND2X1_512 ( .gnd(gnd), .vdd(vdd), .A(_894__bF_buf2), .B(_4159_), .Y(_4160_) );
AOI21X1 AOI21X1_720 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_5_bF_buf0_), .B(micro_hash_ucr_pipe52_bF_buf1), .C(micro_hash_ucr_pipe53_bF_buf0), .Y(_4161_) );
OAI21X1 OAI21X1_1196 ( .gnd(gnd), .vdd(vdd), .A(_893_), .B(micro_hash_ucr_c_1_bF_buf3_), .C(_889__bF_buf4), .Y(_4162_) );
AOI21X1 AOI21X1_721 ( .gnd(gnd), .vdd(vdd), .A(_4161_), .B(_4160_), .C(_4162_), .Y(_4163_) );
NOR2X1 NOR2X1_704 ( .gnd(gnd), .vdd(vdd), .A(_414__bF_buf2), .B(_889__bF_buf3), .Y(_4164_) );
OAI21X1 OAI21X1_1197 ( .gnd(gnd), .vdd(vdd), .A(_4163_), .B(_4164_), .C(_891_), .Y(_4165_) );
NAND3X1 NAND3X1_128 ( .gnd(gnd), .vdd(vdd), .A(_890__bF_buf4), .B(_4084_), .C(_4165_), .Y(_4166_) );
NAND3X1 NAND3X1_129 ( .gnd(gnd), .vdd(vdd), .A(_886_), .B(_4083_), .C(_4166_), .Y(_4167_) );
NAND3X1 NAND3X1_130 ( .gnd(gnd), .vdd(vdd), .A(_888__bF_buf3), .B(_4082_), .C(_4167_), .Y(_4168_) );
NAND3X1 NAND3X1_131 ( .gnd(gnd), .vdd(vdd), .A(_887__bF_buf0), .B(_4081_), .C(_4168_), .Y(_4169_) );
NAND3X1 NAND3X1_132 ( .gnd(gnd), .vdd(vdd), .A(_883__bF_buf3), .B(_4080_), .C(_4169_), .Y(_4170_) );
NAND3X1 NAND3X1_133 ( .gnd(gnd), .vdd(vdd), .A(_885_), .B(_4079_), .C(_4170_), .Y(_4171_) );
NAND3X1 NAND3X1_134 ( .gnd(gnd), .vdd(vdd), .A(_884__bF_buf2), .B(_4078_), .C(_4171_), .Y(_4172_) );
NAND3X1 NAND3X1_135 ( .gnd(gnd), .vdd(vdd), .A(_880__bF_buf3), .B(_4077_), .C(_4172_), .Y(_4173_) );
NAND3X1 NAND3X1_136 ( .gnd(gnd), .vdd(vdd), .A(_882__bF_buf3), .B(_4076_), .C(_4173_), .Y(_4174_) );
NAND3X1 NAND3X1_137 ( .gnd(gnd), .vdd(vdd), .A(_881_), .B(_4075_), .C(_4174_), .Y(_4175_) );
AOI21X1 AOI21X1_722 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_1_bF_buf2_), .B(micro_hash_ucr_pipe65_bF_buf3), .C(micro_hash_ucr_pipe66_bF_buf3), .Y(_4176_) );
NAND2X1 NAND2X1_513 ( .gnd(gnd), .vdd(vdd), .A(_4176_), .B(_4175_), .Y(_4177_) );
AOI21X1 AOI21X1_723 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe66_bF_buf2), .B(_414__bF_buf1), .C(micro_hash_ucr_pipe67), .Y(_4178_) );
OAI21X1 OAI21X1_1198 ( .gnd(gnd), .vdd(vdd), .A(_1058__bF_buf3), .B(_879__bF_buf2), .C(_878__bF_buf0), .Y(_4179_) );
AOI21X1 AOI21X1_724 ( .gnd(gnd), .vdd(vdd), .A(_4178_), .B(_4177_), .C(_4179_), .Y(_4180_) );
OAI21X1 OAI21X1_1199 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_5_bF_buf3_), .B(_878__bF_buf4), .C(_1949_), .Y(_4181_) );
OAI22X1 OAI22X1_64 ( .gnd(gnd), .vdd(vdd), .A(_1058__bF_buf2), .B(_3093_), .C(_4180_), .D(_4181_), .Y(_298__5_) );
NOR2X1 NOR2X1_705 ( .gnd(gnd), .vdd(vdd), .A(_428__bF_buf1), .B(_884__bF_buf1), .Y(_4182_) );
NAND2X1 NAND2X1_514 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_2_bF_buf3_), .B(micro_hash_ucr_pipe61_bF_buf3), .Y(_4183_) );
NOR2X1 NOR2X1_706 ( .gnd(gnd), .vdd(vdd), .A(_428__bF_buf0), .B(_883__bF_buf2), .Y(_4184_) );
NAND2X1 NAND2X1_515 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_2_bF_buf2_), .B(micro_hash_ucr_pipe59), .Y(_4185_) );
NOR2X1 NOR2X1_707 ( .gnd(gnd), .vdd(vdd), .A(_428__bF_buf3), .B(_888__bF_buf2), .Y(_4186_) );
NAND2X1 NAND2X1_516 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_2_bF_buf1_), .B(micro_hash_ucr_pipe57_bF_buf0), .Y(_4187_) );
NOR2X1 NOR2X1_708 ( .gnd(gnd), .vdd(vdd), .A(_428__bF_buf2), .B(_890__bF_buf3), .Y(_4188_) );
NAND2X1 NAND2X1_517 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_2_bF_buf0_), .B(micro_hash_ucr_pipe55), .Y(_4189_) );
NAND2X1 NAND2X1_518 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_2_bF_buf3_), .B(micro_hash_ucr_pipe51), .Y(_4190_) );
NAND2X1 NAND2X1_519 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_2_bF_buf2_), .B(micro_hash_ucr_pipe45_bF_buf3), .Y(_4191_) );
NOR2X1 NOR2X1_709 ( .gnd(gnd), .vdd(vdd), .A(_428__bF_buf1), .B(_908__bF_buf2), .Y(_4192_) );
NAND2X1 NAND2X1_520 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_2_bF_buf1_), .B(micro_hash_ucr_pipe37), .Y(_4193_) );
NOR2X1 NOR2X1_710 ( .gnd(gnd), .vdd(vdd), .A(_1174_), .B(_910_), .Y(_4194_) );
NAND2X1 NAND2X1_521 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_6_bF_buf2_), .B(micro_hash_ucr_pipe32_bF_buf3), .Y(_4195_) );
NOR2X1 NOR2X1_711 ( .gnd(gnd), .vdd(vdd), .A(_1174_), .B(_915__bF_buf1), .Y(_4196_) );
NAND2X1 NAND2X1_522 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_6_bF_buf1_), .B(micro_hash_ucr_pipe30_bF_buf1), .Y(_4197_) );
NOR2X1 NOR2X1_712 ( .gnd(gnd), .vdd(vdd), .A(_1174_), .B(_917_), .Y(_4198_) );
NAND2X1 NAND2X1_523 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_6_bF_buf0_), .B(micro_hash_ucr_pipe28_bF_buf3), .Y(_4199_) );
NOR2X1 NOR2X1_713 ( .gnd(gnd), .vdd(vdd), .A(_1174_), .B(_916_), .Y(_4200_) );
NAND2X1 NAND2X1_524 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_6_bF_buf3_), .B(micro_hash_ucr_pipe26_bF_buf3), .Y(_4201_) );
NOR2X1 NOR2X1_714 ( .gnd(gnd), .vdd(vdd), .A(_1174_), .B(_921__bF_buf0), .Y(_4202_) );
NAND2X1 NAND2X1_525 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_2_bF_buf0_), .B(micro_hash_ucr_pipe21_bF_buf3), .Y(_4203_) );
NOR2X1 NOR2X1_715 ( .gnd(gnd), .vdd(vdd), .A(_428__bF_buf0), .B(_926__bF_buf0), .Y(_4204_) );
NAND2X1 NAND2X1_526 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_2_bF_buf3_), .B(micro_hash_ucr_pipe19_bF_buf0), .Y(_4205_) );
NOR2X1 NOR2X1_716 ( .gnd(gnd), .vdd(vdd), .A(_428__bF_buf3), .B(_925__bF_buf0), .Y(_4206_) );
NAND2X1 NAND2X1_527 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_2_bF_buf2_), .B(micro_hash_ucr_pipe17_bF_buf1), .Y(_4207_) );
NAND2X1 NAND2X1_528 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_2_bF_buf1_), .B(micro_hash_ucr_pipe13), .Y(_4208_) );
NOR2X1 NOR2X1_717 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe11), .B(_425_), .Y(_4209_) );
NAND3X1 NAND3X1_138 ( .gnd(gnd), .vdd(vdd), .A(_4098_), .B(_4209_), .C(_4096_), .Y(_4210_) );
OAI21X1 OAI21X1_1200 ( .gnd(gnd), .vdd(vdd), .A(_1174_), .B(_968_), .C(_4210_), .Y(_4211_) );
AOI22X1 AOI22X1_39 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_6_bF_buf2_), .B(_957_), .C(_4211_), .D(_931_), .Y(_4212_) );
OAI21X1 OAI21X1_1201 ( .gnd(gnd), .vdd(vdd), .A(_4212_), .B(micro_hash_ucr_pipe13), .C(_4208_), .Y(_4213_) );
NAND2X1 NAND2X1_529 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe14_bF_buf1), .B(_428__bF_buf2), .Y(_4214_) );
OAI21X1 OAI21X1_1202 ( .gnd(gnd), .vdd(vdd), .A(_4213_), .B(micro_hash_ucr_pipe14_bF_buf0), .C(_4214_), .Y(_4215_) );
OAI21X1 OAI21X1_1203 ( .gnd(gnd), .vdd(vdd), .A(_928_), .B(micro_hash_ucr_c_2_bF_buf0_), .C(_930__bF_buf1), .Y(_4216_) );
AOI21X1 AOI21X1_725 ( .gnd(gnd), .vdd(vdd), .A(_928_), .B(_4215_), .C(_4216_), .Y(_4217_) );
NOR2X1 NOR2X1_718 ( .gnd(gnd), .vdd(vdd), .A(_428__bF_buf1), .B(_930__bF_buf0), .Y(_4218_) );
OAI21X1 OAI21X1_1204 ( .gnd(gnd), .vdd(vdd), .A(_4217_), .B(_4218_), .C(_929_), .Y(_4219_) );
AOI21X1 AOI21X1_726 ( .gnd(gnd), .vdd(vdd), .A(_4207_), .B(_4219_), .C(micro_hash_ucr_pipe18_bF_buf1), .Y(_4220_) );
OAI21X1 OAI21X1_1205 ( .gnd(gnd), .vdd(vdd), .A(_4220_), .B(_4206_), .C(_927__bF_buf0), .Y(_4221_) );
AOI21X1 AOI21X1_727 ( .gnd(gnd), .vdd(vdd), .A(_4205_), .B(_4221_), .C(micro_hash_ucr_pipe20_bF_buf1), .Y(_4222_) );
OAI21X1 OAI21X1_1206 ( .gnd(gnd), .vdd(vdd), .A(_4222_), .B(_4204_), .C(_922_), .Y(_4223_) );
AOI21X1 AOI21X1_728 ( .gnd(gnd), .vdd(vdd), .A(_4203_), .B(_4223_), .C(micro_hash_ucr_pipe22_bF_buf0), .Y(_4224_) );
OAI21X1 OAI21X1_1207 ( .gnd(gnd), .vdd(vdd), .A(_428__bF_buf0), .B(_924__bF_buf1), .C(_923_), .Y(_4225_) );
AOI21X1 AOI21X1_729 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe23_bF_buf0), .B(_1174_), .C(micro_hash_ucr_pipe24_bF_buf1), .Y(_4226_) );
OAI21X1 OAI21X1_1208 ( .gnd(gnd), .vdd(vdd), .A(_4224_), .B(_4225_), .C(_4226_), .Y(_4227_) );
NAND2X1 NAND2X1_530 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_6_bF_buf1_), .B(micro_hash_ucr_pipe24_bF_buf0), .Y(_4228_) );
AOI21X1 AOI21X1_730 ( .gnd(gnd), .vdd(vdd), .A(_4228_), .B(_4227_), .C(micro_hash_ucr_pipe25), .Y(_4229_) );
OAI21X1 OAI21X1_1209 ( .gnd(gnd), .vdd(vdd), .A(_4229_), .B(_4202_), .C(_920__bF_buf4), .Y(_4230_) );
AOI21X1 AOI21X1_731 ( .gnd(gnd), .vdd(vdd), .A(_4201_), .B(_4230_), .C(micro_hash_ucr_pipe27), .Y(_4231_) );
OAI21X1 OAI21X1_1210 ( .gnd(gnd), .vdd(vdd), .A(_4231_), .B(_4200_), .C(_918__bF_buf3), .Y(_4232_) );
AOI21X1 AOI21X1_732 ( .gnd(gnd), .vdd(vdd), .A(_4199_), .B(_4232_), .C(micro_hash_ucr_pipe29_bF_buf3), .Y(_4233_) );
OAI21X1 OAI21X1_1211 ( .gnd(gnd), .vdd(vdd), .A(_4233_), .B(_4198_), .C(_913__bF_buf0), .Y(_4234_) );
AOI21X1 AOI21X1_733 ( .gnd(gnd), .vdd(vdd), .A(_4197_), .B(_4234_), .C(micro_hash_ucr_pipe31), .Y(_4235_) );
OAI21X1 OAI21X1_1212 ( .gnd(gnd), .vdd(vdd), .A(_4235_), .B(_4196_), .C(_914__bF_buf0), .Y(_4236_) );
AOI21X1 AOI21X1_734 ( .gnd(gnd), .vdd(vdd), .A(_4195_), .B(_4236_), .C(micro_hash_ucr_pipe33_bF_buf1), .Y(_4237_) );
OAI21X1 OAI21X1_1213 ( .gnd(gnd), .vdd(vdd), .A(_4237_), .B(_4194_), .C(_912__bF_buf1), .Y(_4238_) );
AOI21X1 AOI21X1_735 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_6_bF_buf0_), .B(micro_hash_ucr_pipe34_bF_buf1), .C(micro_hash_ucr_pipe35), .Y(_4239_) );
OAI21X1 OAI21X1_1214 ( .gnd(gnd), .vdd(vdd), .A(_911__bF_buf1), .B(micro_hash_ucr_c_2_bF_buf3_), .C(_907__bF_buf1), .Y(_4240_) );
AOI21X1 AOI21X1_736 ( .gnd(gnd), .vdd(vdd), .A(_4239_), .B(_4238_), .C(_4240_), .Y(_4241_) );
NOR2X1 NOR2X1_719 ( .gnd(gnd), .vdd(vdd), .A(_428__bF_buf3), .B(_907__bF_buf0), .Y(_4242_) );
OAI21X1 OAI21X1_1215 ( .gnd(gnd), .vdd(vdd), .A(_4241_), .B(_4242_), .C(_909__bF_buf1), .Y(_4243_) );
AOI21X1 AOI21X1_737 ( .gnd(gnd), .vdd(vdd), .A(_4193_), .B(_4243_), .C(micro_hash_ucr_pipe38_bF_buf1), .Y(_4244_) );
OAI21X1 OAI21X1_1216 ( .gnd(gnd), .vdd(vdd), .A(_4244_), .B(_4192_), .C(_904__bF_buf2), .Y(_4245_) );
AOI21X1 AOI21X1_738 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_2_bF_buf2_), .B(micro_hash_ucr_pipe39), .C(micro_hash_ucr_pipe40_bF_buf2), .Y(_4246_) );
OAI21X1 OAI21X1_1217 ( .gnd(gnd), .vdd(vdd), .A(_906__bF_buf1), .B(micro_hash_ucr_b_6_bF_buf3_), .C(_905__bF_buf0), .Y(_4247_) );
AOI21X1 AOI21X1_739 ( .gnd(gnd), .vdd(vdd), .A(_4246_), .B(_4245_), .C(_4247_), .Y(_4248_) );
OAI21X1 OAI21X1_1218 ( .gnd(gnd), .vdd(vdd), .A(_1174_), .B(_905__bF_buf3), .C(_901__bF_buf1), .Y(_4249_) );
OAI22X1 OAI22X1_65 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_6_bF_buf2_), .B(_901__bF_buf0), .C(_4248_), .D(_4249_), .Y(_4250_) );
OAI21X1 OAI21X1_1219 ( .gnd(gnd), .vdd(vdd), .A(_903__bF_buf3), .B(micro_hash_ucr_c_2_bF_buf1_), .C(_902__bF_buf4), .Y(_4251_) );
AOI21X1 AOI21X1_740 ( .gnd(gnd), .vdd(vdd), .A(_903__bF_buf2), .B(_4250_), .C(_4251_), .Y(_4252_) );
NOR2X1 NOR2X1_720 ( .gnd(gnd), .vdd(vdd), .A(_428__bF_buf2), .B(_902__bF_buf3), .Y(_4253_) );
OAI21X1 OAI21X1_1220 ( .gnd(gnd), .vdd(vdd), .A(_4252_), .B(_4253_), .C(_898_), .Y(_4254_) );
AOI21X1 AOI21X1_741 ( .gnd(gnd), .vdd(vdd), .A(_4191_), .B(_4254_), .C(micro_hash_ucr_pipe46_bF_buf0), .Y(_4255_) );
OAI21X1 OAI21X1_1221 ( .gnd(gnd), .vdd(vdd), .A(_428__bF_buf1), .B(_900__bF_buf1), .C(_899__bF_buf3), .Y(_4256_) );
OAI22X1 OAI22X1_66 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_2_bF_buf0_), .B(_899__bF_buf2), .C(_4255_), .D(_4256_), .Y(_4257_) );
OAI21X1 OAI21X1_1222 ( .gnd(gnd), .vdd(vdd), .A(_895__bF_buf4), .B(micro_hash_ucr_b_6_bF_buf1_), .C(_897__bF_buf2), .Y(_4258_) );
AOI21X1 AOI21X1_742 ( .gnd(gnd), .vdd(vdd), .A(_895__bF_buf3), .B(_4257_), .C(_4258_), .Y(_4259_) );
OAI21X1 OAI21X1_1223 ( .gnd(gnd), .vdd(vdd), .A(_1174_), .B(_897__bF_buf1), .C(_896__bF_buf0), .Y(_4260_) );
OAI22X1 OAI22X1_67 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_6_bF_buf0_), .B(_896__bF_buf4), .C(_4259_), .D(_4260_), .Y(_4261_) );
OAI21X1 OAI21X1_1224 ( .gnd(gnd), .vdd(vdd), .A(_4261_), .B(micro_hash_ucr_pipe51), .C(_4190_), .Y(_4262_) );
NAND2X1 NAND2X1_531 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe52_bF_buf0), .B(_428__bF_buf0), .Y(_4263_) );
OAI21X1 OAI21X1_1225 ( .gnd(gnd), .vdd(vdd), .A(_4262_), .B(micro_hash_ucr_pipe52_bF_buf4), .C(_4263_), .Y(_4264_) );
OAI21X1 OAI21X1_1226 ( .gnd(gnd), .vdd(vdd), .A(_893_), .B(micro_hash_ucr_c_2_bF_buf3_), .C(_889__bF_buf2), .Y(_4265_) );
AOI21X1 AOI21X1_743 ( .gnd(gnd), .vdd(vdd), .A(_893_), .B(_4264_), .C(_4265_), .Y(_4266_) );
NOR2X1 NOR2X1_721 ( .gnd(gnd), .vdd(vdd), .A(_428__bF_buf3), .B(_889__bF_buf1), .Y(_4267_) );
OAI21X1 OAI21X1_1227 ( .gnd(gnd), .vdd(vdd), .A(_4266_), .B(_4267_), .C(_891_), .Y(_4268_) );
AOI21X1 AOI21X1_744 ( .gnd(gnd), .vdd(vdd), .A(_4189_), .B(_4268_), .C(micro_hash_ucr_pipe56_bF_buf3), .Y(_4269_) );
OAI21X1 OAI21X1_1228 ( .gnd(gnd), .vdd(vdd), .A(_4269_), .B(_4188_), .C(_886_), .Y(_4270_) );
AOI21X1 AOI21X1_745 ( .gnd(gnd), .vdd(vdd), .A(_4187_), .B(_4270_), .C(micro_hash_ucr_pipe58_bF_buf0), .Y(_4271_) );
OAI21X1 OAI21X1_1229 ( .gnd(gnd), .vdd(vdd), .A(_4271_), .B(_4186_), .C(_887__bF_buf3), .Y(_4272_) );
AOI21X1 AOI21X1_746 ( .gnd(gnd), .vdd(vdd), .A(_4185_), .B(_4272_), .C(micro_hash_ucr_pipe60_bF_buf0), .Y(_4273_) );
OAI21X1 OAI21X1_1230 ( .gnd(gnd), .vdd(vdd), .A(_4273_), .B(_4184_), .C(_885_), .Y(_4274_) );
AOI21X1 AOI21X1_747 ( .gnd(gnd), .vdd(vdd), .A(_4183_), .B(_4274_), .C(micro_hash_ucr_pipe62_bF_buf1), .Y(_4275_) );
OAI21X1 OAI21X1_1231 ( .gnd(gnd), .vdd(vdd), .A(_4275_), .B(_4182_), .C(_880__bF_buf2), .Y(_4276_) );
OAI21X1 OAI21X1_1232 ( .gnd(gnd), .vdd(vdd), .A(_1174_), .B(_880__bF_buf1), .C(_4276_), .Y(_4277_) );
NAND2X1 NAND2X1_532 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe64_bF_buf0), .B(_428__bF_buf2), .Y(_4278_) );
OAI21X1 OAI21X1_1233 ( .gnd(gnd), .vdd(vdd), .A(_4277_), .B(micro_hash_ucr_pipe64_bF_buf4), .C(_4278_), .Y(_4279_) );
AOI21X1 AOI21X1_748 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_2_bF_buf2_), .B(micro_hash_ucr_pipe65_bF_buf2), .C(micro_hash_ucr_pipe66_bF_buf1), .Y(_4280_) );
OAI21X1 OAI21X1_1234 ( .gnd(gnd), .vdd(vdd), .A(_4279_), .B(micro_hash_ucr_pipe65_bF_buf1), .C(_4280_), .Y(_4281_) );
AOI21X1 AOI21X1_749 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe66_bF_buf0), .B(_428__bF_buf1), .C(micro_hash_ucr_pipe67), .Y(_4282_) );
OAI21X1 OAI21X1_1235 ( .gnd(gnd), .vdd(vdd), .A(_1174_), .B(_879__bF_buf1), .C(_878__bF_buf3), .Y(_4283_) );
AOI21X1 AOI21X1_750 ( .gnd(gnd), .vdd(vdd), .A(_4282_), .B(_4281_), .C(_4283_), .Y(_4284_) );
OAI21X1 OAI21X1_1236 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_6_bF_buf3_), .B(_878__bF_buf2), .C(_1949_), .Y(_4285_) );
OAI22X1 OAI22X1_68 ( .gnd(gnd), .vdd(vdd), .A(_1174_), .B(_3093_), .C(_4284_), .D(_4285_), .Y(_298__6_) );
NAND2X1 NAND2X1_533 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_3_bF_buf1_), .B(_369_), .Y(_4286_) );
NAND2X1 NAND2X1_534 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe66_bF_buf4), .B(_1721__bF_buf2), .Y(_4287_) );
NAND2X1 NAND2X1_535 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_3_bF_buf0_), .B(micro_hash_ucr_pipe65_bF_buf0), .Y(_4288_) );
NAND2X1 NAND2X1_536 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe64_bF_buf3), .B(_1721__bF_buf1), .Y(_4289_) );
NAND2X1 NAND2X1_537 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_3_bF_buf4_), .B(micro_hash_ucr_pipe63), .Y(_4290_) );
NAND2X1 NAND2X1_538 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe62_bF_buf0), .B(_1721__bF_buf0), .Y(_4291_) );
NAND2X1 NAND2X1_539 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_3_bF_buf3_), .B(micro_hash_ucr_pipe61_bF_buf2), .Y(_4292_) );
NAND2X1 NAND2X1_540 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe60_bF_buf4), .B(_1721__bF_buf4), .Y(_4293_) );
NAND2X1 NAND2X1_541 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_3_bF_buf2_), .B(micro_hash_ucr_pipe59), .Y(_4294_) );
NAND2X1 NAND2X1_542 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe58_bF_buf4), .B(_1721__bF_buf3), .Y(_4295_) );
NAND2X1 NAND2X1_543 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_3_bF_buf1_), .B(micro_hash_ucr_pipe57_bF_buf3), .Y(_4296_) );
NAND2X1 NAND2X1_544 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe56_bF_buf2), .B(_1721__bF_buf2), .Y(_4297_) );
NAND2X1 NAND2X1_545 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_3_bF_buf0_), .B(micro_hash_ucr_pipe55), .Y(_4298_) );
NAND2X1 NAND2X1_546 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe51), .B(_4445_), .Y(_4299_) );
NAND2X1 NAND2X1_547 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe46_bF_buf4), .B(_1721__bF_buf1), .Y(_4300_) );
NAND2X1 NAND2X1_548 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_3_bF_buf4_), .B(micro_hash_ucr_pipe45_bF_buf2), .Y(_4301_) );
NAND2X1 NAND2X1_549 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe44), .B(_1721__bF_buf0), .Y(_4302_) );
NAND2X1 NAND2X1_550 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_3_bF_buf3_), .B(micro_hash_ucr_pipe43), .Y(_4303_) );
NAND2X1 NAND2X1_551 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe42_bF_buf1), .B(_1721__bF_buf4), .Y(_4304_) );
NAND2X1 NAND2X1_552 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_3_bF_buf2_), .B(micro_hash_ucr_pipe41), .Y(_4305_) );
NAND2X1 NAND2X1_553 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe34_bF_buf0), .B(_1721__bF_buf3), .Y(_4306_) );
NAND2X1 NAND2X1_554 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_3_bF_buf1_), .B(micro_hash_ucr_pipe33_bF_buf0), .Y(_4307_) );
NAND2X1 NAND2X1_555 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe32_bF_buf2), .B(_1721__bF_buf2), .Y(_4308_) );
NAND2X1 NAND2X1_556 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_3_bF_buf0_), .B(micro_hash_ucr_pipe31), .Y(_4309_) );
NAND2X1 NAND2X1_557 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe30_bF_buf0), .B(_1721__bF_buf1), .Y(_4310_) );
NAND2X1 NAND2X1_558 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_3_bF_buf4_), .B(micro_hash_ucr_pipe29_bF_buf2), .Y(_4311_) );
NAND2X1 NAND2X1_559 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe28_bF_buf2), .B(_1721__bF_buf0), .Y(_4312_) );
NAND2X1 NAND2X1_560 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_3_bF_buf3_), .B(micro_hash_ucr_pipe27), .Y(_4313_) );
NAND2X1 NAND2X1_561 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe26_bF_buf2), .B(_1721__bF_buf4), .Y(_4314_) );
NAND2X1 NAND2X1_562 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_3_bF_buf2_), .B(micro_hash_ucr_pipe25), .Y(_4315_) );
NAND2X1 NAND2X1_563 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe24_bF_buf4), .B(_1721__bF_buf3), .Y(_4316_) );
NAND2X1 NAND2X1_564 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_3_bF_buf1_), .B(micro_hash_ucr_pipe23_bF_buf3), .Y(_4317_) );
NAND2X1 NAND2X1_565 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe22_bF_buf4), .B(_1721__bF_buf2), .Y(_4318_) );
NAND2X1 NAND2X1_566 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_3_bF_buf0_), .B(micro_hash_ucr_pipe21_bF_buf2), .Y(_4319_) );
NAND2X1 NAND2X1_567 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe20_bF_buf0), .B(_1721__bF_buf1), .Y(_4320_) );
NAND2X1 NAND2X1_568 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_3_bF_buf4_), .B(micro_hash_ucr_pipe19_bF_buf3), .Y(_4321_) );
NAND2X1 NAND2X1_569 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe18_bF_buf0), .B(_1721__bF_buf0), .Y(_4322_) );
NAND2X1 NAND2X1_570 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_3_bF_buf3_), .B(micro_hash_ucr_pipe17_bF_buf0), .Y(_4323_) );
NAND2X1 NAND2X1_571 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe16_bF_buf1), .B(_1721__bF_buf4), .Y(_4324_) );
NAND2X1 NAND2X1_572 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_3_bF_buf2_), .B(micro_hash_ucr_pipe15_bF_buf2), .Y(_4325_) );
NAND2X1 NAND2X1_573 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe14_bF_buf4), .B(_1721__bF_buf3), .Y(_4326_) );
NAND2X1 NAND2X1_574 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_3_bF_buf1_), .B(micro_hash_ucr_pipe13), .Y(_4327_) );
NOR2X1 NOR2X1_722 ( .gnd(gnd), .vdd(vdd), .A(H_15_), .B(micro_hash_ucr_pipe11), .Y(_4328_) );
AND2X2 AND2X2_254 ( .gnd(gnd), .vdd(vdd), .A(_4098_), .B(_4328_), .Y(_4329_) );
NAND2X1 NAND2X1_575 ( .gnd(gnd), .vdd(vdd), .A(_4329_), .B(_4096_), .Y(_4330_) );
OAI21X1 OAI21X1_1237 ( .gnd(gnd), .vdd(vdd), .A(_968_), .B(micro_hash_ucr_c_3_bF_buf0_), .C(_4330_), .Y(_4331_) );
NAND2X1 NAND2X1_576 ( .gnd(gnd), .vdd(vdd), .A(_931_), .B(_4331_), .Y(_4332_) );
AOI21X1 AOI21X1_751 ( .gnd(gnd), .vdd(vdd), .A(_1721__bF_buf2), .B(_957_), .C(micro_hash_ucr_pipe13), .Y(_4333_) );
NAND2X1 NAND2X1_577 ( .gnd(gnd), .vdd(vdd), .A(_4332_), .B(_4333_), .Y(_4334_) );
NAND3X1 NAND3X1_139 ( .gnd(gnd), .vdd(vdd), .A(_932_), .B(_4327_), .C(_4334_), .Y(_4335_) );
NAND3X1 NAND3X1_140 ( .gnd(gnd), .vdd(vdd), .A(_928_), .B(_4326_), .C(_4335_), .Y(_4336_) );
NAND3X1 NAND3X1_141 ( .gnd(gnd), .vdd(vdd), .A(_930__bF_buf4), .B(_4325_), .C(_4336_), .Y(_4337_) );
NAND3X1 NAND3X1_142 ( .gnd(gnd), .vdd(vdd), .A(_929_), .B(_4324_), .C(_4337_), .Y(_4338_) );
NAND3X1 NAND3X1_143 ( .gnd(gnd), .vdd(vdd), .A(_925__bF_buf4), .B(_4323_), .C(_4338_), .Y(_4339_) );
NAND3X1 NAND3X1_144 ( .gnd(gnd), .vdd(vdd), .A(_927__bF_buf3), .B(_4322_), .C(_4339_), .Y(_4340_) );
NAND3X1 NAND3X1_145 ( .gnd(gnd), .vdd(vdd), .A(_926__bF_buf4), .B(_4321_), .C(_4340_), .Y(_4341_) );
NAND3X1 NAND3X1_146 ( .gnd(gnd), .vdd(vdd), .A(_922_), .B(_4320_), .C(_4341_), .Y(_4342_) );
NAND3X1 NAND3X1_147 ( .gnd(gnd), .vdd(vdd), .A(_924__bF_buf0), .B(_4319_), .C(_4342_), .Y(_4343_) );
NAND3X1 NAND3X1_148 ( .gnd(gnd), .vdd(vdd), .A(_923_), .B(_4318_), .C(_4343_), .Y(_4344_) );
NAND3X1 NAND3X1_149 ( .gnd(gnd), .vdd(vdd), .A(_919__bF_buf0), .B(_4317_), .C(_4344_), .Y(_4345_) );
NAND3X1 NAND3X1_150 ( .gnd(gnd), .vdd(vdd), .A(_921__bF_buf3), .B(_4316_), .C(_4345_), .Y(_4346_) );
NAND3X1 NAND3X1_151 ( .gnd(gnd), .vdd(vdd), .A(_920__bF_buf3), .B(_4315_), .C(_4346_), .Y(_4347_) );
NAND3X1 NAND3X1_152 ( .gnd(gnd), .vdd(vdd), .A(_916_), .B(_4314_), .C(_4347_), .Y(_4348_) );
NAND3X1 NAND3X1_153 ( .gnd(gnd), .vdd(vdd), .A(_918__bF_buf2), .B(_4313_), .C(_4348_), .Y(_4349_) );
NAND3X1 NAND3X1_154 ( .gnd(gnd), .vdd(vdd), .A(_917_), .B(_4312_), .C(_4349_), .Y(_4350_) );
NAND3X1 NAND3X1_155 ( .gnd(gnd), .vdd(vdd), .A(_913__bF_buf4), .B(_4311_), .C(_4350_), .Y(_4351_) );
NAND3X1 NAND3X1_156 ( .gnd(gnd), .vdd(vdd), .A(_915__bF_buf0), .B(_4310_), .C(_4351_), .Y(_4352_) );
NAND3X1 NAND3X1_157 ( .gnd(gnd), .vdd(vdd), .A(_914__bF_buf4), .B(_4309_), .C(_4352_), .Y(_4353_) );
NAND3X1 NAND3X1_158 ( .gnd(gnd), .vdd(vdd), .A(_910_), .B(_4308_), .C(_4353_), .Y(_4354_) );
NAND3X1 NAND3X1_159 ( .gnd(gnd), .vdd(vdd), .A(_912__bF_buf0), .B(_4307_), .C(_4354_), .Y(_4355_) );
NAND3X1 NAND3X1_160 ( .gnd(gnd), .vdd(vdd), .A(_911__bF_buf0), .B(_4306_), .C(_4355_), .Y(_4356_) );
AOI21X1 AOI21X1_752 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_3_bF_buf4_), .B(micro_hash_ucr_pipe35), .C(micro_hash_ucr_pipe36_bF_buf0), .Y(_4357_) );
OAI21X1 OAI21X1_1238 ( .gnd(gnd), .vdd(vdd), .A(_907__bF_buf4), .B(micro_hash_ucr_b_7_), .C(_909__bF_buf0), .Y(_4358_) );
AOI21X1 AOI21X1_753 ( .gnd(gnd), .vdd(vdd), .A(_4357_), .B(_4356_), .C(_4358_), .Y(_4359_) );
OAI21X1 OAI21X1_1239 ( .gnd(gnd), .vdd(vdd), .A(_4445_), .B(_909__bF_buf3), .C(_908__bF_buf1), .Y(_4360_) );
NAND2X1 NAND2X1_578 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe38_bF_buf0), .B(_1721__bF_buf1), .Y(_4361_) );
OAI21X1 OAI21X1_1240 ( .gnd(gnd), .vdd(vdd), .A(_4359_), .B(_4360_), .C(_4361_), .Y(_4362_) );
OAI21X1 OAI21X1_1241 ( .gnd(gnd), .vdd(vdd), .A(_904__bF_buf1), .B(micro_hash_ucr_c_3_bF_buf3_), .C(_906__bF_buf0), .Y(_4363_) );
AOI21X1 AOI21X1_754 ( .gnd(gnd), .vdd(vdd), .A(_904__bF_buf0), .B(_4362_), .C(_4363_), .Y(_4364_) );
NOR2X1 NOR2X1_723 ( .gnd(gnd), .vdd(vdd), .A(_1721__bF_buf0), .B(_906__bF_buf4), .Y(_4365_) );
OAI21X1 OAI21X1_1242 ( .gnd(gnd), .vdd(vdd), .A(_4364_), .B(_4365_), .C(_905__bF_buf2), .Y(_4366_) );
NAND3X1 NAND3X1_161 ( .gnd(gnd), .vdd(vdd), .A(_901__bF_buf4), .B(_4305_), .C(_4366_), .Y(_4367_) );
NAND3X1 NAND3X1_162 ( .gnd(gnd), .vdd(vdd), .A(_903__bF_buf1), .B(_4304_), .C(_4367_), .Y(_4368_) );
NAND3X1 NAND3X1_163 ( .gnd(gnd), .vdd(vdd), .A(_902__bF_buf2), .B(_4303_), .C(_4368_), .Y(_4369_) );
NAND3X1 NAND3X1_164 ( .gnd(gnd), .vdd(vdd), .A(_898_), .B(_4302_), .C(_4369_), .Y(_4370_) );
NAND3X1 NAND3X1_165 ( .gnd(gnd), .vdd(vdd), .A(_900__bF_buf0), .B(_4301_), .C(_4370_), .Y(_4371_) );
NAND3X1 NAND3X1_166 ( .gnd(gnd), .vdd(vdd), .A(_899__bF_buf1), .B(_4300_), .C(_4371_), .Y(_4372_) );
AOI21X1 AOI21X1_755 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_3_bF_buf2_), .B(micro_hash_ucr_pipe47), .C(micro_hash_ucr_pipe48_bF_buf2), .Y(_4373_) );
OAI21X1 OAI21X1_1243 ( .gnd(gnd), .vdd(vdd), .A(_895__bF_buf2), .B(micro_hash_ucr_b_7_), .C(_897__bF_buf0), .Y(_4374_) );
AOI21X1 AOI21X1_756 ( .gnd(gnd), .vdd(vdd), .A(_4373_), .B(_4372_), .C(_4374_), .Y(_4375_) );
OAI21X1 OAI21X1_1244 ( .gnd(gnd), .vdd(vdd), .A(_4445_), .B(_897__bF_buf3), .C(_896__bF_buf3), .Y(_4376_) );
NAND2X1 NAND2X1_579 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe50_bF_buf2), .B(_1721__bF_buf4), .Y(_4377_) );
OAI21X1 OAI21X1_1245 ( .gnd(gnd), .vdd(vdd), .A(_4375_), .B(_4376_), .C(_4377_), .Y(_4378_) );
NAND2X1 NAND2X1_580 ( .gnd(gnd), .vdd(vdd), .A(_892_), .B(_4378_), .Y(_4379_) );
NAND3X1 NAND3X1_167 ( .gnd(gnd), .vdd(vdd), .A(_894__bF_buf1), .B(_4299_), .C(_4379_), .Y(_4380_) );
AOI21X1 AOI21X1_757 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_7_), .B(micro_hash_ucr_pipe52_bF_buf3), .C(micro_hash_ucr_pipe53_bF_buf3), .Y(_4381_) );
OAI21X1 OAI21X1_1246 ( .gnd(gnd), .vdd(vdd), .A(_893_), .B(micro_hash_ucr_c_3_bF_buf1_), .C(_889__bF_buf0), .Y(_4382_) );
AOI21X1 AOI21X1_758 ( .gnd(gnd), .vdd(vdd), .A(_4381_), .B(_4380_), .C(_4382_), .Y(_4383_) );
NOR2X1 NOR2X1_724 ( .gnd(gnd), .vdd(vdd), .A(_1721__bF_buf3), .B(_889__bF_buf4), .Y(_4384_) );
OAI21X1 OAI21X1_1247 ( .gnd(gnd), .vdd(vdd), .A(_4383_), .B(_4384_), .C(_891_), .Y(_4385_) );
NAND3X1 NAND3X1_168 ( .gnd(gnd), .vdd(vdd), .A(_890__bF_buf2), .B(_4298_), .C(_4385_), .Y(_4386_) );
NAND3X1 NAND3X1_169 ( .gnd(gnd), .vdd(vdd), .A(_886_), .B(_4297_), .C(_4386_), .Y(_4387_) );
NAND3X1 NAND3X1_170 ( .gnd(gnd), .vdd(vdd), .A(_888__bF_buf1), .B(_4296_), .C(_4387_), .Y(_4388_) );
NAND3X1 NAND3X1_171 ( .gnd(gnd), .vdd(vdd), .A(_887__bF_buf2), .B(_4295_), .C(_4388_), .Y(_4389_) );
NAND3X1 NAND3X1_172 ( .gnd(gnd), .vdd(vdd), .A(_883__bF_buf1), .B(_4294_), .C(_4389_), .Y(_4390_) );
NAND3X1 NAND3X1_173 ( .gnd(gnd), .vdd(vdd), .A(_885_), .B(_4293_), .C(_4390_), .Y(_4391_) );
NAND3X1 NAND3X1_174 ( .gnd(gnd), .vdd(vdd), .A(_884__bF_buf0), .B(_4292_), .C(_4391_), .Y(_4392_) );
NAND3X1 NAND3X1_175 ( .gnd(gnd), .vdd(vdd), .A(_880__bF_buf0), .B(_4291_), .C(_4392_), .Y(_4393_) );
NAND3X1 NAND3X1_176 ( .gnd(gnd), .vdd(vdd), .A(_882__bF_buf2), .B(_4290_), .C(_4393_), .Y(_4394_) );
NAND3X1 NAND3X1_177 ( .gnd(gnd), .vdd(vdd), .A(_881_), .B(_4289_), .C(_4394_), .Y(_4395_) );
NAND3X1 NAND3X1_178 ( .gnd(gnd), .vdd(vdd), .A(_877__bF_buf1), .B(_4288_), .C(_4395_), .Y(_4396_) );
NAND3X1 NAND3X1_179 ( .gnd(gnd), .vdd(vdd), .A(_879__bF_buf0), .B(_4287_), .C(_4396_), .Y(_4397_) );
AOI21X1 AOI21X1_759 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_c_3_bF_buf0_), .B(micro_hash_ucr_pipe67), .C(micro_hash_ucr_pipe68), .Y(_4398_) );
AND2X2 AND2X2_255 ( .gnd(gnd), .vdd(vdd), .A(_4397_), .B(_4398_), .Y(_4399_) );
OAI21X1 OAI21X1_1248 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_b_7_), .B(_878__bF_buf1), .C(_1949_), .Y(_4400_) );
OAI21X1 OAI21X1_1249 ( .gnd(gnd), .vdd(vdd), .A(_4399_), .B(_4400_), .C(_4286_), .Y(_298__7_) );
AOI21X1 AOI21X1_760 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_136_), .B(_587_), .C(micro_hash_ucr_Wx_224_), .Y(_4401_) );
OAI21X1 OAI21X1_1250 ( .gnd(gnd), .vdd(vdd), .A(_587_), .B(micro_hash_ucr_Wx_136_), .C(_4401_), .Y(_4402_) );
AND2X2 AND2X2_256 ( .gnd(gnd), .vdd(vdd), .A(_4402_), .B(_302__bF_buf13), .Y(_296__248_) );
OAI21X1 OAI21X1_1251 ( .gnd(gnd), .vdd(vdd), .A(_590_), .B(micro_hash_ucr_Wx_137_), .C(_2524_), .Y(_4403_) );
AOI21X1 AOI21X1_761 ( .gnd(gnd), .vdd(vdd), .A(_590_), .B(micro_hash_ucr_Wx_137_), .C(_4403_), .Y(_4404_) );
NOR2X1 NOR2X1_725 ( .gnd(gnd), .vdd(vdd), .A(_4404_), .B(_400__bF_buf3), .Y(_296__249_) );
OAI21X1 OAI21X1_1252 ( .gnd(gnd), .vdd(vdd), .A(_593_), .B(micro_hash_ucr_Wx_138_), .C(_2527_), .Y(_4405_) );
AOI21X1 AOI21X1_762 ( .gnd(gnd), .vdd(vdd), .A(_593_), .B(micro_hash_ucr_Wx_138_), .C(_4405_), .Y(_4406_) );
NOR2X1 NOR2X1_726 ( .gnd(gnd), .vdd(vdd), .A(_4406_), .B(_400__bF_buf2), .Y(_296__250_) );
OAI21X1 OAI21X1_1253 ( .gnd(gnd), .vdd(vdd), .A(_596_), .B(micro_hash_ucr_Wx_139_), .C(_2813_), .Y(_4407_) );
AOI21X1 AOI21X1_763 ( .gnd(gnd), .vdd(vdd), .A(_596_), .B(micro_hash_ucr_Wx_139_), .C(_4407_), .Y(_4408_) );
NOR2X1 NOR2X1_727 ( .gnd(gnd), .vdd(vdd), .A(_4408_), .B(_400__bF_buf1), .Y(_296__251_) );
AOI21X1 AOI21X1_764 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_140_), .B(_599_), .C(micro_hash_ucr_Wx_228_), .Y(_4409_) );
OAI21X1 OAI21X1_1254 ( .gnd(gnd), .vdd(vdd), .A(_599_), .B(micro_hash_ucr_Wx_140_), .C(_4409_), .Y(_4410_) );
AND2X2 AND2X2_257 ( .gnd(gnd), .vdd(vdd), .A(_4410_), .B(_302__bF_buf12), .Y(_296__252_) );
AOI21X1 AOI21X1_765 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_141_), .B(_602_), .C(micro_hash_ucr_Wx_229_), .Y(_4411_) );
OAI21X1 OAI21X1_1255 ( .gnd(gnd), .vdd(vdd), .A(_602_), .B(micro_hash_ucr_Wx_141_), .C(_4411_), .Y(_4412_) );
AND2X2 AND2X2_258 ( .gnd(gnd), .vdd(vdd), .A(_4412_), .B(_302__bF_buf11), .Y(_296__253_) );
OAI21X1 OAI21X1_1256 ( .gnd(gnd), .vdd(vdd), .A(_605_), .B(micro_hash_ucr_Wx_142_), .C(_3547_), .Y(_4413_) );
AOI21X1 AOI21X1_766 ( .gnd(gnd), .vdd(vdd), .A(_605_), .B(micro_hash_ucr_Wx_142_), .C(_4413_), .Y(_4414_) );
NOR2X1 NOR2X1_728 ( .gnd(gnd), .vdd(vdd), .A(_4414_), .B(_400__bF_buf0), .Y(_296__254_) );
AOI21X1 AOI21X1_767 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_Wx_143_), .B(_608_), .C(micro_hash_ucr_Wx_231_), .Y(_4415_) );
OAI21X1 OAI21X1_1257 ( .gnd(gnd), .vdd(vdd), .A(_608_), .B(micro_hash_ucr_Wx_143_), .C(_4415_), .Y(_4416_) );
AND2X2 AND2X2_259 ( .gnd(gnd), .vdd(vdd), .A(_4416_), .B(_302__bF_buf10), .Y(_296__255_) );
OAI21X1 OAI21X1_1258 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe70_bF_buf1), .B(comparador_valid_hash), .C(_302__bF_buf9), .Y(_4417_) );
NOR2X1 NOR2X1_729 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_pipe71), .B(_4417_), .Y(_374_) );
DFFPOSX1 DFFPOSX1_391 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_300__0_), .Q(H_0_) );
DFFPOSX1 DFFPOSX1_392 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_300__1_), .Q(H_1_) );
DFFPOSX1 DFFPOSX1_393 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_300__2_), .Q(H_2_) );
DFFPOSX1 DFFPOSX1_394 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_300__3_), .Q(H_3_) );
DFFPOSX1 DFFPOSX1_395 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_300__4_), .Q(H_4_) );
DFFPOSX1 DFFPOSX1_396 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_300__5_), .Q(H_5_) );
DFFPOSX1 DFFPOSX1_397 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_300__6_), .Q(H_6_) );
DFFPOSX1 DFFPOSX1_398 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_300__7_), .Q(H_7_) );
DFFPOSX1 DFFPOSX1_399 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_300__8_), .Q(H_8_) );
DFFPOSX1 DFFPOSX1_400 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_300__9_), .Q(H_9_) );
DFFPOSX1 DFFPOSX1_401 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_300__10_), .Q(H_10_) );
DFFPOSX1 DFFPOSX1_402 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_300__11_), .Q(H_11_) );
DFFPOSX1 DFFPOSX1_403 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_300__12_), .Q(H_12_) );
DFFPOSX1 DFFPOSX1_404 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_300__13_), .Q(H_13_) );
DFFPOSX1 DFFPOSX1_405 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_300__14_), .Q(H_14_) );
DFFPOSX1 DFFPOSX1_406 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_300__15_), .Q(H_15_) );
DFFPOSX1 DFFPOSX1_407 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_300__16_), .Q(H_16_) );
DFFPOSX1 DFFPOSX1_408 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_300__17_), .Q(H_17_) );
DFFPOSX1 DFFPOSX1_409 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_300__18_), .Q(H_18_) );
DFFPOSX1 DFFPOSX1_410 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_300__19_), .Q(H_19_) );
DFFPOSX1 DFFPOSX1_411 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_300__20_), .Q(H_20_) );
DFFPOSX1 DFFPOSX1_412 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_300__21_), .Q(H_21_) );
DFFPOSX1 DFFPOSX1_413 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_300__22_), .Q(H_22_) );
DFFPOSX1 DFFPOSX1_414 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_300__23_), .Q(H_23_) );
DFFPOSX1 DFFPOSX1_415 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_374_), .Q(comparador_valid_hash) );
DFFPOSX1 DFFPOSX1_416 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_298__0_), .Q(micro_hash_ucr_b_0_) );
DFFPOSX1 DFFPOSX1_417 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_298__1_), .Q(micro_hash_ucr_b_1_) );
DFFPOSX1 DFFPOSX1_418 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_298__2_), .Q(micro_hash_ucr_b_2_) );
DFFPOSX1 DFFPOSX1_419 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_298__3_), .Q(micro_hash_ucr_b_3_) );
DFFPOSX1 DFFPOSX1_420 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_298__4_), .Q(micro_hash_ucr_b_4_) );
DFFPOSX1 DFFPOSX1_421 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_298__5_), .Q(micro_hash_ucr_b_5_) );
DFFPOSX1 DFFPOSX1_422 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_298__6_), .Q(micro_hash_ucr_b_6_) );
DFFPOSX1 DFFPOSX1_423 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_298__7_), .Q(micro_hash_ucr_b_7_) );
DFFPOSX1 DFFPOSX1_424 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_299__0_), .Q(micro_hash_ucr_c_0_) );
DFFPOSX1 DFFPOSX1_425 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_299__1_), .Q(micro_hash_ucr_c_1_) );
DFFPOSX1 DFFPOSX1_426 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_299__2_), .Q(micro_hash_ucr_c_2_) );
DFFPOSX1 DFFPOSX1_427 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_299__3_), .Q(micro_hash_ucr_c_3_) );
DFFPOSX1 DFFPOSX1_428 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_299__4_), .Q(micro_hash_ucr_c_4_) );
DFFPOSX1 DFFPOSX1_429 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_299__5_), .Q(micro_hash_ucr_c_5_) );
DFFPOSX1 DFFPOSX1_430 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_299__6_), .Q(micro_hash_ucr_c_6_) );
DFFPOSX1 DFFPOSX1_431 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_299__7_), .Q(micro_hash_ucr_c_7_) );
DFFPOSX1 DFFPOSX1_432 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_375__0_), .Q(micro_hash_ucr_x_0_) );
DFFPOSX1 DFFPOSX1_433 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_375__1_), .Q(micro_hash_ucr_x_1_) );
DFFPOSX1 DFFPOSX1_434 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_375__2_), .Q(micro_hash_ucr_x_2_) );
DFFPOSX1 DFFPOSX1_435 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_375__3_), .Q(micro_hash_ucr_x_3_) );
DFFPOSX1 DFFPOSX1_436 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_375__4_), .Q(micro_hash_ucr_x_4_) );
DFFPOSX1 DFFPOSX1_437 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_375__5_), .Q(micro_hash_ucr_x_5_) );
DFFPOSX1 DFFPOSX1_438 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_375__6_), .Q(micro_hash_ucr_x_6_) );
DFFPOSX1 DFFPOSX1_439 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_375__7_), .Q(micro_hash_ucr_x_7_) );
DFFPOSX1 DFFPOSX1_440 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_301__0_), .Q(micro_hash_ucr_k_0_) );
DFFPOSX1 DFFPOSX1_441 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_301__1_), .Q(micro_hash_ucr_k_1_) );
DFFPOSX1 DFFPOSX1_442 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_301__2_), .Q(micro_hash_ucr_k_2_) );
DFFPOSX1 DFFPOSX1_443 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_301__3_), .Q(micro_hash_ucr_k_3_) );
DFFPOSX1 DFFPOSX1_444 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_301__4_), .Q(micro_hash_ucr_k_4_) );
DFFPOSX1 DFFPOSX1_445 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_301__5_), .Q(micro_hash_ucr_k_5_) );
DFFPOSX1 DFFPOSX1_446 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_301__6_), .Q(micro_hash_ucr_k_6_) );
DFFPOSX1 DFFPOSX1_447 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_301__7_), .Q(micro_hash_ucr_k_7_) );
DFFPOSX1 DFFPOSX1_448 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_297__0_), .Q(micro_hash_ucr_a_0_) );
DFFPOSX1 DFFPOSX1_449 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_297__1_), .Q(micro_hash_ucr_a_1_) );
DFFPOSX1 DFFPOSX1_450 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_297__2_), .Q(micro_hash_ucr_a_2_) );
DFFPOSX1 DFFPOSX1_451 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_297__3_), .Q(micro_hash_ucr_a_3_) );
DFFPOSX1 DFFPOSX1_452 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_297__4_), .Q(micro_hash_ucr_a_4_) );
DFFPOSX1 DFFPOSX1_453 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_297__5_), .Q(micro_hash_ucr_a_5_) );
DFFPOSX1 DFFPOSX1_454 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_297__6_), .Q(micro_hash_ucr_a_6_) );
DFFPOSX1 DFFPOSX1_455 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_297__7_), .Q(micro_hash_ucr_a_7_) );
DFFPOSX1 DFFPOSX1_456 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_302__bF_buf8), .Q(micro_hash_ucr_pipe0) );
DFFPOSX1 DFFPOSX1_457 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_296__0_), .Q(micro_hash_ucr_Wx_0_) );
DFFPOSX1 DFFPOSX1_458 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_296__1_), .Q(micro_hash_ucr_Wx_1_) );
DFFPOSX1 DFFPOSX1_459 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_296__2_), .Q(micro_hash_ucr_Wx_2_) );
DFFPOSX1 DFFPOSX1_460 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_296__3_), .Q(micro_hash_ucr_Wx_3_) );
DFFPOSX1 DFFPOSX1_461 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_296__4_), .Q(micro_hash_ucr_Wx_4_) );
DFFPOSX1 DFFPOSX1_462 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_296__5_), .Q(micro_hash_ucr_Wx_5_) );
DFFPOSX1 DFFPOSX1_463 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_296__6_), .Q(micro_hash_ucr_Wx_6_) );
DFFPOSX1 DFFPOSX1_464 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_296__7_), .Q(micro_hash_ucr_Wx_7_) );
DFFPOSX1 DFFPOSX1_465 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_296__8_), .Q(micro_hash_ucr_Wx_8_) );
DFFPOSX1 DFFPOSX1_466 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_296__9_), .Q(micro_hash_ucr_Wx_9_) );
DFFPOSX1 DFFPOSX1_467 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_296__10_), .Q(micro_hash_ucr_Wx_10_) );
DFFPOSX1 DFFPOSX1_468 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_296__11_), .Q(micro_hash_ucr_Wx_11_) );
DFFPOSX1 DFFPOSX1_469 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_296__12_), .Q(micro_hash_ucr_Wx_12_) );
DFFPOSX1 DFFPOSX1_470 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_296__13_), .Q(micro_hash_ucr_Wx_13_) );
DFFPOSX1 DFFPOSX1_471 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_296__14_), .Q(micro_hash_ucr_Wx_14_) );
DFFPOSX1 DFFPOSX1_472 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_296__15_), .Q(micro_hash_ucr_Wx_15_) );
DFFPOSX1 DFFPOSX1_473 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_296__16_), .Q(micro_hash_ucr_Wx_16_) );
DFFPOSX1 DFFPOSX1_474 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_296__17_), .Q(micro_hash_ucr_Wx_17_) );
DFFPOSX1 DFFPOSX1_475 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf157), .D(_296__18_), .Q(micro_hash_ucr_Wx_18_) );
DFFPOSX1 DFFPOSX1_476 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf156), .D(_296__19_), .Q(micro_hash_ucr_Wx_19_) );
DFFPOSX1 DFFPOSX1_477 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf155), .D(_296__20_), .Q(micro_hash_ucr_Wx_20_) );
DFFPOSX1 DFFPOSX1_478 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf154), .D(_296__21_), .Q(micro_hash_ucr_Wx_21_) );
DFFPOSX1 DFFPOSX1_479 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf153), .D(_296__22_), .Q(micro_hash_ucr_Wx_22_) );
DFFPOSX1 DFFPOSX1_480 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf152), .D(_296__23_), .Q(micro_hash_ucr_Wx_23_) );
DFFPOSX1 DFFPOSX1_481 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf151), .D(_296__24_), .Q(micro_hash_ucr_Wx_24_) );
DFFPOSX1 DFFPOSX1_482 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf150), .D(_296__25_), .Q(micro_hash_ucr_Wx_25_) );
DFFPOSX1 DFFPOSX1_483 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf149), .D(_296__26_), .Q(micro_hash_ucr_Wx_26_) );
DFFPOSX1 DFFPOSX1_484 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf148), .D(_296__27_), .Q(micro_hash_ucr_Wx_27_) );
DFFPOSX1 DFFPOSX1_485 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf147), .D(_296__28_), .Q(micro_hash_ucr_Wx_28_) );
DFFPOSX1 DFFPOSX1_486 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf146), .D(_296__29_), .Q(micro_hash_ucr_Wx_29_) );
DFFPOSX1 DFFPOSX1_487 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf145), .D(_296__30_), .Q(micro_hash_ucr_Wx_30_) );
DFFPOSX1 DFFPOSX1_488 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf144), .D(_296__31_), .Q(micro_hash_ucr_Wx_31_) );
DFFPOSX1 DFFPOSX1_489 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf143), .D(_296__32_), .Q(micro_hash_ucr_Wx_32_) );
DFFPOSX1 DFFPOSX1_490 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf142), .D(_296__33_), .Q(micro_hash_ucr_Wx_33_) );
DFFPOSX1 DFFPOSX1_491 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf141), .D(_296__34_), .Q(micro_hash_ucr_Wx_34_) );
DFFPOSX1 DFFPOSX1_492 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf140), .D(_296__35_), .Q(micro_hash_ucr_Wx_35_) );
DFFPOSX1 DFFPOSX1_493 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf139), .D(_296__36_), .Q(micro_hash_ucr_Wx_36_) );
DFFPOSX1 DFFPOSX1_494 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf138), .D(_296__37_), .Q(micro_hash_ucr_Wx_37_) );
DFFPOSX1 DFFPOSX1_495 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf137), .D(_296__38_), .Q(micro_hash_ucr_Wx_38_) );
DFFPOSX1 DFFPOSX1_496 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf136), .D(_296__39_), .Q(micro_hash_ucr_Wx_39_) );
DFFPOSX1 DFFPOSX1_497 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf135), .D(_296__40_), .Q(micro_hash_ucr_Wx_40_) );
DFFPOSX1 DFFPOSX1_498 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf134), .D(_296__41_), .Q(micro_hash_ucr_Wx_41_) );
DFFPOSX1 DFFPOSX1_499 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf133), .D(_296__42_), .Q(micro_hash_ucr_Wx_42_) );
DFFPOSX1 DFFPOSX1_500 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf132), .D(_296__43_), .Q(micro_hash_ucr_Wx_43_) );
DFFPOSX1 DFFPOSX1_501 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf131), .D(_296__44_), .Q(micro_hash_ucr_Wx_44_) );
DFFPOSX1 DFFPOSX1_502 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf130), .D(_296__45_), .Q(micro_hash_ucr_Wx_45_) );
DFFPOSX1 DFFPOSX1_503 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf129), .D(_296__46_), .Q(micro_hash_ucr_Wx_46_) );
DFFPOSX1 DFFPOSX1_504 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf128), .D(_296__47_), .Q(micro_hash_ucr_Wx_47_) );
DFFPOSX1 DFFPOSX1_505 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf127), .D(_296__48_), .Q(micro_hash_ucr_Wx_48_) );
DFFPOSX1 DFFPOSX1_506 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf126), .D(_296__49_), .Q(micro_hash_ucr_Wx_49_) );
DFFPOSX1 DFFPOSX1_507 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf125), .D(_296__50_), .Q(micro_hash_ucr_Wx_50_) );
DFFPOSX1 DFFPOSX1_508 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf124), .D(_296__51_), .Q(micro_hash_ucr_Wx_51_) );
DFFPOSX1 DFFPOSX1_509 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf123), .D(_296__52_), .Q(micro_hash_ucr_Wx_52_) );
DFFPOSX1 DFFPOSX1_510 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf122), .D(_296__53_), .Q(micro_hash_ucr_Wx_53_) );
DFFPOSX1 DFFPOSX1_511 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf121), .D(_296__54_), .Q(micro_hash_ucr_Wx_54_) );
DFFPOSX1 DFFPOSX1_512 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf120), .D(_296__55_), .Q(micro_hash_ucr_Wx_55_) );
DFFPOSX1 DFFPOSX1_513 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf119), .D(_296__56_), .Q(micro_hash_ucr_Wx_56_) );
DFFPOSX1 DFFPOSX1_514 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf118), .D(_296__57_), .Q(micro_hash_ucr_Wx_57_) );
DFFPOSX1 DFFPOSX1_515 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf117), .D(_296__58_), .Q(micro_hash_ucr_Wx_58_) );
DFFPOSX1 DFFPOSX1_516 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf116), .D(_296__59_), .Q(micro_hash_ucr_Wx_59_) );
DFFPOSX1 DFFPOSX1_517 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf115), .D(_296__60_), .Q(micro_hash_ucr_Wx_60_) );
DFFPOSX1 DFFPOSX1_518 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf114), .D(_296__61_), .Q(micro_hash_ucr_Wx_61_) );
DFFPOSX1 DFFPOSX1_519 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf113), .D(_296__62_), .Q(micro_hash_ucr_Wx_62_) );
DFFPOSX1 DFFPOSX1_520 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf112), .D(_296__63_), .Q(micro_hash_ucr_Wx_63_) );
DFFPOSX1 DFFPOSX1_521 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf111), .D(_296__64_), .Q(micro_hash_ucr_Wx_64_) );
DFFPOSX1 DFFPOSX1_522 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf110), .D(_296__65_), .Q(micro_hash_ucr_Wx_65_) );
DFFPOSX1 DFFPOSX1_523 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf109), .D(_296__66_), .Q(micro_hash_ucr_Wx_66_) );
DFFPOSX1 DFFPOSX1_524 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf108), .D(_296__67_), .Q(micro_hash_ucr_Wx_67_) );
DFFPOSX1 DFFPOSX1_525 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf107), .D(_296__68_), .Q(micro_hash_ucr_Wx_68_) );
DFFPOSX1 DFFPOSX1_526 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(_296__69_), .Q(micro_hash_ucr_Wx_69_) );
DFFPOSX1 DFFPOSX1_527 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(_296__70_), .Q(micro_hash_ucr_Wx_70_) );
DFFPOSX1 DFFPOSX1_528 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(_296__71_), .Q(micro_hash_ucr_Wx_71_) );
DFFPOSX1 DFFPOSX1_529 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(_296__72_), .Q(micro_hash_ucr_Wx_72_) );
DFFPOSX1 DFFPOSX1_530 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(_296__73_), .Q(micro_hash_ucr_Wx_73_) );
DFFPOSX1 DFFPOSX1_531 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(_296__74_), .Q(micro_hash_ucr_Wx_74_) );
DFFPOSX1 DFFPOSX1_532 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(_296__75_), .Q(micro_hash_ucr_Wx_75_) );
DFFPOSX1 DFFPOSX1_533 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(_296__76_), .Q(micro_hash_ucr_Wx_76_) );
DFFPOSX1 DFFPOSX1_534 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_296__77_), .Q(micro_hash_ucr_Wx_77_) );
DFFPOSX1 DFFPOSX1_535 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_296__78_), .Q(micro_hash_ucr_Wx_78_) );
DFFPOSX1 DFFPOSX1_536 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_296__79_), .Q(micro_hash_ucr_Wx_79_) );
DFFPOSX1 DFFPOSX1_537 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_296__80_), .Q(micro_hash_ucr_Wx_80_) );
DFFPOSX1 DFFPOSX1_538 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_296__81_), .Q(micro_hash_ucr_Wx_81_) );
DFFPOSX1 DFFPOSX1_539 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_296__82_), .Q(micro_hash_ucr_Wx_82_) );
DFFPOSX1 DFFPOSX1_540 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_296__83_), .Q(micro_hash_ucr_Wx_83_) );
DFFPOSX1 DFFPOSX1_541 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_296__84_), .Q(micro_hash_ucr_Wx_84_) );
DFFPOSX1 DFFPOSX1_542 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_296__85_), .Q(micro_hash_ucr_Wx_85_) );
DFFPOSX1 DFFPOSX1_543 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_296__86_), .Q(micro_hash_ucr_Wx_86_) );
DFFPOSX1 DFFPOSX1_544 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_296__87_), .Q(micro_hash_ucr_Wx_87_) );
DFFPOSX1 DFFPOSX1_545 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_296__88_), .Q(micro_hash_ucr_Wx_88_) );
DFFPOSX1 DFFPOSX1_546 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_296__89_), .Q(micro_hash_ucr_Wx_89_) );
DFFPOSX1 DFFPOSX1_547 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_296__90_), .Q(micro_hash_ucr_Wx_90_) );
DFFPOSX1 DFFPOSX1_548 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_296__91_), .Q(micro_hash_ucr_Wx_91_) );
DFFPOSX1 DFFPOSX1_549 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_296__92_), .Q(micro_hash_ucr_Wx_92_) );
DFFPOSX1 DFFPOSX1_550 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_296__93_), .Q(micro_hash_ucr_Wx_93_) );
DFFPOSX1 DFFPOSX1_551 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_296__94_), .Q(micro_hash_ucr_Wx_94_) );
DFFPOSX1 DFFPOSX1_552 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_296__95_), .Q(micro_hash_ucr_Wx_95_) );
DFFPOSX1 DFFPOSX1_553 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_296__96_), .Q(micro_hash_ucr_Wx_96_) );
DFFPOSX1 DFFPOSX1_554 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_296__97_), .Q(micro_hash_ucr_Wx_97_) );
DFFPOSX1 DFFPOSX1_555 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_296__98_), .Q(micro_hash_ucr_Wx_98_) );
DFFPOSX1 DFFPOSX1_556 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_296__99_), .Q(micro_hash_ucr_Wx_99_) );
DFFPOSX1 DFFPOSX1_557 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_296__100_), .Q(micro_hash_ucr_Wx_100_) );
DFFPOSX1 DFFPOSX1_558 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_296__101_), .Q(micro_hash_ucr_Wx_101_) );
DFFPOSX1 DFFPOSX1_559 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_296__102_), .Q(micro_hash_ucr_Wx_102_) );
DFFPOSX1 DFFPOSX1_560 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_296__103_), .Q(micro_hash_ucr_Wx_103_) );
DFFPOSX1 DFFPOSX1_561 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_296__104_), .Q(micro_hash_ucr_Wx_104_) );
DFFPOSX1 DFFPOSX1_562 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_296__105_), .Q(micro_hash_ucr_Wx_105_) );
DFFPOSX1 DFFPOSX1_563 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_296__106_), .Q(micro_hash_ucr_Wx_106_) );
DFFPOSX1 DFFPOSX1_564 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_296__107_), .Q(micro_hash_ucr_Wx_107_) );
DFFPOSX1 DFFPOSX1_565 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_296__108_), .Q(micro_hash_ucr_Wx_108_) );
DFFPOSX1 DFFPOSX1_566 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_296__109_), .Q(micro_hash_ucr_Wx_109_) );
DFFPOSX1 DFFPOSX1_567 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_296__110_), .Q(micro_hash_ucr_Wx_110_) );
DFFPOSX1 DFFPOSX1_568 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_296__111_), .Q(micro_hash_ucr_Wx_111_) );
DFFPOSX1 DFFPOSX1_569 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_296__112_), .Q(micro_hash_ucr_Wx_112_) );
DFFPOSX1 DFFPOSX1_570 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_296__113_), .Q(micro_hash_ucr_Wx_113_) );
DFFPOSX1 DFFPOSX1_571 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_296__114_), .Q(micro_hash_ucr_Wx_114_) );
DFFPOSX1 DFFPOSX1_572 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_296__115_), .Q(micro_hash_ucr_Wx_115_) );
DFFPOSX1 DFFPOSX1_573 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_296__116_), .Q(micro_hash_ucr_Wx_116_) );
DFFPOSX1 DFFPOSX1_574 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_296__117_), .Q(micro_hash_ucr_Wx_117_) );
DFFPOSX1 DFFPOSX1_575 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_296__118_), .Q(micro_hash_ucr_Wx_118_) );
DFFPOSX1 DFFPOSX1_576 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_296__119_), .Q(micro_hash_ucr_Wx_119_) );
DFFPOSX1 DFFPOSX1_577 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_296__120_), .Q(micro_hash_ucr_Wx_120_) );
DFFPOSX1 DFFPOSX1_578 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_296__121_), .Q(micro_hash_ucr_Wx_121_) );
DFFPOSX1 DFFPOSX1_579 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_296__122_), .Q(micro_hash_ucr_Wx_122_) );
DFFPOSX1 DFFPOSX1_580 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_296__123_), .Q(micro_hash_ucr_Wx_123_) );
DFFPOSX1 DFFPOSX1_581 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_296__124_), .Q(micro_hash_ucr_Wx_124_) );
DFFPOSX1 DFFPOSX1_582 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_296__125_), .Q(micro_hash_ucr_Wx_125_) );
DFFPOSX1 DFFPOSX1_583 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_296__126_), .Q(micro_hash_ucr_Wx_126_) );
DFFPOSX1 DFFPOSX1_584 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_296__127_), .Q(micro_hash_ucr_Wx_127_) );
DFFPOSX1 DFFPOSX1_585 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_296__128_), .Q(micro_hash_ucr_Wx_128_) );
DFFPOSX1 DFFPOSX1_586 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_296__129_), .Q(micro_hash_ucr_Wx_129_) );
DFFPOSX1 DFFPOSX1_587 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_296__130_), .Q(micro_hash_ucr_Wx_130_) );
DFFPOSX1 DFFPOSX1_588 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_296__131_), .Q(micro_hash_ucr_Wx_131_) );
DFFPOSX1 DFFPOSX1_589 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_296__132_), .Q(micro_hash_ucr_Wx_132_) );
DFFPOSX1 DFFPOSX1_590 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_296__133_), .Q(micro_hash_ucr_Wx_133_) );
DFFPOSX1 DFFPOSX1_591 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_296__134_), .Q(micro_hash_ucr_Wx_134_) );
DFFPOSX1 DFFPOSX1_592 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_296__135_), .Q(micro_hash_ucr_Wx_135_) );
DFFPOSX1 DFFPOSX1_593 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_296__136_), .Q(micro_hash_ucr_Wx_136_) );
DFFPOSX1 DFFPOSX1_594 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_296__137_), .Q(micro_hash_ucr_Wx_137_) );
DFFPOSX1 DFFPOSX1_595 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_296__138_), .Q(micro_hash_ucr_Wx_138_) );
DFFPOSX1 DFFPOSX1_596 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_296__139_), .Q(micro_hash_ucr_Wx_139_) );
DFFPOSX1 DFFPOSX1_597 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_296__140_), .Q(micro_hash_ucr_Wx_140_) );
DFFPOSX1 DFFPOSX1_598 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_296__141_), .Q(micro_hash_ucr_Wx_141_) );
DFFPOSX1 DFFPOSX1_599 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_296__142_), .Q(micro_hash_ucr_Wx_142_) );
DFFPOSX1 DFFPOSX1_600 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_296__143_), .Q(micro_hash_ucr_Wx_143_) );
DFFPOSX1 DFFPOSX1_601 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_296__144_), .Q(micro_hash_ucr_Wx_144_) );
DFFPOSX1 DFFPOSX1_602 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_296__145_), .Q(micro_hash_ucr_Wx_145_) );
DFFPOSX1 DFFPOSX1_603 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_296__146_), .Q(micro_hash_ucr_Wx_146_) );
DFFPOSX1 DFFPOSX1_604 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_296__147_), .Q(micro_hash_ucr_Wx_147_) );
DFFPOSX1 DFFPOSX1_605 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_296__148_), .Q(micro_hash_ucr_Wx_148_) );
DFFPOSX1 DFFPOSX1_606 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_296__149_), .Q(micro_hash_ucr_Wx_149_) );
DFFPOSX1 DFFPOSX1_607 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_296__150_), .Q(micro_hash_ucr_Wx_150_) );
DFFPOSX1 DFFPOSX1_608 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_296__151_), .Q(micro_hash_ucr_Wx_151_) );
DFFPOSX1 DFFPOSX1_609 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_296__152_), .Q(micro_hash_ucr_Wx_152_) );
DFFPOSX1 DFFPOSX1_610 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_296__153_), .Q(micro_hash_ucr_Wx_153_) );
DFFPOSX1 DFFPOSX1_611 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_296__154_), .Q(micro_hash_ucr_Wx_154_) );
DFFPOSX1 DFFPOSX1_612 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_296__155_), .Q(micro_hash_ucr_Wx_155_) );
DFFPOSX1 DFFPOSX1_613 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_296__156_), .Q(micro_hash_ucr_Wx_156_) );
DFFPOSX1 DFFPOSX1_614 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_296__157_), .Q(micro_hash_ucr_Wx_157_) );
DFFPOSX1 DFFPOSX1_615 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_296__158_), .Q(micro_hash_ucr_Wx_158_) );
DFFPOSX1 DFFPOSX1_616 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_296__159_), .Q(micro_hash_ucr_Wx_159_) );
DFFPOSX1 DFFPOSX1_617 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_296__160_), .Q(micro_hash_ucr_Wx_160_) );
DFFPOSX1 DFFPOSX1_618 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_296__161_), .Q(micro_hash_ucr_Wx_161_) );
DFFPOSX1 DFFPOSX1_619 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_296__162_), .Q(micro_hash_ucr_Wx_162_) );
DFFPOSX1 DFFPOSX1_620 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_296__163_), .Q(micro_hash_ucr_Wx_163_) );
DFFPOSX1 DFFPOSX1_621 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_296__164_), .Q(micro_hash_ucr_Wx_164_) );
DFFPOSX1 DFFPOSX1_622 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_296__165_), .Q(micro_hash_ucr_Wx_165_) );
DFFPOSX1 DFFPOSX1_623 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_296__166_), .Q(micro_hash_ucr_Wx_166_) );
DFFPOSX1 DFFPOSX1_624 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_296__167_), .Q(micro_hash_ucr_Wx_167_) );
DFFPOSX1 DFFPOSX1_625 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_296__168_), .Q(micro_hash_ucr_Wx_168_) );
DFFPOSX1 DFFPOSX1_626 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_296__169_), .Q(micro_hash_ucr_Wx_169_) );
DFFPOSX1 DFFPOSX1_627 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_296__170_), .Q(micro_hash_ucr_Wx_170_) );
DFFPOSX1 DFFPOSX1_628 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_296__171_), .Q(micro_hash_ucr_Wx_171_) );
DFFPOSX1 DFFPOSX1_629 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_296__172_), .Q(micro_hash_ucr_Wx_172_) );
DFFPOSX1 DFFPOSX1_630 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_296__173_), .Q(micro_hash_ucr_Wx_173_) );
DFFPOSX1 DFFPOSX1_631 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_296__174_), .Q(micro_hash_ucr_Wx_174_) );
DFFPOSX1 DFFPOSX1_632 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_296__175_), .Q(micro_hash_ucr_Wx_175_) );
DFFPOSX1 DFFPOSX1_633 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf157), .D(_296__176_), .Q(micro_hash_ucr_Wx_176_) );
DFFPOSX1 DFFPOSX1_634 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf156), .D(_296__177_), .Q(micro_hash_ucr_Wx_177_) );
DFFPOSX1 DFFPOSX1_635 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf155), .D(_296__178_), .Q(micro_hash_ucr_Wx_178_) );
DFFPOSX1 DFFPOSX1_636 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf154), .D(_296__179_), .Q(micro_hash_ucr_Wx_179_) );
DFFPOSX1 DFFPOSX1_637 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf153), .D(_296__180_), .Q(micro_hash_ucr_Wx_180_) );
DFFPOSX1 DFFPOSX1_638 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf152), .D(_296__181_), .Q(micro_hash_ucr_Wx_181_) );
DFFPOSX1 DFFPOSX1_639 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf151), .D(_296__182_), .Q(micro_hash_ucr_Wx_182_) );
DFFPOSX1 DFFPOSX1_640 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf150), .D(_296__183_), .Q(micro_hash_ucr_Wx_183_) );
DFFPOSX1 DFFPOSX1_641 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf149), .D(_296__184_), .Q(micro_hash_ucr_Wx_184_) );
DFFPOSX1 DFFPOSX1_642 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf148), .D(_296__185_), .Q(micro_hash_ucr_Wx_185_) );
DFFPOSX1 DFFPOSX1_643 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf147), .D(_296__186_), .Q(micro_hash_ucr_Wx_186_) );
DFFPOSX1 DFFPOSX1_644 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf146), .D(_296__187_), .Q(micro_hash_ucr_Wx_187_) );
DFFPOSX1 DFFPOSX1_645 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf145), .D(_296__188_), .Q(micro_hash_ucr_Wx_188_) );
DFFPOSX1 DFFPOSX1_646 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf144), .D(_296__189_), .Q(micro_hash_ucr_Wx_189_) );
DFFPOSX1 DFFPOSX1_647 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf143), .D(_296__190_), .Q(micro_hash_ucr_Wx_190_) );
DFFPOSX1 DFFPOSX1_648 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf142), .D(_296__191_), .Q(micro_hash_ucr_Wx_191_) );
DFFPOSX1 DFFPOSX1_649 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf141), .D(_296__192_), .Q(micro_hash_ucr_Wx_192_) );
DFFPOSX1 DFFPOSX1_650 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf140), .D(_296__193_), .Q(micro_hash_ucr_Wx_193_) );
DFFPOSX1 DFFPOSX1_651 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf139), .D(_296__194_), .Q(micro_hash_ucr_Wx_194_) );
DFFPOSX1 DFFPOSX1_652 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf138), .D(_296__195_), .Q(micro_hash_ucr_Wx_195_) );
DFFPOSX1 DFFPOSX1_653 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf137), .D(_296__196_), .Q(micro_hash_ucr_Wx_196_) );
DFFPOSX1 DFFPOSX1_654 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf136), .D(_296__197_), .Q(micro_hash_ucr_Wx_197_) );
DFFPOSX1 DFFPOSX1_655 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf135), .D(_296__198_), .Q(micro_hash_ucr_Wx_198_) );
DFFPOSX1 DFFPOSX1_656 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf134), .D(_296__199_), .Q(micro_hash_ucr_Wx_199_) );
DFFPOSX1 DFFPOSX1_657 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf133), .D(_296__200_), .Q(micro_hash_ucr_Wx_200_) );
DFFPOSX1 DFFPOSX1_658 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf132), .D(_296__201_), .Q(micro_hash_ucr_Wx_201_) );
DFFPOSX1 DFFPOSX1_659 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf131), .D(_296__202_), .Q(micro_hash_ucr_Wx_202_) );
DFFPOSX1 DFFPOSX1_660 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf130), .D(_296__203_), .Q(micro_hash_ucr_Wx_203_) );
DFFPOSX1 DFFPOSX1_661 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf129), .D(_296__204_), .Q(micro_hash_ucr_Wx_204_) );
DFFPOSX1 DFFPOSX1_662 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf128), .D(_296__205_), .Q(micro_hash_ucr_Wx_205_) );
DFFPOSX1 DFFPOSX1_663 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf127), .D(_296__206_), .Q(micro_hash_ucr_Wx_206_) );
DFFPOSX1 DFFPOSX1_664 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf126), .D(_296__207_), .Q(micro_hash_ucr_Wx_207_) );
DFFPOSX1 DFFPOSX1_665 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf125), .D(_296__208_), .Q(micro_hash_ucr_Wx_208_) );
DFFPOSX1 DFFPOSX1_666 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf124), .D(_296__209_), .Q(micro_hash_ucr_Wx_209_) );
DFFPOSX1 DFFPOSX1_667 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf123), .D(_296__210_), .Q(micro_hash_ucr_Wx_210_) );
DFFPOSX1 DFFPOSX1_668 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf122), .D(_296__211_), .Q(micro_hash_ucr_Wx_211_) );
DFFPOSX1 DFFPOSX1_669 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf121), .D(_296__212_), .Q(micro_hash_ucr_Wx_212_) );
DFFPOSX1 DFFPOSX1_670 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf120), .D(_296__213_), .Q(micro_hash_ucr_Wx_213_) );
DFFPOSX1 DFFPOSX1_671 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf119), .D(_296__214_), .Q(micro_hash_ucr_Wx_214_) );
DFFPOSX1 DFFPOSX1_672 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf118), .D(_296__215_), .Q(micro_hash_ucr_Wx_215_) );
DFFPOSX1 DFFPOSX1_673 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf117), .D(_296__216_), .Q(micro_hash_ucr_Wx_216_) );
DFFPOSX1 DFFPOSX1_674 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf116), .D(_296__217_), .Q(micro_hash_ucr_Wx_217_) );
DFFPOSX1 DFFPOSX1_675 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf115), .D(_296__218_), .Q(micro_hash_ucr_Wx_218_) );
DFFPOSX1 DFFPOSX1_676 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf114), .D(_296__219_), .Q(micro_hash_ucr_Wx_219_) );
DFFPOSX1 DFFPOSX1_677 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf113), .D(_296__220_), .Q(micro_hash_ucr_Wx_220_) );
DFFPOSX1 DFFPOSX1_678 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf112), .D(_296__221_), .Q(micro_hash_ucr_Wx_221_) );
DFFPOSX1 DFFPOSX1_679 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf111), .D(_296__222_), .Q(micro_hash_ucr_Wx_222_) );
DFFPOSX1 DFFPOSX1_680 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf110), .D(_296__223_), .Q(micro_hash_ucr_Wx_223_) );
DFFPOSX1 DFFPOSX1_681 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf109), .D(_296__224_), .Q(micro_hash_ucr_Wx_224_) );
DFFPOSX1 DFFPOSX1_682 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf108), .D(_296__225_), .Q(micro_hash_ucr_Wx_225_) );
DFFPOSX1 DFFPOSX1_683 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf107), .D(_296__226_), .Q(micro_hash_ucr_Wx_226_) );
DFFPOSX1 DFFPOSX1_684 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(_296__227_), .Q(micro_hash_ucr_Wx_227_) );
DFFPOSX1 DFFPOSX1_685 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(_296__228_), .Q(micro_hash_ucr_Wx_228_) );
DFFPOSX1 DFFPOSX1_686 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(_296__229_), .Q(micro_hash_ucr_Wx_229_) );
DFFPOSX1 DFFPOSX1_687 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(_296__230_), .Q(micro_hash_ucr_Wx_230_) );
DFFPOSX1 DFFPOSX1_688 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(_296__231_), .Q(micro_hash_ucr_Wx_231_) );
DFFPOSX1 DFFPOSX1_689 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(_296__232_), .Q(micro_hash_ucr_Wx_232_) );
DFFPOSX1 DFFPOSX1_690 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(_296__233_), .Q(micro_hash_ucr_Wx_233_) );
DFFPOSX1 DFFPOSX1_691 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(_296__234_), .Q(micro_hash_ucr_Wx_234_) );
DFFPOSX1 DFFPOSX1_692 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_296__235_), .Q(micro_hash_ucr_Wx_235_) );
DFFPOSX1 DFFPOSX1_693 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_296__236_), .Q(micro_hash_ucr_Wx_236_) );
DFFPOSX1 DFFPOSX1_694 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_296__237_), .Q(micro_hash_ucr_Wx_237_) );
DFFPOSX1 DFFPOSX1_695 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_296__238_), .Q(micro_hash_ucr_Wx_238_) );
DFFPOSX1 DFFPOSX1_696 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_296__239_), .Q(micro_hash_ucr_Wx_239_) );
DFFPOSX1 DFFPOSX1_697 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_296__240_), .Q(micro_hash_ucr_Wx_240_) );
DFFPOSX1 DFFPOSX1_698 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_296__241_), .Q(micro_hash_ucr_Wx_241_) );
DFFPOSX1 DFFPOSX1_699 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_296__242_), .Q(micro_hash_ucr_Wx_242_) );
DFFPOSX1 DFFPOSX1_700 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_296__243_), .Q(micro_hash_ucr_Wx_243_) );
DFFPOSX1 DFFPOSX1_701 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_296__244_), .Q(micro_hash_ucr_Wx_244_) );
DFFPOSX1 DFFPOSX1_702 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_296__245_), .Q(micro_hash_ucr_Wx_245_) );
DFFPOSX1 DFFPOSX1_703 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_296__246_), .Q(micro_hash_ucr_Wx_246_) );
DFFPOSX1 DFFPOSX1_704 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_296__247_), .Q(micro_hash_ucr_Wx_247_) );
DFFPOSX1 DFFPOSX1_705 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_296__248_), .Q(micro_hash_ucr_Wx_248_) );
DFFPOSX1 DFFPOSX1_706 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_296__249_), .Q(micro_hash_ucr_Wx_249_) );
DFFPOSX1 DFFPOSX1_707 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_296__250_), .Q(micro_hash_ucr_Wx_250_) );
DFFPOSX1 DFFPOSX1_708 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_296__251_), .Q(micro_hash_ucr_Wx_251_) );
DFFPOSX1 DFFPOSX1_709 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_296__252_), .Q(micro_hash_ucr_Wx_252_) );
DFFPOSX1 DFFPOSX1_710 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_296__253_), .Q(micro_hash_ucr_Wx_253_) );
DFFPOSX1 DFFPOSX1_711 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_296__254_), .Q(micro_hash_ucr_Wx_254_) );
DFFPOSX1 DFFPOSX1_712 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_296__255_), .Q(micro_hash_ucr_Wx_255_) );
DFFPOSX1 DFFPOSX1_713 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_313_), .Q(micro_hash_ucr_pipe1) );
DFFPOSX1 DFFPOSX1_714 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_324_), .Q(micro_hash_ucr_pipe2) );
DFFPOSX1 DFFPOSX1_715 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_335_), .Q(micro_hash_ucr_pipe3) );
DFFPOSX1 DFFPOSX1_716 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_346_), .Q(micro_hash_ucr_pipe4) );
DFFPOSX1 DFFPOSX1_717 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_357_), .Q(micro_hash_ucr_pipe5) );
DFFPOSX1 DFFPOSX1_718 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_368_), .Q(micro_hash_ucr_pipe6) );
DFFPOSX1 DFFPOSX1_719 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_371_), .Q(micro_hash_ucr_pipe7) );
DFFPOSX1 DFFPOSX1_720 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_372_), .Q(micro_hash_ucr_pipe8) );
DFFPOSX1 DFFPOSX1_721 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_373_), .Q(micro_hash_ucr_pipe9) );
DFFPOSX1 DFFPOSX1_722 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_303_), .Q(micro_hash_ucr_pipe10) );
DFFPOSX1 DFFPOSX1_723 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_304_), .Q(micro_hash_ucr_pipe11) );
DFFPOSX1 DFFPOSX1_724 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_305_), .Q(micro_hash_ucr_pipe12) );
DFFPOSX1 DFFPOSX1_725 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_306_), .Q(micro_hash_ucr_pipe13) );
DFFPOSX1 DFFPOSX1_726 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_307_), .Q(micro_hash_ucr_pipe14) );
DFFPOSX1 DFFPOSX1_727 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_308_), .Q(micro_hash_ucr_pipe15) );
DFFPOSX1 DFFPOSX1_728 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_309_), .Q(micro_hash_ucr_pipe16) );
DFFPOSX1 DFFPOSX1_729 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_310_), .Q(micro_hash_ucr_pipe17) );
DFFPOSX1 DFFPOSX1_730 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_311_), .Q(micro_hash_ucr_pipe18) );
DFFPOSX1 DFFPOSX1_731 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_312_), .Q(micro_hash_ucr_pipe19) );
DFFPOSX1 DFFPOSX1_732 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_314_), .Q(micro_hash_ucr_pipe20) );
DFFPOSX1 DFFPOSX1_733 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_315_), .Q(micro_hash_ucr_pipe21) );
DFFPOSX1 DFFPOSX1_734 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_316_), .Q(micro_hash_ucr_pipe22) );
DFFPOSX1 DFFPOSX1_735 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_317_), .Q(micro_hash_ucr_pipe23) );
DFFPOSX1 DFFPOSX1_736 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_318_), .Q(micro_hash_ucr_pipe24) );
DFFPOSX1 DFFPOSX1_737 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_319_), .Q(micro_hash_ucr_pipe25) );
DFFPOSX1 DFFPOSX1_738 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_320_), .Q(micro_hash_ucr_pipe26) );
DFFPOSX1 DFFPOSX1_739 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_321_), .Q(micro_hash_ucr_pipe27) );
DFFPOSX1 DFFPOSX1_740 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_322_), .Q(micro_hash_ucr_pipe28) );
DFFPOSX1 DFFPOSX1_741 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_323_), .Q(micro_hash_ucr_pipe29) );
DFFPOSX1 DFFPOSX1_742 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_325_), .Q(micro_hash_ucr_pipe30) );
DFFPOSX1 DFFPOSX1_743 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_326_), .Q(micro_hash_ucr_pipe31) );
DFFPOSX1 DFFPOSX1_744 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_327_), .Q(micro_hash_ucr_pipe32) );
DFFPOSX1 DFFPOSX1_745 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_328_), .Q(micro_hash_ucr_pipe33) );
DFFPOSX1 DFFPOSX1_746 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_329_), .Q(micro_hash_ucr_pipe34) );
DFFPOSX1 DFFPOSX1_747 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_330_), .Q(micro_hash_ucr_pipe35) );
DFFPOSX1 DFFPOSX1_748 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_331_), .Q(micro_hash_ucr_pipe36) );
DFFPOSX1 DFFPOSX1_749 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_332_), .Q(micro_hash_ucr_pipe37) );
DFFPOSX1 DFFPOSX1_750 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_333_), .Q(micro_hash_ucr_pipe38) );
DFFPOSX1 DFFPOSX1_751 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_334_), .Q(micro_hash_ucr_pipe39) );
DFFPOSX1 DFFPOSX1_752 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_336_), .Q(micro_hash_ucr_pipe40) );
DFFPOSX1 DFFPOSX1_753 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_337_), .Q(micro_hash_ucr_pipe41) );
DFFPOSX1 DFFPOSX1_754 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_338_), .Q(micro_hash_ucr_pipe42) );
DFFPOSX1 DFFPOSX1_755 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_339_), .Q(micro_hash_ucr_pipe43) );
DFFPOSX1 DFFPOSX1_756 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_340_), .Q(micro_hash_ucr_pipe44) );
DFFPOSX1 DFFPOSX1_757 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_341_), .Q(micro_hash_ucr_pipe45) );
DFFPOSX1 DFFPOSX1_758 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_342_), .Q(micro_hash_ucr_pipe46) );
DFFPOSX1 DFFPOSX1_759 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_343_), .Q(micro_hash_ucr_pipe47) );
DFFPOSX1 DFFPOSX1_760 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_344_), .Q(micro_hash_ucr_pipe48) );
DFFPOSX1 DFFPOSX1_761 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_345_), .Q(micro_hash_ucr_pipe49) );
DFFPOSX1 DFFPOSX1_762 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_347_), .Q(micro_hash_ucr_pipe50) );
DFFPOSX1 DFFPOSX1_763 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_348_), .Q(micro_hash_ucr_pipe51) );
DFFPOSX1 DFFPOSX1_764 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_349_), .Q(micro_hash_ucr_pipe52) );
DFFPOSX1 DFFPOSX1_765 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_350_), .Q(micro_hash_ucr_pipe53) );
DFFPOSX1 DFFPOSX1_766 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_351_), .Q(micro_hash_ucr_pipe54) );
DFFPOSX1 DFFPOSX1_767 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_352_), .Q(micro_hash_ucr_pipe55) );
DFFPOSX1 DFFPOSX1_768 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_353_), .Q(micro_hash_ucr_pipe56) );
DFFPOSX1 DFFPOSX1_769 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_354_), .Q(micro_hash_ucr_pipe57) );
DFFPOSX1 DFFPOSX1_770 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_355_), .Q(micro_hash_ucr_pipe58) );
DFFPOSX1 DFFPOSX1_771 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_356_), .Q(micro_hash_ucr_pipe59) );
DFFPOSX1 DFFPOSX1_772 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_358_), .Q(micro_hash_ucr_pipe60) );
DFFPOSX1 DFFPOSX1_773 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_359_), .Q(micro_hash_ucr_pipe61) );
DFFPOSX1 DFFPOSX1_774 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_360_), .Q(micro_hash_ucr_pipe62) );
DFFPOSX1 DFFPOSX1_775 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_361_), .Q(micro_hash_ucr_pipe63) );
DFFPOSX1 DFFPOSX1_776 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_362_), .Q(micro_hash_ucr_pipe64) );
DFFPOSX1 DFFPOSX1_777 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_363_), .Q(micro_hash_ucr_pipe65) );
DFFPOSX1 DFFPOSX1_778 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_364_), .Q(micro_hash_ucr_pipe66) );
DFFPOSX1 DFFPOSX1_779 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_365_), .Q(micro_hash_ucr_pipe67) );
DFFPOSX1 DFFPOSX1_780 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_366_), .Q(micro_hash_ucr_pipe68) );
DFFPOSX1 DFFPOSX1_781 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_367_), .Q(micro_hash_ucr_pipe69) );
DFFPOSX1 DFFPOSX1_782 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_369_), .Q(micro_hash_ucr_pipe70) );
DFFPOSX1 DFFPOSX1_783 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_370_), .Q(micro_hash_ucr_pipe71) );
INVX1 INVX1_316 ( .gnd(gnd), .vdd(vdd), .A(_0__bF_buf7), .Y(_8627_) );
NAND2X1 NAND2X1_581 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf6), .B(_8627_), .Y(_8628_) );
NOR2X1 NOR2X1_730 ( .gnd(gnd), .vdd(vdd), .A(comparador_next_bF_buf2), .B(_8628_), .Y(_4496_) );
NOR2X1 NOR2X1_731 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe70_bF_buf3), .B(micro_hash_ucr_2_pipe5), .Y(_8629_) );
NAND2X1 NAND2X1_582 ( .gnd(gnd), .vdd(vdd), .A(H_2_16_), .B(_8629_), .Y(_8630_) );
INVX1 INVX1_317 ( .gnd(gnd), .vdd(vdd), .A(H_2_16_), .Y(_8631_) );
INVX8 INVX8_96 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_0_bF_buf3_), .Y(_8632_) );
OAI21X1 OAI21X1_1259 ( .gnd(gnd), .vdd(vdd), .A(_8631_), .B(_8632__bF_buf3), .C(micro_hash_ucr_2_pipe70_bF_buf2), .Y(_8633_) );
OAI21X1 OAI21X1_1260 ( .gnd(gnd), .vdd(vdd), .A(H_2_16_), .B(micro_hash_ucr_2_c_0_bF_buf2_), .C(_4496__bF_buf13), .Y(_8634_) );
AOI21X1 AOI21X1_768 ( .gnd(gnd), .vdd(vdd), .A(_8630_), .B(_8633_), .C(_8634_), .Y(_4494__16_) );
NOR2X1 NOR2X1_732 ( .gnd(gnd), .vdd(vdd), .A(_8631_), .B(_8632__bF_buf2), .Y(_8635_) );
NOR2X1 NOR2X1_733 ( .gnd(gnd), .vdd(vdd), .A(H_2_17_), .B(micro_hash_ucr_2_c_1_bF_buf3_), .Y(_8636_) );
NAND2X1 NAND2X1_583 ( .gnd(gnd), .vdd(vdd), .A(H_2_17_), .B(micro_hash_ucr_2_c_1_bF_buf2_), .Y(_8637_) );
INVX1 INVX1_318 ( .gnd(gnd), .vdd(vdd), .A(_8637_), .Y(_8638_) );
NOR2X1 NOR2X1_734 ( .gnd(gnd), .vdd(vdd), .A(_8636_), .B(_8638_), .Y(_8639_) );
XNOR2X1 XNOR2X1_195 ( .gnd(gnd), .vdd(vdd), .A(_8639_), .B(_8635_), .Y(_8640_) );
INVX8 INVX8_97 ( .gnd(gnd), .vdd(vdd), .A(_8629_), .Y(_8641_) );
OAI21X1 OAI21X1_1261 ( .gnd(gnd), .vdd(vdd), .A(H_2_17_), .B(_8641_), .C(_4496__bF_buf12), .Y(_8642_) );
AOI21X1 AOI21X1_769 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe70_bF_buf1), .B(_8640_), .C(_8642_), .Y(_4494__17_) );
INVX1 INVX1_319 ( .gnd(gnd), .vdd(vdd), .A(_8635_), .Y(_8643_) );
OAI21X1 OAI21X1_1262 ( .gnd(gnd), .vdd(vdd), .A(_8643_), .B(_8636_), .C(_8637_), .Y(_8644_) );
XOR2X1 XOR2X1_77 ( .gnd(gnd), .vdd(vdd), .A(H_2_18_), .B(micro_hash_ucr_2_c_2_bF_buf3_), .Y(_8645_) );
XNOR2X1 XNOR2X1_196 ( .gnd(gnd), .vdd(vdd), .A(_8644_), .B(_8645_), .Y(_8646_) );
OAI21X1 OAI21X1_1263 ( .gnd(gnd), .vdd(vdd), .A(H_2_18_), .B(_8641_), .C(_4496__bF_buf11), .Y(_8647_) );
AOI21X1 AOI21X1_770 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe70_bF_buf0), .B(_8646_), .C(_8647_), .Y(_4494__18_) );
INVX1 INVX1_320 ( .gnd(gnd), .vdd(vdd), .A(_8644_), .Y(_8648_) );
INVX1 INVX1_321 ( .gnd(gnd), .vdd(vdd), .A(_8645_), .Y(_8649_) );
NOR2X1 NOR2X1_735 ( .gnd(gnd), .vdd(vdd), .A(_8649_), .B(_8648_), .Y(_8650_) );
AOI21X1 AOI21X1_771 ( .gnd(gnd), .vdd(vdd), .A(H_2_18_), .B(micro_hash_ucr_2_c_2_bF_buf2_), .C(_8650_), .Y(_8651_) );
NOR2X1 NOR2X1_736 ( .gnd(gnd), .vdd(vdd), .A(H_2_19_), .B(micro_hash_ucr_2_c_3_bF_buf3_), .Y(_8652_) );
INVX1 INVX1_322 ( .gnd(gnd), .vdd(vdd), .A(H_2_19_), .Y(_8653_) );
INVX8 INVX8_98 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_3_bF_buf2_), .Y(_8654_) );
NOR2X1 NOR2X1_737 ( .gnd(gnd), .vdd(vdd), .A(_8653_), .B(_8654_), .Y(_8655_) );
OR2X2 OR2X2_44 ( .gnd(gnd), .vdd(vdd), .A(_8655_), .B(_8652_), .Y(_8656_) );
XNOR2X1 XNOR2X1_197 ( .gnd(gnd), .vdd(vdd), .A(_8651_), .B(_8656_), .Y(_8657_) );
OAI21X1 OAI21X1_1264 ( .gnd(gnd), .vdd(vdd), .A(H_2_19_), .B(_8641_), .C(_4496__bF_buf10), .Y(_8658_) );
AOI21X1 AOI21X1_772 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe70_bF_buf3), .B(_8657_), .C(_8658_), .Y(_4494__19_) );
NOR2X1 NOR2X1_738 ( .gnd(gnd), .vdd(vdd), .A(H_2_20_), .B(micro_hash_ucr_2_c_4_), .Y(_8659_) );
AND2X2 AND2X2_260 ( .gnd(gnd), .vdd(vdd), .A(H_2_20_), .B(micro_hash_ucr_2_c_4_), .Y(_8660_) );
NOR2X1 NOR2X1_739 ( .gnd(gnd), .vdd(vdd), .A(_8659_), .B(_8660_), .Y(_8661_) );
INVX1 INVX1_323 ( .gnd(gnd), .vdd(vdd), .A(_8655_), .Y(_8662_) );
OAI21X1 OAI21X1_1265 ( .gnd(gnd), .vdd(vdd), .A(_8651_), .B(_8652_), .C(_8662_), .Y(_8663_) );
XNOR2X1 XNOR2X1_198 ( .gnd(gnd), .vdd(vdd), .A(_8663_), .B(_8661_), .Y(_8664_) );
OAI21X1 OAI21X1_1266 ( .gnd(gnd), .vdd(vdd), .A(H_2_20_), .B(_8641_), .C(_4496__bF_buf9), .Y(_8665_) );
AOI21X1 AOI21X1_773 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe70_bF_buf2), .B(_8664_), .C(_8665_), .Y(_4494__20_) );
AOI21X1 AOI21X1_774 ( .gnd(gnd), .vdd(vdd), .A(_8661_), .B(_8663_), .C(_8660_), .Y(_8666_) );
NOR2X1 NOR2X1_740 ( .gnd(gnd), .vdd(vdd), .A(H_2_21_), .B(micro_hash_ucr_2_c_5_), .Y(_8667_) );
INVX1 INVX1_324 ( .gnd(gnd), .vdd(vdd), .A(H_2_21_), .Y(_8668_) );
INVX1 INVX1_325 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_5_), .Y(_8669_) );
NOR2X1 NOR2X1_741 ( .gnd(gnd), .vdd(vdd), .A(_8668_), .B(_8669_), .Y(_8670_) );
NOR2X1 NOR2X1_742 ( .gnd(gnd), .vdd(vdd), .A(_8667_), .B(_8670_), .Y(_8671_) );
OAI21X1 OAI21X1_1267 ( .gnd(gnd), .vdd(vdd), .A(_8666_), .B(_8671_), .C(micro_hash_ucr_2_pipe70_bF_buf1), .Y(_8672_) );
AOI21X1 AOI21X1_775 ( .gnd(gnd), .vdd(vdd), .A(_8666_), .B(_8671_), .C(_8672_), .Y(_8673_) );
OAI21X1 OAI21X1_1268 ( .gnd(gnd), .vdd(vdd), .A(H_2_21_), .B(_8641_), .C(_4496__bF_buf8), .Y(_8674_) );
NOR2X1 NOR2X1_743 ( .gnd(gnd), .vdd(vdd), .A(_8674_), .B(_8673_), .Y(_4494__21_) );
XOR2X1 XOR2X1_78 ( .gnd(gnd), .vdd(vdd), .A(H_2_22_), .B(micro_hash_ucr_2_c_6_), .Y(_8675_) );
INVX1 INVX1_326 ( .gnd(gnd), .vdd(vdd), .A(_8670_), .Y(_8676_) );
OAI21X1 OAI21X1_1269 ( .gnd(gnd), .vdd(vdd), .A(_8666_), .B(_8667_), .C(_8676_), .Y(_8677_) );
XNOR2X1 XNOR2X1_199 ( .gnd(gnd), .vdd(vdd), .A(_8677_), .B(_8675_), .Y(_8678_) );
OAI21X1 OAI21X1_1270 ( .gnd(gnd), .vdd(vdd), .A(H_2_22_), .B(_8641_), .C(_4496__bF_buf7), .Y(_8679_) );
AOI21X1 AOI21X1_776 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe70_bF_buf0), .B(_8678_), .C(_8679_), .Y(_4494__22_) );
INVX1 INVX1_327 ( .gnd(gnd), .vdd(vdd), .A(H_2_22_), .Y(_8680_) );
INVX2 INVX2_125 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_6_), .Y(_8681_) );
NAND2X1 NAND2X1_584 ( .gnd(gnd), .vdd(vdd), .A(_8675_), .B(_8677_), .Y(_8682_) );
OAI21X1 OAI21X1_1271 ( .gnd(gnd), .vdd(vdd), .A(_8680_), .B(_8681_), .C(_8682_), .Y(_8683_) );
XOR2X1 XOR2X1_79 ( .gnd(gnd), .vdd(vdd), .A(H_2_23_), .B(micro_hash_ucr_2_c_7_), .Y(_8684_) );
XNOR2X1 XNOR2X1_200 ( .gnd(gnd), .vdd(vdd), .A(_8683_), .B(_8684_), .Y(_8685_) );
OAI21X1 OAI21X1_1272 ( .gnd(gnd), .vdd(vdd), .A(H_2_23_), .B(_8641_), .C(_4496__bF_buf6), .Y(_8686_) );
AOI21X1 AOI21X1_777 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe70_bF_buf3), .B(_8685_), .C(_8686_), .Y(_4494__23_) );
INVX2 INVX2_126 ( .gnd(gnd), .vdd(vdd), .A(H_2_8_), .Y(_8687_) );
INVX8 INVX8_99 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe70_bF_buf2), .Y(_8688_) );
OAI21X1 OAI21X1_1273 ( .gnd(gnd), .vdd(vdd), .A(_8688__bF_buf3), .B(micro_hash_ucr_2_b_0_bF_buf3_), .C(_8641_), .Y(_8689_) );
INVX8 INVX8_100 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_0_bF_buf2_), .Y(_8690_) );
NOR2X1 NOR2X1_744 ( .gnd(gnd), .vdd(vdd), .A(_8687_), .B(_8690_), .Y(_8691_) );
INVX1 INVX1_328 ( .gnd(gnd), .vdd(vdd), .A(_8691_), .Y(_8692_) );
OAI21X1 OAI21X1_1274 ( .gnd(gnd), .vdd(vdd), .A(_8692_), .B(_8688__bF_buf2), .C(_4496__bF_buf5), .Y(_8693_) );
AOI21X1 AOI21X1_778 ( .gnd(gnd), .vdd(vdd), .A(_8687_), .B(_8689_), .C(_8693_), .Y(_4494__8_) );
INVX2 INVX2_127 ( .gnd(gnd), .vdd(vdd), .A(H_2_9_), .Y(_8694_) );
NOR2X1 NOR2X1_745 ( .gnd(gnd), .vdd(vdd), .A(H_2_9_), .B(micro_hash_ucr_2_b_1_bF_buf3_), .Y(_8695_) );
INVX8 INVX8_101 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_1_bF_buf2_), .Y(_8696_) );
NOR2X1 NOR2X1_746 ( .gnd(gnd), .vdd(vdd), .A(_8694_), .B(_8696_), .Y(_8697_) );
NOR2X1 NOR2X1_747 ( .gnd(gnd), .vdd(vdd), .A(_8695_), .B(_8697_), .Y(_8698_) );
AOI21X1 AOI21X1_779 ( .gnd(gnd), .vdd(vdd), .A(_8691_), .B(_8698_), .C(_8688__bF_buf1), .Y(_4570_) );
OAI21X1 OAI21X1_1275 ( .gnd(gnd), .vdd(vdd), .A(_8691_), .B(_8698_), .C(_4570_), .Y(_4571_) );
OAI21X1 OAI21X1_1276 ( .gnd(gnd), .vdd(vdd), .A(_8694_), .B(_8641_), .C(_4571_), .Y(_4572_) );
AND2X2 AND2X2_261 ( .gnd(gnd), .vdd(vdd), .A(_4572_), .B(_4496__bF_buf4), .Y(_4494__9_) );
INVX2 INVX2_128 ( .gnd(gnd), .vdd(vdd), .A(H_2_10_), .Y(_4573_) );
INVX1 INVX1_329 ( .gnd(gnd), .vdd(vdd), .A(_8697_), .Y(_4574_) );
OAI21X1 OAI21X1_1277 ( .gnd(gnd), .vdd(vdd), .A(_8692_), .B(_8695_), .C(_4574_), .Y(_4575_) );
XOR2X1 XOR2X1_80 ( .gnd(gnd), .vdd(vdd), .A(H_2_10_), .B(micro_hash_ucr_2_b_2_bF_buf3_), .Y(_4576_) );
INVX1 INVX1_330 ( .gnd(gnd), .vdd(vdd), .A(_4575_), .Y(_4577_) );
INVX1 INVX1_331 ( .gnd(gnd), .vdd(vdd), .A(_4576_), .Y(_4578_) );
NOR2X1 NOR2X1_748 ( .gnd(gnd), .vdd(vdd), .A(_4578_), .B(_4577_), .Y(_4579_) );
NOR2X1 NOR2X1_749 ( .gnd(gnd), .vdd(vdd), .A(_8688__bF_buf0), .B(_4579_), .Y(_4580_) );
OAI21X1 OAI21X1_1278 ( .gnd(gnd), .vdd(vdd), .A(_4575_), .B(_4576_), .C(_4580_), .Y(_4581_) );
OAI21X1 OAI21X1_1279 ( .gnd(gnd), .vdd(vdd), .A(_4573_), .B(_8641_), .C(_4581_), .Y(_4582_) );
AND2X2 AND2X2_262 ( .gnd(gnd), .vdd(vdd), .A(_4582_), .B(_4496__bF_buf3), .Y(_4494__10_) );
INVX8 INVX8_102 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_2_bF_buf2_), .Y(_4583_) );
INVX1 INVX1_332 ( .gnd(gnd), .vdd(vdd), .A(_4579_), .Y(_4584_) );
OAI21X1 OAI21X1_1280 ( .gnd(gnd), .vdd(vdd), .A(_4573_), .B(_4583_), .C(_4584_), .Y(_4585_) );
NOR2X1 NOR2X1_750 ( .gnd(gnd), .vdd(vdd), .A(H_2_11_), .B(micro_hash_ucr_2_b_3_bF_buf3_), .Y(_4586_) );
INVX1 INVX1_333 ( .gnd(gnd), .vdd(vdd), .A(H_2_11_), .Y(_4587_) );
INVX8 INVX8_103 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_3_bF_buf2_), .Y(_4588_) );
NOR2X1 NOR2X1_751 ( .gnd(gnd), .vdd(vdd), .A(_4587_), .B(_4588_), .Y(_4589_) );
OR2X2 OR2X2_45 ( .gnd(gnd), .vdd(vdd), .A(_4589_), .B(_4586_), .Y(_4590_) );
OAI21X1 OAI21X1_1281 ( .gnd(gnd), .vdd(vdd), .A(_4585_), .B(_4590_), .C(micro_hash_ucr_2_pipe70_bF_buf1), .Y(_4591_) );
AOI21X1 AOI21X1_780 ( .gnd(gnd), .vdd(vdd), .A(_4585_), .B(_4590_), .C(_4591_), .Y(_4592_) );
OAI21X1 OAI21X1_1282 ( .gnd(gnd), .vdd(vdd), .A(H_2_11_), .B(_8641_), .C(_4496__bF_buf2), .Y(_4593_) );
NOR2X1 NOR2X1_752 ( .gnd(gnd), .vdd(vdd), .A(_4593_), .B(_4592_), .Y(_4494__11_) );
INVX8 INVX8_104 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf1), .Y(_4594_) );
XOR2X1 XOR2X1_81 ( .gnd(gnd), .vdd(vdd), .A(H_2_12_), .B(micro_hash_ucr_2_b_4_bF_buf3_), .Y(_4595_) );
INVX1 INVX1_334 ( .gnd(gnd), .vdd(vdd), .A(_4586_), .Y(_4596_) );
AOI21X1 AOI21X1_781 ( .gnd(gnd), .vdd(vdd), .A(_4596_), .B(_4585_), .C(_4589_), .Y(_4597_) );
XNOR2X1 XNOR2X1_201 ( .gnd(gnd), .vdd(vdd), .A(_4597_), .B(_4595_), .Y(_4598_) );
INVX1 INVX1_335 ( .gnd(gnd), .vdd(vdd), .A(H_2_12_), .Y(_4599_) );
OAI21X1 OAI21X1_1283 ( .gnd(gnd), .vdd(vdd), .A(_4599_), .B(micro_hash_ucr_2_pipe5), .C(_8688__bF_buf3), .Y(_4600_) );
OAI21X1 OAI21X1_1284 ( .gnd(gnd), .vdd(vdd), .A(_4598_), .B(_8688__bF_buf2), .C(_4600_), .Y(_4601_) );
NOR2X1 NOR2X1_753 ( .gnd(gnd), .vdd(vdd), .A(_4594__bF_buf12), .B(_4601_), .Y(_4494__12_) );
NAND2X1 NAND2X1_585 ( .gnd(gnd), .vdd(vdd), .A(H_2_12_), .B(micro_hash_ucr_2_b_4_bF_buf2_), .Y(_4602_) );
INVX1 INVX1_336 ( .gnd(gnd), .vdd(vdd), .A(_4595_), .Y(_4603_) );
OAI21X1 OAI21X1_1285 ( .gnd(gnd), .vdd(vdd), .A(_4597_), .B(_4603_), .C(_4602_), .Y(_4604_) );
INVX2 INVX2_129 ( .gnd(gnd), .vdd(vdd), .A(_4604_), .Y(_4605_) );
NOR2X1 NOR2X1_754 ( .gnd(gnd), .vdd(vdd), .A(H_2_13_), .B(micro_hash_ucr_2_b_5_bF_buf3_), .Y(_4606_) );
INVX2 INVX2_130 ( .gnd(gnd), .vdd(vdd), .A(H_2_13_), .Y(_4607_) );
INVX8 INVX8_105 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_5_bF_buf2_), .Y(_4608_) );
NOR2X1 NOR2X1_755 ( .gnd(gnd), .vdd(vdd), .A(_4607_), .B(_4608__bF_buf3), .Y(_4609_) );
NOR2X1 NOR2X1_756 ( .gnd(gnd), .vdd(vdd), .A(_4606_), .B(_4609_), .Y(_4610_) );
AND2X2 AND2X2_263 ( .gnd(gnd), .vdd(vdd), .A(_4605_), .B(_4610_), .Y(_4611_) );
OAI21X1 OAI21X1_1286 ( .gnd(gnd), .vdd(vdd), .A(_4605_), .B(_4610_), .C(micro_hash_ucr_2_pipe70_bF_buf0), .Y(_4612_) );
OAI21X1 OAI21X1_1287 ( .gnd(gnd), .vdd(vdd), .A(_4607_), .B(micro_hash_ucr_2_pipe5), .C(_8688__bF_buf1), .Y(_4613_) );
OAI21X1 OAI21X1_1288 ( .gnd(gnd), .vdd(vdd), .A(_4611_), .B(_4612_), .C(_4613_), .Y(_4614_) );
NOR2X1 NOR2X1_757 ( .gnd(gnd), .vdd(vdd), .A(_4594__bF_buf11), .B(_4614_), .Y(_4494__13_) );
XOR2X1 XOR2X1_82 ( .gnd(gnd), .vdd(vdd), .A(H_2_14_), .B(micro_hash_ucr_2_b_6_), .Y(_4615_) );
INVX1 INVX1_337 ( .gnd(gnd), .vdd(vdd), .A(_4609_), .Y(_4616_) );
OAI21X1 OAI21X1_1289 ( .gnd(gnd), .vdd(vdd), .A(_4605_), .B(_4606_), .C(_4616_), .Y(_4617_) );
XNOR2X1 XNOR2X1_202 ( .gnd(gnd), .vdd(vdd), .A(_4617_), .B(_4615_), .Y(_4618_) );
INVX1 INVX1_338 ( .gnd(gnd), .vdd(vdd), .A(H_2_14_), .Y(_4619_) );
OAI21X1 OAI21X1_1290 ( .gnd(gnd), .vdd(vdd), .A(_4619_), .B(micro_hash_ucr_2_pipe5), .C(_8688__bF_buf0), .Y(_4620_) );
NAND2X1 NAND2X1_586 ( .gnd(gnd), .vdd(vdd), .A(_4620_), .B(_4496__bF_buf0), .Y(_4621_) );
AOI21X1 AOI21X1_782 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe70_bF_buf3), .B(_4618_), .C(_4621_), .Y(_4494__14_) );
INVX8 INVX8_106 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_6_), .Y(_4622_) );
NAND2X1 NAND2X1_587 ( .gnd(gnd), .vdd(vdd), .A(_4615_), .B(_4617_), .Y(_4623_) );
OAI21X1 OAI21X1_1291 ( .gnd(gnd), .vdd(vdd), .A(_4619_), .B(_4622__bF_buf3), .C(_4623_), .Y(_4624_) );
XOR2X1 XOR2X1_83 ( .gnd(gnd), .vdd(vdd), .A(H_2_15_), .B(micro_hash_ucr_2_b_7_bF_buf3_), .Y(_4625_) );
XNOR2X1 XNOR2X1_203 ( .gnd(gnd), .vdd(vdd), .A(_4624_), .B(_4625_), .Y(_4626_) );
OAI21X1 OAI21X1_1292 ( .gnd(gnd), .vdd(vdd), .A(H_2_15_), .B(_8641_), .C(_4496__bF_buf13), .Y(_4627_) );
AOI21X1 AOI21X1_783 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe70_bF_buf2), .B(_4626_), .C(_4627_), .Y(_4494__15_) );
INVX2 INVX2_131 ( .gnd(gnd), .vdd(vdd), .A(H_2_0_), .Y(_4628_) );
OAI21X1 OAI21X1_1293 ( .gnd(gnd), .vdd(vdd), .A(_8688__bF_buf3), .B(micro_hash_ucr_2_a_0_), .C(_8641_), .Y(_4629_) );
INVX8 INVX8_107 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_0_), .Y(_4630_) );
NOR2X1 NOR2X1_758 ( .gnd(gnd), .vdd(vdd), .A(_4628_), .B(_4630_), .Y(_4631_) );
INVX1 INVX1_339 ( .gnd(gnd), .vdd(vdd), .A(_4631_), .Y(_4632_) );
OAI21X1 OAI21X1_1294 ( .gnd(gnd), .vdd(vdd), .A(_4632_), .B(_8688__bF_buf2), .C(_4496__bF_buf12), .Y(_4633_) );
AOI21X1 AOI21X1_784 ( .gnd(gnd), .vdd(vdd), .A(_4628_), .B(_4629_), .C(_4633_), .Y(_4494__0_) );
INVX1 INVX1_340 ( .gnd(gnd), .vdd(vdd), .A(H_2_1_), .Y(_4634_) );
NOR2X1 NOR2X1_759 ( .gnd(gnd), .vdd(vdd), .A(H_2_1_), .B(micro_hash_ucr_2_a_1_bF_buf3_), .Y(_4635_) );
INVX8 INVX8_108 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_1_bF_buf2_), .Y(_4636_) );
NOR2X1 NOR2X1_760 ( .gnd(gnd), .vdd(vdd), .A(_4634_), .B(_4636_), .Y(_4637_) );
NOR2X1 NOR2X1_761 ( .gnd(gnd), .vdd(vdd), .A(_4635_), .B(_4637_), .Y(_4638_) );
AOI21X1 AOI21X1_785 ( .gnd(gnd), .vdd(vdd), .A(_4631_), .B(_4638_), .C(_8688__bF_buf1), .Y(_4639_) );
OAI21X1 OAI21X1_1295 ( .gnd(gnd), .vdd(vdd), .A(_4631_), .B(_4638_), .C(_4639_), .Y(_4640_) );
OAI21X1 OAI21X1_1296 ( .gnd(gnd), .vdd(vdd), .A(_4634_), .B(_8641_), .C(_4640_), .Y(_4641_) );
AND2X2 AND2X2_264 ( .gnd(gnd), .vdd(vdd), .A(_4641_), .B(_4496__bF_buf11), .Y(_4494__1_) );
INVX1 INVX1_341 ( .gnd(gnd), .vdd(vdd), .A(_4637_), .Y(_4642_) );
OAI21X1 OAI21X1_1297 ( .gnd(gnd), .vdd(vdd), .A(_4632_), .B(_4635_), .C(_4642_), .Y(_4643_) );
XOR2X1 XOR2X1_84 ( .gnd(gnd), .vdd(vdd), .A(H_2_2_), .B(micro_hash_ucr_2_a_2_), .Y(_4644_) );
INVX1 INVX1_342 ( .gnd(gnd), .vdd(vdd), .A(_4643_), .Y(_4645_) );
INVX1 INVX1_343 ( .gnd(gnd), .vdd(vdd), .A(_4644_), .Y(_4646_) );
NOR2X1 NOR2X1_762 ( .gnd(gnd), .vdd(vdd), .A(_4646_), .B(_4645_), .Y(_4647_) );
NOR2X1 NOR2X1_763 ( .gnd(gnd), .vdd(vdd), .A(_8688__bF_buf0), .B(_4647_), .Y(_4648_) );
OAI21X1 OAI21X1_1298 ( .gnd(gnd), .vdd(vdd), .A(_4643_), .B(_4644_), .C(_4648_), .Y(_4649_) );
NAND2X1 NAND2X1_588 ( .gnd(gnd), .vdd(vdd), .A(H_2_2_), .B(_8629_), .Y(_4650_) );
AOI21X1 AOI21X1_786 ( .gnd(gnd), .vdd(vdd), .A(_4650_), .B(_4649_), .C(_4594__bF_buf10), .Y(_4494__2_) );
AOI21X1 AOI21X1_787 ( .gnd(gnd), .vdd(vdd), .A(H_2_2_), .B(micro_hash_ucr_2_a_2_), .C(_4647_), .Y(_4651_) );
NOR2X1 NOR2X1_764 ( .gnd(gnd), .vdd(vdd), .A(H_2_3_), .B(micro_hash_ucr_2_a_3_), .Y(_4652_) );
INVX2 INVX2_132 ( .gnd(gnd), .vdd(vdd), .A(H_2_3_), .Y(_4653_) );
INVX8 INVX8_109 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_3_), .Y(_4654_) );
NOR2X1 NOR2X1_765 ( .gnd(gnd), .vdd(vdd), .A(_4653_), .B(_4654__bF_buf3), .Y(_4655_) );
NOR2X1 NOR2X1_766 ( .gnd(gnd), .vdd(vdd), .A(_4652_), .B(_4655_), .Y(_4656_) );
AND2X2 AND2X2_265 ( .gnd(gnd), .vdd(vdd), .A(_4651_), .B(_4656_), .Y(_4657_) );
OAI21X1 OAI21X1_1299 ( .gnd(gnd), .vdd(vdd), .A(_4651_), .B(_4656_), .C(micro_hash_ucr_2_pipe70_bF_buf1), .Y(_4658_) );
OAI21X1 OAI21X1_1300 ( .gnd(gnd), .vdd(vdd), .A(_4653_), .B(micro_hash_ucr_2_pipe5), .C(_8688__bF_buf3), .Y(_4659_) );
OAI21X1 OAI21X1_1301 ( .gnd(gnd), .vdd(vdd), .A(_4657_), .B(_4658_), .C(_4659_), .Y(_4660_) );
NOR2X1 NOR2X1_767 ( .gnd(gnd), .vdd(vdd), .A(_4594__bF_buf9), .B(_4660_), .Y(_4494__3_) );
XOR2X1 XOR2X1_85 ( .gnd(gnd), .vdd(vdd), .A(H_2_4_), .B(micro_hash_ucr_2_a_4_), .Y(_4661_) );
INVX1 INVX1_344 ( .gnd(gnd), .vdd(vdd), .A(_4655_), .Y(_4662_) );
OAI21X1 OAI21X1_1302 ( .gnd(gnd), .vdd(vdd), .A(_4651_), .B(_4652_), .C(_4662_), .Y(_4663_) );
XNOR2X1 XNOR2X1_204 ( .gnd(gnd), .vdd(vdd), .A(_4663_), .B(_4661_), .Y(_4664_) );
INVX2 INVX2_133 ( .gnd(gnd), .vdd(vdd), .A(H_2_4_), .Y(_4665_) );
OAI21X1 OAI21X1_1303 ( .gnd(gnd), .vdd(vdd), .A(_4665_), .B(micro_hash_ucr_2_pipe5), .C(_8688__bF_buf2), .Y(_4666_) );
NAND2X1 NAND2X1_589 ( .gnd(gnd), .vdd(vdd), .A(_4666_), .B(_4496__bF_buf10), .Y(_4667_) );
AOI21X1 AOI21X1_788 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe70_bF_buf0), .B(_4664_), .C(_4667_), .Y(_4494__4_) );
INVX8 INVX8_110 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_4_), .Y(_4668_) );
NAND2X1 NAND2X1_590 ( .gnd(gnd), .vdd(vdd), .A(_4661_), .B(_4663_), .Y(_4669_) );
OAI21X1 OAI21X1_1304 ( .gnd(gnd), .vdd(vdd), .A(_4665_), .B(_4668__bF_buf3), .C(_4669_), .Y(_4670_) );
INVX2 INVX2_134 ( .gnd(gnd), .vdd(vdd), .A(_4670_), .Y(_4671_) );
NOR2X1 NOR2X1_768 ( .gnd(gnd), .vdd(vdd), .A(H_2_5_), .B(micro_hash_ucr_2_a_5_bF_buf3_), .Y(_4672_) );
INVX2 INVX2_135 ( .gnd(gnd), .vdd(vdd), .A(H_2_5_), .Y(_4673_) );
INVX8 INVX8_111 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_5_bF_buf2_), .Y(_4674_) );
NOR2X1 NOR2X1_769 ( .gnd(gnd), .vdd(vdd), .A(_4673_), .B(_4674__bF_buf3), .Y(_4675_) );
NOR2X1 NOR2X1_770 ( .gnd(gnd), .vdd(vdd), .A(_4672_), .B(_4675_), .Y(_4676_) );
AND2X2 AND2X2_266 ( .gnd(gnd), .vdd(vdd), .A(_4671_), .B(_4676_), .Y(_4677_) );
OAI21X1 OAI21X1_1305 ( .gnd(gnd), .vdd(vdd), .A(_4671_), .B(_4676_), .C(micro_hash_ucr_2_pipe70_bF_buf3), .Y(_4678_) );
OAI21X1 OAI21X1_1306 ( .gnd(gnd), .vdd(vdd), .A(_4673_), .B(micro_hash_ucr_2_pipe5), .C(_8688__bF_buf1), .Y(_4679_) );
OAI21X1 OAI21X1_1307 ( .gnd(gnd), .vdd(vdd), .A(_4677_), .B(_4678_), .C(_4679_), .Y(_4680_) );
NOR2X1 NOR2X1_771 ( .gnd(gnd), .vdd(vdd), .A(_4594__bF_buf8), .B(_4680_), .Y(_4494__5_) );
XOR2X1 XOR2X1_86 ( .gnd(gnd), .vdd(vdd), .A(H_2_6_), .B(micro_hash_ucr_2_a_6_bF_buf3_), .Y(_4681_) );
INVX1 INVX1_345 ( .gnd(gnd), .vdd(vdd), .A(_4675_), .Y(_4682_) );
OAI21X1 OAI21X1_1308 ( .gnd(gnd), .vdd(vdd), .A(_4671_), .B(_4672_), .C(_4682_), .Y(_4683_) );
XOR2X1 XOR2X1_87 ( .gnd(gnd), .vdd(vdd), .A(_4683_), .B(_4681_), .Y(_4684_) );
INVX1 INVX1_346 ( .gnd(gnd), .vdd(vdd), .A(H_2_6_), .Y(_4685_) );
OAI21X1 OAI21X1_1309 ( .gnd(gnd), .vdd(vdd), .A(_4685_), .B(micro_hash_ucr_2_pipe5), .C(_8688__bF_buf0), .Y(_4686_) );
OAI21X1 OAI21X1_1310 ( .gnd(gnd), .vdd(vdd), .A(_4684_), .B(_8688__bF_buf3), .C(_4686_), .Y(_4687_) );
NOR2X1 NOR2X1_772 ( .gnd(gnd), .vdd(vdd), .A(_4594__bF_buf7), .B(_4687_), .Y(_4494__6_) );
INVX8 INVX8_112 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_6_bF_buf2_), .Y(_4688_) );
NAND2X1 NAND2X1_591 ( .gnd(gnd), .vdd(vdd), .A(_4681_), .B(_4683_), .Y(_4689_) );
OAI21X1 OAI21X1_1311 ( .gnd(gnd), .vdd(vdd), .A(_4685_), .B(_4688_), .C(_4689_), .Y(_4690_) );
XNOR2X1 XNOR2X1_205 ( .gnd(gnd), .vdd(vdd), .A(H_2_7_), .B(micro_hash_ucr_2_a_7_), .Y(_4691_) );
AND2X2 AND2X2_267 ( .gnd(gnd), .vdd(vdd), .A(_4690_), .B(_4691_), .Y(_4692_) );
OAI21X1 OAI21X1_1312 ( .gnd(gnd), .vdd(vdd), .A(_4690_), .B(_4691_), .C(micro_hash_ucr_2_pipe70_bF_buf2), .Y(_4693_) );
INVX1 INVX1_347 ( .gnd(gnd), .vdd(vdd), .A(H_2_7_), .Y(_4694_) );
OAI21X1 OAI21X1_1313 ( .gnd(gnd), .vdd(vdd), .A(_4694_), .B(micro_hash_ucr_2_pipe5), .C(_8688__bF_buf2), .Y(_4695_) );
OAI21X1 OAI21X1_1314 ( .gnd(gnd), .vdd(vdd), .A(_4692_), .B(_4693_), .C(_4695_), .Y(_4696_) );
NOR2X1 NOR2X1_773 ( .gnd(gnd), .vdd(vdd), .A(_4594__bF_buf6), .B(_4696_), .Y(_4494__7_) );
INVX2 INVX2_136 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_152_), .Y(_4697_) );
INVX1 INVX1_348 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_200_), .Y(_4698_) );
OAI21X1 OAI21X1_1315 ( .gnd(gnd), .vdd(vdd), .A(_4697_), .B(micro_hash_ucr_2_Wx_112_), .C(_4698_), .Y(_4699_) );
AOI21X1 AOI21X1_789 ( .gnd(gnd), .vdd(vdd), .A(_4697_), .B(micro_hash_ucr_2_Wx_112_), .C(_4699_), .Y(_4700_) );
NOR2X1 NOR2X1_774 ( .gnd(gnd), .vdd(vdd), .A(_4700_), .B(_4594__bF_buf5), .Y(_4490__224_) );
INVX4 INVX4_57 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_153_), .Y(_4701_) );
INVX2 INVX2_137 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_201_), .Y(_4702_) );
OAI21X1 OAI21X1_1316 ( .gnd(gnd), .vdd(vdd), .A(_4701_), .B(micro_hash_ucr_2_Wx_113_), .C(_4702_), .Y(_4703_) );
AOI21X1 AOI21X1_790 ( .gnd(gnd), .vdd(vdd), .A(_4701_), .B(micro_hash_ucr_2_Wx_113_), .C(_4703_), .Y(_4704_) );
NOR2X1 NOR2X1_775 ( .gnd(gnd), .vdd(vdd), .A(_4704_), .B(_4594__bF_buf4), .Y(_4490__225_) );
INVX2 INVX2_138 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_154_), .Y(_4705_) );
INVX2 INVX2_139 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_202_), .Y(_4706_) );
OAI21X1 OAI21X1_1317 ( .gnd(gnd), .vdd(vdd), .A(_4705_), .B(micro_hash_ucr_2_Wx_114_), .C(_4706_), .Y(_4707_) );
AOI21X1 AOI21X1_791 ( .gnd(gnd), .vdd(vdd), .A(_4705_), .B(micro_hash_ucr_2_Wx_114_), .C(_4707_), .Y(_4708_) );
NOR2X1 NOR2X1_776 ( .gnd(gnd), .vdd(vdd), .A(_4708_), .B(_4594__bF_buf3), .Y(_4490__226_) );
INVX2 INVX2_140 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_155_), .Y(_4709_) );
INVX1 INVX1_349 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_203_), .Y(_4710_) );
OAI21X1 OAI21X1_1318 ( .gnd(gnd), .vdd(vdd), .A(_4709_), .B(micro_hash_ucr_2_Wx_115_), .C(_4710_), .Y(_4711_) );
AOI21X1 AOI21X1_792 ( .gnd(gnd), .vdd(vdd), .A(_4709_), .B(micro_hash_ucr_2_Wx_115_), .C(_4711_), .Y(_4712_) );
NOR2X1 NOR2X1_777 ( .gnd(gnd), .vdd(vdd), .A(_4712_), .B(_4594__bF_buf2), .Y(_4490__227_) );
INVX2 INVX2_141 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_156_), .Y(_4713_) );
AOI21X1 AOI21X1_793 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_116_), .B(_4713_), .C(micro_hash_ucr_2_Wx_204_), .Y(_4714_) );
OAI21X1 OAI21X1_1319 ( .gnd(gnd), .vdd(vdd), .A(_4713_), .B(micro_hash_ucr_2_Wx_116_), .C(_4714_), .Y(_4715_) );
AND2X2 AND2X2_268 ( .gnd(gnd), .vdd(vdd), .A(_4715_), .B(_4496__bF_buf9), .Y(_4490__228_) );
INVX2 INVX2_142 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_157_), .Y(_4716_) );
AOI21X1 AOI21X1_794 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_117_), .B(_4716_), .C(micro_hash_ucr_2_Wx_205_), .Y(_4717_) );
OAI21X1 OAI21X1_1320 ( .gnd(gnd), .vdd(vdd), .A(_4716_), .B(micro_hash_ucr_2_Wx_117_), .C(_4717_), .Y(_4718_) );
AND2X2 AND2X2_269 ( .gnd(gnd), .vdd(vdd), .A(_4718_), .B(_4496__bF_buf8), .Y(_4490__229_) );
INVX4 INVX4_58 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_158_), .Y(_4719_) );
INVX2 INVX2_143 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_206_), .Y(_4720_) );
OAI21X1 OAI21X1_1321 ( .gnd(gnd), .vdd(vdd), .A(_4719_), .B(micro_hash_ucr_2_Wx_118_), .C(_4720_), .Y(_4721_) );
AOI21X1 AOI21X1_795 ( .gnd(gnd), .vdd(vdd), .A(_4719_), .B(micro_hash_ucr_2_Wx_118_), .C(_4721_), .Y(_4722_) );
NOR2X1 NOR2X1_778 ( .gnd(gnd), .vdd(vdd), .A(_4722_), .B(_4594__bF_buf1), .Y(_4490__230_) );
INVX2 INVX2_144 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_159_), .Y(_4723_) );
AOI21X1 AOI21X1_796 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_119_), .B(_4723_), .C(micro_hash_ucr_2_Wx_207_), .Y(_4724_) );
OAI21X1 OAI21X1_1322 ( .gnd(gnd), .vdd(vdd), .A(_4723_), .B(micro_hash_ucr_2_Wx_119_), .C(_4724_), .Y(_4725_) );
AND2X2 AND2X2_270 ( .gnd(gnd), .vdd(vdd), .A(_4725_), .B(_4496__bF_buf7), .Y(_4490__231_) );
INVX1 INVX1_350 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_216_), .Y(_4726_) );
XNOR2X1 XNOR2X1_206 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_168_), .B(micro_hash_ucr_2_Wx_128_), .Y(_4727_) );
AOI21X1 AOI21X1_797 ( .gnd(gnd), .vdd(vdd), .A(_4726_), .B(_4727_), .C(_4594__bF_buf0), .Y(_4490__240_) );
INVX2 INVX2_145 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_169_), .Y(_4728_) );
INVX1 INVX1_351 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_217_), .Y(_4729_) );
OAI21X1 OAI21X1_1323 ( .gnd(gnd), .vdd(vdd), .A(_4728_), .B(micro_hash_ucr_2_Wx_129_), .C(_4729_), .Y(_4730_) );
AOI21X1 AOI21X1_798 ( .gnd(gnd), .vdd(vdd), .A(_4728_), .B(micro_hash_ucr_2_Wx_129_), .C(_4730_), .Y(_4731_) );
NOR2X1 NOR2X1_779 ( .gnd(gnd), .vdd(vdd), .A(_4731_), .B(_4594__bF_buf12), .Y(_4490__241_) );
INVX4 INVX4_59 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_170_), .Y(_4732_) );
INVX2 INVX2_146 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_218_), .Y(_4733_) );
OAI21X1 OAI21X1_1324 ( .gnd(gnd), .vdd(vdd), .A(_4732_), .B(micro_hash_ucr_2_Wx_130_), .C(_4733_), .Y(_4734_) );
AOI21X1 AOI21X1_799 ( .gnd(gnd), .vdd(vdd), .A(_4732_), .B(micro_hash_ucr_2_Wx_130_), .C(_4734_), .Y(_4735_) );
NOR2X1 NOR2X1_780 ( .gnd(gnd), .vdd(vdd), .A(_4735_), .B(_4594__bF_buf11), .Y(_4490__242_) );
INVX2 INVX2_147 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_171_), .Y(_4736_) );
INVX1 INVX1_352 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_219_), .Y(_4737_) );
OAI21X1 OAI21X1_1325 ( .gnd(gnd), .vdd(vdd), .A(_4736_), .B(micro_hash_ucr_2_Wx_131_), .C(_4737_), .Y(_4738_) );
AOI21X1 AOI21X1_800 ( .gnd(gnd), .vdd(vdd), .A(_4736_), .B(micro_hash_ucr_2_Wx_131_), .C(_4738_), .Y(_4739_) );
NOR2X1 NOR2X1_781 ( .gnd(gnd), .vdd(vdd), .A(_4739_), .B(_4594__bF_buf10), .Y(_4490__243_) );
INVX2 INVX2_148 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_172_), .Y(_4740_) );
AOI21X1 AOI21X1_801 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_132_), .B(_4740_), .C(micro_hash_ucr_2_Wx_220_), .Y(_4741_) );
OAI21X1 OAI21X1_1326 ( .gnd(gnd), .vdd(vdd), .A(_4740_), .B(micro_hash_ucr_2_Wx_132_), .C(_4741_), .Y(_4742_) );
AND2X2 AND2X2_271 ( .gnd(gnd), .vdd(vdd), .A(_4742_), .B(_4496__bF_buf6), .Y(_4490__244_) );
INVX2 INVX2_149 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_173_), .Y(_4743_) );
INVX1 INVX1_353 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_221_), .Y(_4744_) );
OAI21X1 OAI21X1_1327 ( .gnd(gnd), .vdd(vdd), .A(_4743_), .B(micro_hash_ucr_2_Wx_133_), .C(_4744_), .Y(_4745_) );
AOI21X1 AOI21X1_802 ( .gnd(gnd), .vdd(vdd), .A(_4743_), .B(micro_hash_ucr_2_Wx_133_), .C(_4745_), .Y(_4746_) );
NOR2X1 NOR2X1_782 ( .gnd(gnd), .vdd(vdd), .A(_4746_), .B(_4594__bF_buf9), .Y(_4490__245_) );
INVX2 INVX2_150 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_174_), .Y(_4747_) );
INVX2 INVX2_151 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_222_), .Y(_4748_) );
OAI21X1 OAI21X1_1328 ( .gnd(gnd), .vdd(vdd), .A(_4747_), .B(micro_hash_ucr_2_Wx_134_), .C(_4748_), .Y(_4749_) );
AOI21X1 AOI21X1_803 ( .gnd(gnd), .vdd(vdd), .A(_4747_), .B(micro_hash_ucr_2_Wx_134_), .C(_4749_), .Y(_4750_) );
NOR2X1 NOR2X1_783 ( .gnd(gnd), .vdd(vdd), .A(_4750_), .B(_4594__bF_buf8), .Y(_4490__246_) );
INVX4 INVX4_60 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_175_), .Y(_4751_) );
AOI21X1 AOI21X1_804 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_135_), .B(_4751_), .C(micro_hash_ucr_2_Wx_223_), .Y(_4752_) );
OAI21X1 OAI21X1_1329 ( .gnd(gnd), .vdd(vdd), .A(_4751_), .B(micro_hash_ucr_2_Wx_135_), .C(_4752_), .Y(_4753_) );
AND2X2 AND2X2_272 ( .gnd(gnd), .vdd(vdd), .A(_4753_), .B(_4496__bF_buf5), .Y(_4490__247_) );
INVX4 INVX4_61 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_120_), .Y(_4754_) );
AOI21X1 AOI21X1_805 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_160_), .B(_4754_), .C(micro_hash_ucr_2_Wx_208_), .Y(_4755_) );
OAI21X1 OAI21X1_1330 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_160_), .B(_4754_), .C(_4755_), .Y(_4756_) );
AND2X2 AND2X2_273 ( .gnd(gnd), .vdd(vdd), .A(_4756_), .B(_4496__bF_buf4), .Y(_4490__232_) );
INVX2 INVX2_152 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_161_), .Y(_4757_) );
AOI21X1 AOI21X1_806 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_121_), .B(_4757_), .C(micro_hash_ucr_2_Wx_209_), .Y(_4758_) );
OAI21X1 OAI21X1_1331 ( .gnd(gnd), .vdd(vdd), .A(_4757_), .B(micro_hash_ucr_2_Wx_121_), .C(_4758_), .Y(_4759_) );
AND2X2 AND2X2_274 ( .gnd(gnd), .vdd(vdd), .A(_4759_), .B(_4496__bF_buf3), .Y(_4490__233_) );
INVX4 INVX4_62 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_162_), .Y(_4760_) );
INVX1 INVX1_354 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_210_), .Y(_4761_) );
OAI21X1 OAI21X1_1332 ( .gnd(gnd), .vdd(vdd), .A(_4760_), .B(micro_hash_ucr_2_Wx_122_), .C(_4761_), .Y(_4762_) );
AOI21X1 AOI21X1_807 ( .gnd(gnd), .vdd(vdd), .A(_4760_), .B(micro_hash_ucr_2_Wx_122_), .C(_4762_), .Y(_4763_) );
NOR2X1 NOR2X1_784 ( .gnd(gnd), .vdd(vdd), .A(_4763_), .B(_4594__bF_buf7), .Y(_4490__234_) );
INVX2 INVX2_153 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_163_), .Y(_4764_) );
INVX1 INVX1_355 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_211_), .Y(_4765_) );
OAI21X1 OAI21X1_1333 ( .gnd(gnd), .vdd(vdd), .A(_4764_), .B(micro_hash_ucr_2_Wx_123_), .C(_4765_), .Y(_4766_) );
AOI21X1 AOI21X1_808 ( .gnd(gnd), .vdd(vdd), .A(_4764_), .B(micro_hash_ucr_2_Wx_123_), .C(_4766_), .Y(_4767_) );
NOR2X1 NOR2X1_785 ( .gnd(gnd), .vdd(vdd), .A(_4767_), .B(_4594__bF_buf6), .Y(_4490__235_) );
INVX4 INVX4_63 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_124_), .Y(_4768_) );
AOI21X1 AOI21X1_809 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_164_), .B(_4768_), .C(micro_hash_ucr_2_Wx_212_), .Y(_4769_) );
OAI21X1 OAI21X1_1334 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_164_), .B(_4768_), .C(_4769_), .Y(_4770_) );
AND2X2 AND2X2_275 ( .gnd(gnd), .vdd(vdd), .A(_4770_), .B(_4496__bF_buf2), .Y(_4490__236_) );
INVX2 INVX2_154 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_165_), .Y(_4771_) );
AOI21X1 AOI21X1_810 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_125_), .B(_4771_), .C(micro_hash_ucr_2_Wx_213_), .Y(_4772_) );
OAI21X1 OAI21X1_1335 ( .gnd(gnd), .vdd(vdd), .A(_4771_), .B(micro_hash_ucr_2_Wx_125_), .C(_4772_), .Y(_4773_) );
AND2X2 AND2X2_276 ( .gnd(gnd), .vdd(vdd), .A(_4773_), .B(_4496__bF_buf1), .Y(_4490__237_) );
INVX4 INVX4_64 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_166_), .Y(_4774_) );
INVX2 INVX2_155 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_214_), .Y(_4775_) );
OAI21X1 OAI21X1_1336 ( .gnd(gnd), .vdd(vdd), .A(_4774_), .B(micro_hash_ucr_2_Wx_126_), .C(_4775_), .Y(_4776_) );
AOI21X1 AOI21X1_811 ( .gnd(gnd), .vdd(vdd), .A(_4774_), .B(micro_hash_ucr_2_Wx_126_), .C(_4776_), .Y(_4777_) );
NOR2X1 NOR2X1_786 ( .gnd(gnd), .vdd(vdd), .A(_4777_), .B(_4594__bF_buf5), .Y(_4490__238_) );
INVX2 INVX2_156 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_167_), .Y(_4778_) );
AOI21X1 AOI21X1_812 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_127_), .B(_4778_), .C(micro_hash_ucr_2_Wx_215_), .Y(_4779_) );
OAI21X1 OAI21X1_1337 ( .gnd(gnd), .vdd(vdd), .A(_4778_), .B(micro_hash_ucr_2_Wx_127_), .C(_4779_), .Y(_4780_) );
AND2X2 AND2X2_277 ( .gnd(gnd), .vdd(vdd), .A(_4780_), .B(_4496__bF_buf0), .Y(_4490__239_) );
INVX2 INVX2_157 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_128_), .Y(_4781_) );
INVX2 INVX2_158 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_176_), .Y(_4782_) );
OAI21X1 OAI21X1_1338 ( .gnd(gnd), .vdd(vdd), .A(_4781_), .B(micro_hash_ucr_2_Wx_88_), .C(_4782_), .Y(_4783_) );
AOI21X1 AOI21X1_813 ( .gnd(gnd), .vdd(vdd), .A(_4781_), .B(micro_hash_ucr_2_Wx_88_), .C(_4783_), .Y(_4784_) );
NOR2X1 NOR2X1_787 ( .gnd(gnd), .vdd(vdd), .A(_4784_), .B(_4594__bF_buf4), .Y(_4490__200_) );
INVX4 INVX4_65 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_129_), .Y(_4785_) );
INVX4 INVX4_66 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_177_), .Y(_4786_) );
OAI21X1 OAI21X1_1339 ( .gnd(gnd), .vdd(vdd), .A(_4785_), .B(micro_hash_ucr_2_Wx_89_), .C(_4786_), .Y(_4787_) );
AOI21X1 AOI21X1_814 ( .gnd(gnd), .vdd(vdd), .A(_4785_), .B(micro_hash_ucr_2_Wx_89_), .C(_4787_), .Y(_4788_) );
NOR2X1 NOR2X1_788 ( .gnd(gnd), .vdd(vdd), .A(_4788_), .B(_4594__bF_buf3), .Y(_4490__201_) );
INVX4 INVX4_67 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_130_), .Y(_4789_) );
INVX4 INVX4_68 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_178_), .Y(_4790_) );
OAI21X1 OAI21X1_1340 ( .gnd(gnd), .vdd(vdd), .A(_4789_), .B(micro_hash_ucr_2_Wx_90_), .C(_4790_), .Y(_4791_) );
AOI21X1 AOI21X1_815 ( .gnd(gnd), .vdd(vdd), .A(_4789_), .B(micro_hash_ucr_2_Wx_90_), .C(_4791_), .Y(_4792_) );
NOR2X1 NOR2X1_789 ( .gnd(gnd), .vdd(vdd), .A(_4792_), .B(_4594__bF_buf2), .Y(_4490__202_) );
INVX2 INVX2_159 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_131_), .Y(_4793_) );
INVX2 INVX2_160 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_179_), .Y(_4794_) );
OAI21X1 OAI21X1_1341 ( .gnd(gnd), .vdd(vdd), .A(_4793_), .B(micro_hash_ucr_2_Wx_91_), .C(_4794_), .Y(_4795_) );
AOI21X1 AOI21X1_816 ( .gnd(gnd), .vdd(vdd), .A(_4793_), .B(micro_hash_ucr_2_Wx_91_), .C(_4795_), .Y(_4796_) );
NOR2X1 NOR2X1_790 ( .gnd(gnd), .vdd(vdd), .A(_4796_), .B(_4594__bF_buf1), .Y(_4490__203_) );
INVX2 INVX2_161 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_132_), .Y(_4797_) );
INVX4 INVX4_69 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_180_), .Y(_4798_) );
OAI21X1 OAI21X1_1342 ( .gnd(gnd), .vdd(vdd), .A(_4797_), .B(micro_hash_ucr_2_Wx_92_), .C(_4798_), .Y(_4799_) );
AOI21X1 AOI21X1_817 ( .gnd(gnd), .vdd(vdd), .A(_4797_), .B(micro_hash_ucr_2_Wx_92_), .C(_4799_), .Y(_4800_) );
NOR2X1 NOR2X1_791 ( .gnd(gnd), .vdd(vdd), .A(_4800_), .B(_4594__bF_buf0), .Y(_4490__204_) );
INVX2 INVX2_162 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_133_), .Y(_4801_) );
INVX2 INVX2_163 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_181_), .Y(_4802_) );
OAI21X1 OAI21X1_1343 ( .gnd(gnd), .vdd(vdd), .A(_4801_), .B(micro_hash_ucr_2_Wx_93_), .C(_4802_), .Y(_4803_) );
AOI21X1 AOI21X1_818 ( .gnd(gnd), .vdd(vdd), .A(_4801_), .B(micro_hash_ucr_2_Wx_93_), .C(_4803_), .Y(_4804_) );
NOR2X1 NOR2X1_792 ( .gnd(gnd), .vdd(vdd), .A(_4804_), .B(_4594__bF_buf12), .Y(_4490__205_) );
INVX4 INVX4_70 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_134_), .Y(_4805_) );
INVX2 INVX2_164 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_182_), .Y(_4806_) );
OAI21X1 OAI21X1_1344 ( .gnd(gnd), .vdd(vdd), .A(_4805_), .B(micro_hash_ucr_2_Wx_94_), .C(_4806_), .Y(_4807_) );
AOI21X1 AOI21X1_819 ( .gnd(gnd), .vdd(vdd), .A(_4805_), .B(micro_hash_ucr_2_Wx_94_), .C(_4807_), .Y(_4808_) );
NOR2X1 NOR2X1_793 ( .gnd(gnd), .vdd(vdd), .A(_4808_), .B(_4594__bF_buf11), .Y(_4490__206_) );
INVX4 INVX4_71 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_183_), .Y(_4809_) );
XNOR2X1 XNOR2X1_207 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_135_), .B(micro_hash_ucr_2_Wx_95_), .Y(_4810_) );
AOI21X1 AOI21X1_820 ( .gnd(gnd), .vdd(vdd), .A(_4809_), .B(_4810_), .C(_4594__bF_buf10), .Y(_4490__207_) );
INVX2 INVX2_165 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_144_), .Y(_4811_) );
INVX1 INVX1_356 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_192_), .Y(_4812_) );
OAI21X1 OAI21X1_1345 ( .gnd(gnd), .vdd(vdd), .A(_4811_), .B(micro_hash_ucr_2_Wx_104_), .C(_4812_), .Y(_4813_) );
AOI21X1 AOI21X1_821 ( .gnd(gnd), .vdd(vdd), .A(_4811_), .B(micro_hash_ucr_2_Wx_104_), .C(_4813_), .Y(_4814_) );
NOR2X1 NOR2X1_794 ( .gnd(gnd), .vdd(vdd), .A(_4814_), .B(_4594__bF_buf9), .Y(_4490__216_) );
INVX4 INVX4_72 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_145_), .Y(_4815_) );
INVX2 INVX2_166 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_193_), .Y(_4816_) );
OAI21X1 OAI21X1_1346 ( .gnd(gnd), .vdd(vdd), .A(_4815_), .B(micro_hash_ucr_2_Wx_105_), .C(_4816_), .Y(_4817_) );
AOI21X1 AOI21X1_822 ( .gnd(gnd), .vdd(vdd), .A(_4815_), .B(micro_hash_ucr_2_Wx_105_), .C(_4817_), .Y(_4818_) );
NOR2X1 NOR2X1_795 ( .gnd(gnd), .vdd(vdd), .A(_4818_), .B(_4594__bF_buf8), .Y(_4490__217_) );
INVX4 INVX4_73 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_146_), .Y(_4819_) );
INVX2 INVX2_167 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_194_), .Y(_4820_) );
OAI21X1 OAI21X1_1347 ( .gnd(gnd), .vdd(vdd), .A(_4819_), .B(micro_hash_ucr_2_Wx_106_), .C(_4820_), .Y(_4821_) );
AOI21X1 AOI21X1_823 ( .gnd(gnd), .vdd(vdd), .A(_4819_), .B(micro_hash_ucr_2_Wx_106_), .C(_4821_), .Y(_4822_) );
NOR2X1 NOR2X1_796 ( .gnd(gnd), .vdd(vdd), .A(_4822_), .B(_4594__bF_buf7), .Y(_4490__218_) );
INVX2 INVX2_168 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_147_), .Y(_4823_) );
INVX1 INVX1_357 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_195_), .Y(_4824_) );
OAI21X1 OAI21X1_1348 ( .gnd(gnd), .vdd(vdd), .A(_4823_), .B(micro_hash_ucr_2_Wx_107_), .C(_4824_), .Y(_4825_) );
AOI21X1 AOI21X1_824 ( .gnd(gnd), .vdd(vdd), .A(_4823_), .B(micro_hash_ucr_2_Wx_107_), .C(_4825_), .Y(_4826_) );
NOR2X1 NOR2X1_797 ( .gnd(gnd), .vdd(vdd), .A(_4826_), .B(_4594__bF_buf6), .Y(_4490__219_) );
INVX2 INVX2_169 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_148_), .Y(_4827_) );
AOI21X1 AOI21X1_825 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_108_), .B(_4827_), .C(micro_hash_ucr_2_Wx_196_), .Y(_4828_) );
OAI21X1 OAI21X1_1349 ( .gnd(gnd), .vdd(vdd), .A(_4827_), .B(micro_hash_ucr_2_Wx_108_), .C(_4828_), .Y(_4829_) );
AND2X2 AND2X2_278 ( .gnd(gnd), .vdd(vdd), .A(_4829_), .B(_4496__bF_buf13), .Y(_4490__220_) );
INVX2 INVX2_170 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_149_), .Y(_4830_) );
AOI21X1 AOI21X1_826 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_109_), .B(_4830_), .C(micro_hash_ucr_2_Wx_197_), .Y(_4831_) );
OAI21X1 OAI21X1_1350 ( .gnd(gnd), .vdd(vdd), .A(_4830_), .B(micro_hash_ucr_2_Wx_109_), .C(_4831_), .Y(_4832_) );
AND2X2 AND2X2_279 ( .gnd(gnd), .vdd(vdd), .A(_4832_), .B(_4496__bF_buf12), .Y(_4490__221_) );
INVX4 INVX4_74 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_150_), .Y(_4833_) );
INVX1 INVX1_358 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_198_), .Y(_4834_) );
OAI21X1 OAI21X1_1351 ( .gnd(gnd), .vdd(vdd), .A(_4833_), .B(micro_hash_ucr_2_Wx_110_), .C(_4834_), .Y(_4835_) );
AOI21X1 AOI21X1_827 ( .gnd(gnd), .vdd(vdd), .A(_4833_), .B(micro_hash_ucr_2_Wx_110_), .C(_4835_), .Y(_4836_) );
NOR2X1 NOR2X1_798 ( .gnd(gnd), .vdd(vdd), .A(_4836_), .B(_4594__bF_buf5), .Y(_4490__222_) );
INVX4 INVX4_75 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_151_), .Y(_4837_) );
AOI21X1 AOI21X1_828 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_111_), .B(_4837_), .C(micro_hash_ucr_2_Wx_199_), .Y(_4838_) );
OAI21X1 OAI21X1_1352 ( .gnd(gnd), .vdd(vdd), .A(_4837_), .B(micro_hash_ucr_2_Wx_111_), .C(_4838_), .Y(_4839_) );
AND2X2 AND2X2_280 ( .gnd(gnd), .vdd(vdd), .A(_4839_), .B(_4496__bF_buf11), .Y(_4490__223_) );
INVX4 INVX4_76 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_96_), .Y(_4840_) );
AOI21X1 AOI21X1_829 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_136_), .B(_4840_), .C(micro_hash_ucr_2_Wx_184_), .Y(_4841_) );
OAI21X1 OAI21X1_1353 ( .gnd(gnd), .vdd(vdd), .A(_4840_), .B(micro_hash_ucr_2_Wx_136_), .C(_4841_), .Y(_4842_) );
AND2X2 AND2X2_281 ( .gnd(gnd), .vdd(vdd), .A(_4842_), .B(_4496__bF_buf10), .Y(_4490__208_) );
INVX4 INVX4_77 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_97_), .Y(_4843_) );
INVX2 INVX2_171 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_185_), .Y(_4844_) );
OAI21X1 OAI21X1_1354 ( .gnd(gnd), .vdd(vdd), .A(_4843_), .B(micro_hash_ucr_2_Wx_137_), .C(_4844_), .Y(_4845_) );
AOI21X1 AOI21X1_830 ( .gnd(gnd), .vdd(vdd), .A(_4843_), .B(micro_hash_ucr_2_Wx_137_), .C(_4845_), .Y(_4846_) );
NOR2X1 NOR2X1_799 ( .gnd(gnd), .vdd(vdd), .A(_4846_), .B(_4594__bF_buf4), .Y(_4490__209_) );
INVX4 INVX4_78 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_98_), .Y(_4847_) );
INVX1 INVX1_359 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_186_), .Y(_4848_) );
OAI21X1 OAI21X1_1355 ( .gnd(gnd), .vdd(vdd), .A(_4847_), .B(micro_hash_ucr_2_Wx_138_), .C(_4848_), .Y(_4849_) );
AOI21X1 AOI21X1_831 ( .gnd(gnd), .vdd(vdd), .A(_4847_), .B(micro_hash_ucr_2_Wx_138_), .C(_4849_), .Y(_4850_) );
NOR2X1 NOR2X1_800 ( .gnd(gnd), .vdd(vdd), .A(_4850_), .B(_4594__bF_buf3), .Y(_4490__210_) );
INVX4 INVX4_79 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_99_), .Y(_4851_) );
INVX1 INVX1_360 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_187_), .Y(_4852_) );
OAI21X1 OAI21X1_1356 ( .gnd(gnd), .vdd(vdd), .A(_4851_), .B(micro_hash_ucr_2_Wx_139_), .C(_4852_), .Y(_4853_) );
AOI21X1 AOI21X1_832 ( .gnd(gnd), .vdd(vdd), .A(_4851_), .B(micro_hash_ucr_2_Wx_139_), .C(_4853_), .Y(_4854_) );
NOR2X1 NOR2X1_801 ( .gnd(gnd), .vdd(vdd), .A(_4854_), .B(_4594__bF_buf2), .Y(_4490__211_) );
INVX2 INVX2_172 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_100_), .Y(_4855_) );
AOI21X1 AOI21X1_833 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_140_), .B(_4855_), .C(micro_hash_ucr_2_Wx_188_), .Y(_4856_) );
OAI21X1 OAI21X1_1357 ( .gnd(gnd), .vdd(vdd), .A(_4855_), .B(micro_hash_ucr_2_Wx_140_), .C(_4856_), .Y(_4857_) );
AND2X2 AND2X2_282 ( .gnd(gnd), .vdd(vdd), .A(_4857_), .B(_4496__bF_buf9), .Y(_4490__212_) );
INVX4 INVX4_80 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_101_), .Y(_4858_) );
INVX1 INVX1_361 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_189_), .Y(_4859_) );
OAI21X1 OAI21X1_1358 ( .gnd(gnd), .vdd(vdd), .A(_4858_), .B(micro_hash_ucr_2_Wx_141_), .C(_4859_), .Y(_4860_) );
AOI21X1 AOI21X1_834 ( .gnd(gnd), .vdd(vdd), .A(_4858_), .B(micro_hash_ucr_2_Wx_141_), .C(_4860_), .Y(_4861_) );
NOR2X1 NOR2X1_802 ( .gnd(gnd), .vdd(vdd), .A(_4861_), .B(_4594__bF_buf1), .Y(_4490__213_) );
INVX4 INVX4_81 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_102_), .Y(_4862_) );
INVX2 INVX2_173 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_190_), .Y(_4863_) );
OAI21X1 OAI21X1_1359 ( .gnd(gnd), .vdd(vdd), .A(_4862_), .B(micro_hash_ucr_2_Wx_142_), .C(_4863_), .Y(_4864_) );
AOI21X1 AOI21X1_835 ( .gnd(gnd), .vdd(vdd), .A(_4862_), .B(micro_hash_ucr_2_Wx_142_), .C(_4864_), .Y(_4865_) );
NOR2X1 NOR2X1_803 ( .gnd(gnd), .vdd(vdd), .A(_4865_), .B(_4594__bF_buf0), .Y(_4490__214_) );
INVX4 INVX4_82 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_103_), .Y(_4866_) );
AOI21X1 AOI21X1_836 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_143_), .B(_4866_), .C(micro_hash_ucr_2_Wx_191_), .Y(_4867_) );
OAI21X1 OAI21X1_1360 ( .gnd(gnd), .vdd(vdd), .A(_4866_), .B(micro_hash_ucr_2_Wx_143_), .C(_4867_), .Y(_4868_) );
AND2X2 AND2X2_283 ( .gnd(gnd), .vdd(vdd), .A(_4868_), .B(_4496__bF_buf8), .Y(_4490__215_) );
INVX2 INVX2_174 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_104_), .Y(_4869_) );
OAI21X1 OAI21X1_1361 ( .gnd(gnd), .vdd(vdd), .A(_4869_), .B(micro_hash_ucr_2_Wx_64_), .C(_4697_), .Y(_4870_) );
AOI21X1 AOI21X1_837 ( .gnd(gnd), .vdd(vdd), .A(_4869_), .B(micro_hash_ucr_2_Wx_64_), .C(_4870_), .Y(_4871_) );
NOR2X1 NOR2X1_804 ( .gnd(gnd), .vdd(vdd), .A(_4871_), .B(_4594__bF_buf12), .Y(_4490__176_) );
INVX2 INVX2_175 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_105_), .Y(_4872_) );
OAI21X1 OAI21X1_1362 ( .gnd(gnd), .vdd(vdd), .A(_4872_), .B(micro_hash_ucr_2_Wx_65_), .C(_4701_), .Y(_4873_) );
AOI21X1 AOI21X1_838 ( .gnd(gnd), .vdd(vdd), .A(_4872_), .B(micro_hash_ucr_2_Wx_65_), .C(_4873_), .Y(_4874_) );
NOR2X1 NOR2X1_805 ( .gnd(gnd), .vdd(vdd), .A(_4874_), .B(_4594__bF_buf11), .Y(_4490__177_) );
INVX4 INVX4_83 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_106_), .Y(_4875_) );
OAI21X1 OAI21X1_1363 ( .gnd(gnd), .vdd(vdd), .A(_4875_), .B(micro_hash_ucr_2_Wx_66_), .C(_4705_), .Y(_4876_) );
AOI21X1 AOI21X1_839 ( .gnd(gnd), .vdd(vdd), .A(_4875_), .B(micro_hash_ucr_2_Wx_66_), .C(_4876_), .Y(_4877_) );
NOR2X1 NOR2X1_806 ( .gnd(gnd), .vdd(vdd), .A(_4877_), .B(_4594__bF_buf10), .Y(_4490__178_) );
INVX2 INVX2_176 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_107_), .Y(_4878_) );
OAI21X1 OAI21X1_1364 ( .gnd(gnd), .vdd(vdd), .A(_4878_), .B(micro_hash_ucr_2_Wx_67_), .C(_4709_), .Y(_4879_) );
AOI21X1 AOI21X1_840 ( .gnd(gnd), .vdd(vdd), .A(_4878_), .B(micro_hash_ucr_2_Wx_67_), .C(_4879_), .Y(_4880_) );
NOR2X1 NOR2X1_807 ( .gnd(gnd), .vdd(vdd), .A(_4880_), .B(_4594__bF_buf9), .Y(_4490__179_) );
INVX2 INVX2_177 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_108_), .Y(_4881_) );
OAI21X1 OAI21X1_1365 ( .gnd(gnd), .vdd(vdd), .A(_4881_), .B(micro_hash_ucr_2_Wx_68_), .C(_4713_), .Y(_4882_) );
AOI21X1 AOI21X1_841 ( .gnd(gnd), .vdd(vdd), .A(_4881_), .B(micro_hash_ucr_2_Wx_68_), .C(_4882_), .Y(_4883_) );
NOR2X1 NOR2X1_808 ( .gnd(gnd), .vdd(vdd), .A(_4883_), .B(_4594__bF_buf8), .Y(_4490__180_) );
INVX2 INVX2_178 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_109_), .Y(_4884_) );
OAI21X1 OAI21X1_1366 ( .gnd(gnd), .vdd(vdd), .A(_4884_), .B(micro_hash_ucr_2_Wx_69_), .C(_4716_), .Y(_4885_) );
AOI21X1 AOI21X1_842 ( .gnd(gnd), .vdd(vdd), .A(_4884_), .B(micro_hash_ucr_2_Wx_69_), .C(_4885_), .Y(_4886_) );
NOR2X1 NOR2X1_809 ( .gnd(gnd), .vdd(vdd), .A(_4886_), .B(_4594__bF_buf7), .Y(_4490__181_) );
INVX4 INVX4_84 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_70_), .Y(_4887_) );
OAI21X1 OAI21X1_1367 ( .gnd(gnd), .vdd(vdd), .A(_4887_), .B(micro_hash_ucr_2_Wx_110_), .C(_4719_), .Y(_4888_) );
AOI21X1 AOI21X1_843 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_110_), .B(_4887_), .C(_4888_), .Y(_4889_) );
NOR2X1 NOR2X1_810 ( .gnd(gnd), .vdd(vdd), .A(_4889_), .B(_4594__bF_buf6), .Y(_4490__182_) );
INVX4 INVX4_85 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_111_), .Y(_4890_) );
OAI21X1 OAI21X1_1368 ( .gnd(gnd), .vdd(vdd), .A(_4890_), .B(micro_hash_ucr_2_Wx_71_), .C(_4723_), .Y(_4891_) );
AOI21X1 AOI21X1_844 ( .gnd(gnd), .vdd(vdd), .A(_4890_), .B(micro_hash_ucr_2_Wx_71_), .C(_4891_), .Y(_4892_) );
NOR2X1 NOR2X1_811 ( .gnd(gnd), .vdd(vdd), .A(_4892_), .B(_4594__bF_buf5), .Y(_4490__183_) );
AOI21X1 AOI21X1_845 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_80_), .B(_4754_), .C(micro_hash_ucr_2_Wx_168_), .Y(_4893_) );
OAI21X1 OAI21X1_1369 ( .gnd(gnd), .vdd(vdd), .A(_4754_), .B(micro_hash_ucr_2_Wx_80_), .C(_4893_), .Y(_4894_) );
AND2X2 AND2X2_284 ( .gnd(gnd), .vdd(vdd), .A(_4894_), .B(_4496__bF_buf7), .Y(_4490__192_) );
INVX2 INVX2_179 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_121_), .Y(_4895_) );
OAI21X1 OAI21X1_1370 ( .gnd(gnd), .vdd(vdd), .A(_4895_), .B(micro_hash_ucr_2_Wx_81_), .C(_4728_), .Y(_4896_) );
AOI21X1 AOI21X1_846 ( .gnd(gnd), .vdd(vdd), .A(_4895_), .B(micro_hash_ucr_2_Wx_81_), .C(_4896_), .Y(_4897_) );
NOR2X1 NOR2X1_812 ( .gnd(gnd), .vdd(vdd), .A(_4897_), .B(_4594__bF_buf4), .Y(_4490__193_) );
INVX4 INVX4_86 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_122_), .Y(_4898_) );
OAI21X1 OAI21X1_1371 ( .gnd(gnd), .vdd(vdd), .A(_4898_), .B(micro_hash_ucr_2_Wx_82_), .C(_4732_), .Y(_4899_) );
AOI21X1 AOI21X1_847 ( .gnd(gnd), .vdd(vdd), .A(_4898_), .B(micro_hash_ucr_2_Wx_82_), .C(_4899_), .Y(_4900_) );
NOR2X1 NOR2X1_813 ( .gnd(gnd), .vdd(vdd), .A(_4900_), .B(_4594__bF_buf3), .Y(_4490__194_) );
INVX2 INVX2_180 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_123_), .Y(_4901_) );
OAI21X1 OAI21X1_1372 ( .gnd(gnd), .vdd(vdd), .A(_4901_), .B(micro_hash_ucr_2_Wx_83_), .C(_4736_), .Y(_4902_) );
AOI21X1 AOI21X1_848 ( .gnd(gnd), .vdd(vdd), .A(_4901_), .B(micro_hash_ucr_2_Wx_83_), .C(_4902_), .Y(_4903_) );
NOR2X1 NOR2X1_814 ( .gnd(gnd), .vdd(vdd), .A(_4903_), .B(_4594__bF_buf2), .Y(_4490__195_) );
OAI21X1 OAI21X1_1373 ( .gnd(gnd), .vdd(vdd), .A(_4768_), .B(micro_hash_ucr_2_Wx_84_), .C(_4740_), .Y(_4904_) );
AOI21X1 AOI21X1_849 ( .gnd(gnd), .vdd(vdd), .A(_4768_), .B(micro_hash_ucr_2_Wx_84_), .C(_4904_), .Y(_4905_) );
NOR2X1 NOR2X1_815 ( .gnd(gnd), .vdd(vdd), .A(_4905_), .B(_4594__bF_buf1), .Y(_4490__196_) );
INVX2 INVX2_181 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_125_), .Y(_4906_) );
OAI21X1 OAI21X1_1374 ( .gnd(gnd), .vdd(vdd), .A(_4906_), .B(micro_hash_ucr_2_Wx_85_), .C(_4743_), .Y(_4907_) );
AOI21X1 AOI21X1_850 ( .gnd(gnd), .vdd(vdd), .A(_4906_), .B(micro_hash_ucr_2_Wx_85_), .C(_4907_), .Y(_4908_) );
NOR2X1 NOR2X1_816 ( .gnd(gnd), .vdd(vdd), .A(_4908_), .B(_4594__bF_buf0), .Y(_4490__197_) );
INVX4 INVX4_87 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_126_), .Y(_4909_) );
OAI21X1 OAI21X1_1375 ( .gnd(gnd), .vdd(vdd), .A(_4909_), .B(micro_hash_ucr_2_Wx_86_), .C(_4747_), .Y(_4910_) );
AOI21X1 AOI21X1_851 ( .gnd(gnd), .vdd(vdd), .A(_4909_), .B(micro_hash_ucr_2_Wx_86_), .C(_4910_), .Y(_4911_) );
NOR2X1 NOR2X1_817 ( .gnd(gnd), .vdd(vdd), .A(_4911_), .B(_4594__bF_buf12), .Y(_4490__198_) );
XNOR2X1 XNOR2X1_208 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_127_), .B(micro_hash_ucr_2_Wx_87_), .Y(_4912_) );
AOI21X1 AOI21X1_852 ( .gnd(gnd), .vdd(vdd), .A(_4751_), .B(_4912_), .C(_4594__bF_buf11), .Y(_4490__199_) );
INVX2 INVX2_182 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_112_), .Y(_4913_) );
AOI21X1 AOI21X1_853 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_72_), .B(_4913_), .C(micro_hash_ucr_2_Wx_160_), .Y(_4914_) );
OAI21X1 OAI21X1_1376 ( .gnd(gnd), .vdd(vdd), .A(_4913_), .B(micro_hash_ucr_2_Wx_72_), .C(_4914_), .Y(_4915_) );
AND2X2 AND2X2_285 ( .gnd(gnd), .vdd(vdd), .A(_4915_), .B(_4496__bF_buf6), .Y(_4490__184_) );
INVX4 INVX4_88 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_113_), .Y(_4916_) );
OAI21X1 OAI21X1_1377 ( .gnd(gnd), .vdd(vdd), .A(_4916_), .B(micro_hash_ucr_2_Wx_73_), .C(_4757_), .Y(_4917_) );
AOI21X1 AOI21X1_854 ( .gnd(gnd), .vdd(vdd), .A(_4916_), .B(micro_hash_ucr_2_Wx_73_), .C(_4917_), .Y(_4918_) );
NOR2X1 NOR2X1_818 ( .gnd(gnd), .vdd(vdd), .A(_4918_), .B(_4594__bF_buf10), .Y(_4490__185_) );
INVX4 INVX4_89 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_114_), .Y(_4919_) );
OAI21X1 OAI21X1_1378 ( .gnd(gnd), .vdd(vdd), .A(_4919_), .B(micro_hash_ucr_2_Wx_74_), .C(_4760_), .Y(_4920_) );
AOI21X1 AOI21X1_855 ( .gnd(gnd), .vdd(vdd), .A(_4919_), .B(micro_hash_ucr_2_Wx_74_), .C(_4920_), .Y(_4921_) );
NOR2X1 NOR2X1_819 ( .gnd(gnd), .vdd(vdd), .A(_4921_), .B(_4594__bF_buf9), .Y(_4490__186_) );
INVX2 INVX2_183 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_115_), .Y(_4922_) );
OAI21X1 OAI21X1_1379 ( .gnd(gnd), .vdd(vdd), .A(_4922_), .B(micro_hash_ucr_2_Wx_75_), .C(_4764_), .Y(_4923_) );
AOI21X1 AOI21X1_856 ( .gnd(gnd), .vdd(vdd), .A(_4922_), .B(micro_hash_ucr_2_Wx_75_), .C(_4923_), .Y(_4924_) );
NOR2X1 NOR2X1_820 ( .gnd(gnd), .vdd(vdd), .A(_4924_), .B(_4594__bF_buf8), .Y(_4490__187_) );
INVX2 INVX2_184 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_116_), .Y(_4925_) );
AOI21X1 AOI21X1_857 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_76_), .B(_4925_), .C(micro_hash_ucr_2_Wx_164_), .Y(_4926_) );
OAI21X1 OAI21X1_1380 ( .gnd(gnd), .vdd(vdd), .A(_4925_), .B(micro_hash_ucr_2_Wx_76_), .C(_4926_), .Y(_4927_) );
AND2X2 AND2X2_286 ( .gnd(gnd), .vdd(vdd), .A(_4927_), .B(_4496__bF_buf5), .Y(_4490__188_) );
INVX2 INVX2_185 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_117_), .Y(_4928_) );
OAI21X1 OAI21X1_1381 ( .gnd(gnd), .vdd(vdd), .A(_4928_), .B(micro_hash_ucr_2_Wx_77_), .C(_4771_), .Y(_4929_) );
AOI21X1 AOI21X1_858 ( .gnd(gnd), .vdd(vdd), .A(_4928_), .B(micro_hash_ucr_2_Wx_77_), .C(_4929_), .Y(_4930_) );
NOR2X1 NOR2X1_821 ( .gnd(gnd), .vdd(vdd), .A(_4930_), .B(_4594__bF_buf7), .Y(_4490__189_) );
INVX2 INVX2_186 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_118_), .Y(_4931_) );
OAI21X1 OAI21X1_1382 ( .gnd(gnd), .vdd(vdd), .A(_4931_), .B(micro_hash_ucr_2_Wx_78_), .C(_4774_), .Y(_4932_) );
AOI21X1 AOI21X1_859 ( .gnd(gnd), .vdd(vdd), .A(_4931_), .B(micro_hash_ucr_2_Wx_78_), .C(_4932_), .Y(_4933_) );
NOR2X1 NOR2X1_822 ( .gnd(gnd), .vdd(vdd), .A(_4933_), .B(_4594__bF_buf6), .Y(_4490__190_) );
XNOR2X1 XNOR2X1_209 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_119_), .B(micro_hash_ucr_2_Wx_79_), .Y(_4934_) );
AOI21X1 AOI21X1_860 ( .gnd(gnd), .vdd(vdd), .A(_4778_), .B(_4934_), .C(_4594__bF_buf5), .Y(_4490__191_) );
INVX2 INVX2_187 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_80_), .Y(_4935_) );
OAI21X1 OAI21X1_1383 ( .gnd(gnd), .vdd(vdd), .A(_4935_), .B(micro_hash_ucr_2_Wx_40_), .C(_4781_), .Y(_4936_) );
AOI21X1 AOI21X1_861 ( .gnd(gnd), .vdd(vdd), .A(_4935_), .B(micro_hash_ucr_2_Wx_40_), .C(_4936_), .Y(_4937_) );
NOR2X1 NOR2X1_823 ( .gnd(gnd), .vdd(vdd), .A(_4937_), .B(_4594__bF_buf4), .Y(_4490__152_) );
INVX4 INVX4_90 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_81_), .Y(_4938_) );
OAI21X1 OAI21X1_1384 ( .gnd(gnd), .vdd(vdd), .A(_4938_), .B(micro_hash_ucr_2_Wx_41_), .C(_4785_), .Y(_4939_) );
AOI21X1 AOI21X1_862 ( .gnd(gnd), .vdd(vdd), .A(_4938_), .B(micro_hash_ucr_2_Wx_41_), .C(_4939_), .Y(_4940_) );
NOR2X1 NOR2X1_824 ( .gnd(gnd), .vdd(vdd), .A(_4940_), .B(_4594__bF_buf3), .Y(_4490__153_) );
INVX2 INVX2_188 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_82_), .Y(_4941_) );
OAI21X1 OAI21X1_1385 ( .gnd(gnd), .vdd(vdd), .A(_4941_), .B(micro_hash_ucr_2_Wx_42_), .C(_4789_), .Y(_4942_) );
AOI21X1 AOI21X1_863 ( .gnd(gnd), .vdd(vdd), .A(_4941_), .B(micro_hash_ucr_2_Wx_42_), .C(_4942_), .Y(_4943_) );
NOR2X1 NOR2X1_825 ( .gnd(gnd), .vdd(vdd), .A(_4943_), .B(_4594__bF_buf2), .Y(_4490__154_) );
INVX2 INVX2_189 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_83_), .Y(_4944_) );
OAI21X1 OAI21X1_1386 ( .gnd(gnd), .vdd(vdd), .A(_4944_), .B(micro_hash_ucr_2_Wx_43_), .C(_4793_), .Y(_4945_) );
AOI21X1 AOI21X1_864 ( .gnd(gnd), .vdd(vdd), .A(_4944_), .B(micro_hash_ucr_2_Wx_43_), .C(_4945_), .Y(_4946_) );
NOR2X1 NOR2X1_826 ( .gnd(gnd), .vdd(vdd), .A(_4946_), .B(_4594__bF_buf1), .Y(_4490__155_) );
INVX2 INVX2_190 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_84_), .Y(_4947_) );
OAI21X1 OAI21X1_1387 ( .gnd(gnd), .vdd(vdd), .A(_4947_), .B(micro_hash_ucr_2_Wx_44_), .C(_4797_), .Y(_4948_) );
AOI21X1 AOI21X1_865 ( .gnd(gnd), .vdd(vdd), .A(_4947_), .B(micro_hash_ucr_2_Wx_44_), .C(_4948_), .Y(_4949_) );
NOR2X1 NOR2X1_827 ( .gnd(gnd), .vdd(vdd), .A(_4949_), .B(_4594__bF_buf0), .Y(_4490__156_) );
INVX2 INVX2_191 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_85_), .Y(_4950_) );
OAI21X1 OAI21X1_1388 ( .gnd(gnd), .vdd(vdd), .A(_4950_), .B(micro_hash_ucr_2_Wx_45_), .C(_4801_), .Y(_4951_) );
AOI21X1 AOI21X1_866 ( .gnd(gnd), .vdd(vdd), .A(_4950_), .B(micro_hash_ucr_2_Wx_45_), .C(_4951_), .Y(_4952_) );
NOR2X1 NOR2X1_828 ( .gnd(gnd), .vdd(vdd), .A(_4952_), .B(_4594__bF_buf12), .Y(_4490__157_) );
INVX4 INVX4_91 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_86_), .Y(_4953_) );
OAI21X1 OAI21X1_1389 ( .gnd(gnd), .vdd(vdd), .A(_4953_), .B(micro_hash_ucr_2_Wx_46_), .C(_4805_), .Y(_4954_) );
AOI21X1 AOI21X1_867 ( .gnd(gnd), .vdd(vdd), .A(_4953_), .B(micro_hash_ucr_2_Wx_46_), .C(_4954_), .Y(_4955_) );
NOR2X1 NOR2X1_829 ( .gnd(gnd), .vdd(vdd), .A(_4955_), .B(_4594__bF_buf11), .Y(_4490__158_) );
INVX1 INVX1_362 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_87_), .Y(_4956_) );
AOI21X1 AOI21X1_868 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_47_), .B(_4956_), .C(micro_hash_ucr_2_Wx_135_), .Y(_4957_) );
OAI21X1 OAI21X1_1390 ( .gnd(gnd), .vdd(vdd), .A(_4956_), .B(micro_hash_ucr_2_Wx_47_), .C(_4957_), .Y(_4958_) );
AND2X2 AND2X2_287 ( .gnd(gnd), .vdd(vdd), .A(_4958_), .B(_4496__bF_buf4), .Y(_4490__159_) );
OAI21X1 OAI21X1_1391 ( .gnd(gnd), .vdd(vdd), .A(_4840_), .B(micro_hash_ucr_2_Wx_56_), .C(_4811_), .Y(_4959_) );
AOI21X1 AOI21X1_869 ( .gnd(gnd), .vdd(vdd), .A(_4840_), .B(micro_hash_ucr_2_Wx_56_), .C(_4959_), .Y(_4960_) );
NOR2X1 NOR2X1_830 ( .gnd(gnd), .vdd(vdd), .A(_4960_), .B(_4594__bF_buf10), .Y(_4490__168_) );
OAI21X1 OAI21X1_1392 ( .gnd(gnd), .vdd(vdd), .A(_4843_), .B(micro_hash_ucr_2_Wx_57_), .C(_4815_), .Y(_4961_) );
AOI21X1 AOI21X1_870 ( .gnd(gnd), .vdd(vdd), .A(_4843_), .B(micro_hash_ucr_2_Wx_57_), .C(_4961_), .Y(_4962_) );
NOR2X1 NOR2X1_831 ( .gnd(gnd), .vdd(vdd), .A(_4962_), .B(_4594__bF_buf9), .Y(_4490__169_) );
OAI21X1 OAI21X1_1393 ( .gnd(gnd), .vdd(vdd), .A(_4847_), .B(micro_hash_ucr_2_Wx_58_), .C(_4819_), .Y(_4963_) );
AOI21X1 AOI21X1_871 ( .gnd(gnd), .vdd(vdd), .A(_4847_), .B(micro_hash_ucr_2_Wx_58_), .C(_4963_), .Y(_4964_) );
NOR2X1 NOR2X1_832 ( .gnd(gnd), .vdd(vdd), .A(_4964_), .B(_4594__bF_buf8), .Y(_4490__170_) );
OAI21X1 OAI21X1_1394 ( .gnd(gnd), .vdd(vdd), .A(_4851_), .B(micro_hash_ucr_2_Wx_59_), .C(_4823_), .Y(_4965_) );
AOI21X1 AOI21X1_872 ( .gnd(gnd), .vdd(vdd), .A(_4851_), .B(micro_hash_ucr_2_Wx_59_), .C(_4965_), .Y(_4966_) );
NOR2X1 NOR2X1_833 ( .gnd(gnd), .vdd(vdd), .A(_4966_), .B(_4594__bF_buf7), .Y(_4490__171_) );
OAI21X1 OAI21X1_1395 ( .gnd(gnd), .vdd(vdd), .A(_4855_), .B(micro_hash_ucr_2_Wx_60_), .C(_4827_), .Y(_4967_) );
AOI21X1 AOI21X1_873 ( .gnd(gnd), .vdd(vdd), .A(_4855_), .B(micro_hash_ucr_2_Wx_60_), .C(_4967_), .Y(_4968_) );
NOR2X1 NOR2X1_834 ( .gnd(gnd), .vdd(vdd), .A(_4968_), .B(_4594__bF_buf6), .Y(_4490__172_) );
OAI21X1 OAI21X1_1396 ( .gnd(gnd), .vdd(vdd), .A(_4858_), .B(micro_hash_ucr_2_Wx_61_), .C(_4830_), .Y(_4969_) );
AOI21X1 AOI21X1_874 ( .gnd(gnd), .vdd(vdd), .A(_4858_), .B(micro_hash_ucr_2_Wx_61_), .C(_4969_), .Y(_4970_) );
NOR2X1 NOR2X1_835 ( .gnd(gnd), .vdd(vdd), .A(_4970_), .B(_4594__bF_buf5), .Y(_4490__173_) );
OAI21X1 OAI21X1_1397 ( .gnd(gnd), .vdd(vdd), .A(_4862_), .B(micro_hash_ucr_2_Wx_62_), .C(_4833_), .Y(_4971_) );
AOI21X1 AOI21X1_875 ( .gnd(gnd), .vdd(vdd), .A(_4862_), .B(micro_hash_ucr_2_Wx_62_), .C(_4971_), .Y(_4972_) );
NOR2X1 NOR2X1_836 ( .gnd(gnd), .vdd(vdd), .A(_4972_), .B(_4594__bF_buf4), .Y(_4490__174_) );
OAI21X1 OAI21X1_1398 ( .gnd(gnd), .vdd(vdd), .A(_4866_), .B(micro_hash_ucr_2_Wx_63_), .C(_4837_), .Y(_4973_) );
AOI21X1 AOI21X1_876 ( .gnd(gnd), .vdd(vdd), .A(_4866_), .B(micro_hash_ucr_2_Wx_63_), .C(_4973_), .Y(_4974_) );
NOR2X1 NOR2X1_837 ( .gnd(gnd), .vdd(vdd), .A(_4974_), .B(_4594__bF_buf3), .Y(_4490__175_) );
INVX2 INVX2_192 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_88_), .Y(_4975_) );
INVX1 INVX1_363 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_136_), .Y(_4976_) );
OAI21X1 OAI21X1_1399 ( .gnd(gnd), .vdd(vdd), .A(_4975_), .B(micro_hash_ucr_2_Wx_48_), .C(_4976_), .Y(_4977_) );
AOI21X1 AOI21X1_877 ( .gnd(gnd), .vdd(vdd), .A(_4975_), .B(micro_hash_ucr_2_Wx_48_), .C(_4977_), .Y(_4978_) );
NOR2X1 NOR2X1_838 ( .gnd(gnd), .vdd(vdd), .A(_4978_), .B(_4594__bF_buf2), .Y(_4490__160_) );
INVX2 INVX2_193 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_89_), .Y(_4979_) );
INVX2 INVX2_194 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_137_), .Y(_4980_) );
OAI21X1 OAI21X1_1400 ( .gnd(gnd), .vdd(vdd), .A(_4979_), .B(micro_hash_ucr_2_Wx_49_), .C(_4980_), .Y(_4981_) );
AOI21X1 AOI21X1_878 ( .gnd(gnd), .vdd(vdd), .A(_4979_), .B(micro_hash_ucr_2_Wx_49_), .C(_4981_), .Y(_4982_) );
NOR2X1 NOR2X1_839 ( .gnd(gnd), .vdd(vdd), .A(_4982_), .B(_4594__bF_buf1), .Y(_4490__161_) );
INVX4 INVX4_92 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_90_), .Y(_4983_) );
INVX2 INVX2_195 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_138_), .Y(_4984_) );
OAI21X1 OAI21X1_1401 ( .gnd(gnd), .vdd(vdd), .A(_4983_), .B(micro_hash_ucr_2_Wx_50_), .C(_4984_), .Y(_4985_) );
AOI21X1 AOI21X1_879 ( .gnd(gnd), .vdd(vdd), .A(_4983_), .B(micro_hash_ucr_2_Wx_50_), .C(_4985_), .Y(_4986_) );
NOR2X1 NOR2X1_840 ( .gnd(gnd), .vdd(vdd), .A(_4986_), .B(_4594__bF_buf0), .Y(_4490__162_) );
INVX2 INVX2_196 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_91_), .Y(_4987_) );
INVX1 INVX1_364 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_139_), .Y(_4988_) );
OAI21X1 OAI21X1_1402 ( .gnd(gnd), .vdd(vdd), .A(_4987_), .B(micro_hash_ucr_2_Wx_51_), .C(_4988_), .Y(_4989_) );
AOI21X1 AOI21X1_880 ( .gnd(gnd), .vdd(vdd), .A(_4987_), .B(micro_hash_ucr_2_Wx_51_), .C(_4989_), .Y(_4990_) );
NOR2X1 NOR2X1_841 ( .gnd(gnd), .vdd(vdd), .A(_4990_), .B(_4594__bF_buf12), .Y(_4490__163_) );
INVX2 INVX2_197 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_92_), .Y(_4991_) );
AOI21X1 AOI21X1_881 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_52_), .B(_4991_), .C(micro_hash_ucr_2_Wx_140_), .Y(_4992_) );
OAI21X1 OAI21X1_1403 ( .gnd(gnd), .vdd(vdd), .A(_4991_), .B(micro_hash_ucr_2_Wx_52_), .C(_4992_), .Y(_4993_) );
AND2X2 AND2X2_288 ( .gnd(gnd), .vdd(vdd), .A(_4993_), .B(_4496__bF_buf3), .Y(_4490__164_) );
INVX2 INVX2_198 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_93_), .Y(_4994_) );
INVX1 INVX1_365 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_141_), .Y(_4995_) );
OAI21X1 OAI21X1_1404 ( .gnd(gnd), .vdd(vdd), .A(_4994_), .B(micro_hash_ucr_2_Wx_53_), .C(_4995_), .Y(_4996_) );
AOI21X1 AOI21X1_882 ( .gnd(gnd), .vdd(vdd), .A(_4994_), .B(micro_hash_ucr_2_Wx_53_), .C(_4996_), .Y(_4997_) );
NOR2X1 NOR2X1_842 ( .gnd(gnd), .vdd(vdd), .A(_4997_), .B(_4594__bF_buf11), .Y(_4490__165_) );
INVX4 INVX4_93 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_94_), .Y(_4998_) );
INVX2 INVX2_199 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_142_), .Y(_4999_) );
OAI21X1 OAI21X1_1405 ( .gnd(gnd), .vdd(vdd), .A(_4998_), .B(micro_hash_ucr_2_Wx_54_), .C(_4999_), .Y(_5000_) );
AOI21X1 AOI21X1_883 ( .gnd(gnd), .vdd(vdd), .A(_4998_), .B(micro_hash_ucr_2_Wx_54_), .C(_5000_), .Y(_5001_) );
NOR2X1 NOR2X1_843 ( .gnd(gnd), .vdd(vdd), .A(_5001_), .B(_4594__bF_buf10), .Y(_4490__166_) );
INVX1 INVX1_366 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_143_), .Y(_5002_) );
XNOR2X1 XNOR2X1_210 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_95_), .B(micro_hash_ucr_2_Wx_55_), .Y(_5003_) );
AOI21X1 AOI21X1_884 ( .gnd(gnd), .vdd(vdd), .A(_5002_), .B(_5003_), .C(_4594__bF_buf9), .Y(_4490__167_) );
INVX2 INVX2_200 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_56_), .Y(_5004_) );
OAI21X1 OAI21X1_1406 ( .gnd(gnd), .vdd(vdd), .A(_5004_), .B(micro_hash_ucr_2_Wx_16_), .C(_4869_), .Y(_5005_) );
AOI21X1 AOI21X1_885 ( .gnd(gnd), .vdd(vdd), .A(_5004_), .B(micro_hash_ucr_2_Wx_16_), .C(_5005_), .Y(_5006_) );
NOR2X1 NOR2X1_844 ( .gnd(gnd), .vdd(vdd), .A(_5006_), .B(_4594__bF_buf8), .Y(_4490__128_) );
INVX2 INVX2_201 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_57_), .Y(_5007_) );
OAI21X1 OAI21X1_1407 ( .gnd(gnd), .vdd(vdd), .A(_5007_), .B(micro_hash_ucr_2_Wx_17_), .C(_4872_), .Y(_5008_) );
AOI21X1 AOI21X1_886 ( .gnd(gnd), .vdd(vdd), .A(_5007_), .B(micro_hash_ucr_2_Wx_17_), .C(_5008_), .Y(_5009_) );
NOR2X1 NOR2X1_845 ( .gnd(gnd), .vdd(vdd), .A(_5009_), .B(_4594__bF_buf7), .Y(_4490__129_) );
INVX4 INVX4_94 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_58_), .Y(_5010_) );
OAI21X1 OAI21X1_1408 ( .gnd(gnd), .vdd(vdd), .A(_5010_), .B(micro_hash_ucr_2_Wx_18_), .C(_4875_), .Y(_5011_) );
AOI21X1 AOI21X1_887 ( .gnd(gnd), .vdd(vdd), .A(_5010_), .B(micro_hash_ucr_2_Wx_18_), .C(_5011_), .Y(_5012_) );
NOR2X1 NOR2X1_846 ( .gnd(gnd), .vdd(vdd), .A(_5012_), .B(_4594__bF_buf6), .Y(_4490__130_) );
INVX2 INVX2_202 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_59_), .Y(_5013_) );
OAI21X1 OAI21X1_1409 ( .gnd(gnd), .vdd(vdd), .A(_5013_), .B(micro_hash_ucr_2_Wx_19_), .C(_4878_), .Y(_5014_) );
AOI21X1 AOI21X1_888 ( .gnd(gnd), .vdd(vdd), .A(_5013_), .B(micro_hash_ucr_2_Wx_19_), .C(_5014_), .Y(_5015_) );
NOR2X1 NOR2X1_847 ( .gnd(gnd), .vdd(vdd), .A(_5015_), .B(_4594__bF_buf5), .Y(_4490__131_) );
INVX2 INVX2_203 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_60_), .Y(_5016_) );
OAI21X1 OAI21X1_1410 ( .gnd(gnd), .vdd(vdd), .A(_5016_), .B(micro_hash_ucr_2_Wx_20_), .C(_4881_), .Y(_5017_) );
AOI21X1 AOI21X1_889 ( .gnd(gnd), .vdd(vdd), .A(_5016_), .B(micro_hash_ucr_2_Wx_20_), .C(_5017_), .Y(_5018_) );
NOR2X1 NOR2X1_848 ( .gnd(gnd), .vdd(vdd), .A(_5018_), .B(_4594__bF_buf4), .Y(_4490__132_) );
INVX2 INVX2_204 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_61_), .Y(_5019_) );
OAI21X1 OAI21X1_1411 ( .gnd(gnd), .vdd(vdd), .A(_5019_), .B(micro_hash_ucr_2_Wx_21_), .C(_4884_), .Y(_5020_) );
AOI21X1 AOI21X1_890 ( .gnd(gnd), .vdd(vdd), .A(_5019_), .B(micro_hash_ucr_2_Wx_21_), .C(_5020_), .Y(_5021_) );
NOR2X1 NOR2X1_849 ( .gnd(gnd), .vdd(vdd), .A(_5021_), .B(_4594__bF_buf3), .Y(_4490__133_) );
INVX4 INVX4_95 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_62_), .Y(_5022_) );
AOI21X1 AOI21X1_891 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_22_), .B(_5022_), .C(micro_hash_ucr_2_Wx_110_), .Y(_5023_) );
OAI21X1 OAI21X1_1412 ( .gnd(gnd), .vdd(vdd), .A(_5022_), .B(micro_hash_ucr_2_Wx_22_), .C(_5023_), .Y(_5024_) );
AND2X2 AND2X2_289 ( .gnd(gnd), .vdd(vdd), .A(_5024_), .B(_4496__bF_buf2), .Y(_4490__134_) );
XNOR2X1 XNOR2X1_211 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_63_), .B(micro_hash_ucr_2_Wx_23_), .Y(_5025_) );
AOI21X1 AOI21X1_892 ( .gnd(gnd), .vdd(vdd), .A(_4890_), .B(_5025_), .C(_4594__bF_buf2), .Y(_4490__135_) );
INVX2 INVX2_205 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_72_), .Y(_5026_) );
OAI21X1 OAI21X1_1413 ( .gnd(gnd), .vdd(vdd), .A(_5026_), .B(micro_hash_ucr_2_Wx_32_), .C(_4754_), .Y(_5027_) );
AOI21X1 AOI21X1_893 ( .gnd(gnd), .vdd(vdd), .A(_5026_), .B(micro_hash_ucr_2_Wx_32_), .C(_5027_), .Y(_5028_) );
NOR2X1 NOR2X1_850 ( .gnd(gnd), .vdd(vdd), .A(_5028_), .B(_4594__bF_buf1), .Y(_4490__144_) );
INVX2 INVX2_206 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_73_), .Y(_5029_) );
OAI21X1 OAI21X1_1414 ( .gnd(gnd), .vdd(vdd), .A(_5029_), .B(micro_hash_ucr_2_Wx_33_), .C(_4895_), .Y(_5030_) );
AOI21X1 AOI21X1_894 ( .gnd(gnd), .vdd(vdd), .A(_5029_), .B(micro_hash_ucr_2_Wx_33_), .C(_5030_), .Y(_5031_) );
NOR2X1 NOR2X1_851 ( .gnd(gnd), .vdd(vdd), .A(_5031_), .B(_4594__bF_buf0), .Y(_4490__145_) );
INVX2 INVX2_207 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_74_), .Y(_5032_) );
OAI21X1 OAI21X1_1415 ( .gnd(gnd), .vdd(vdd), .A(_5032_), .B(micro_hash_ucr_2_Wx_34_), .C(_4898_), .Y(_5033_) );
AOI21X1 AOI21X1_895 ( .gnd(gnd), .vdd(vdd), .A(_5032_), .B(micro_hash_ucr_2_Wx_34_), .C(_5033_), .Y(_5034_) );
NOR2X1 NOR2X1_852 ( .gnd(gnd), .vdd(vdd), .A(_5034_), .B(_4594__bF_buf12), .Y(_4490__146_) );
INVX2 INVX2_208 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_75_), .Y(_5035_) );
OAI21X1 OAI21X1_1416 ( .gnd(gnd), .vdd(vdd), .A(_5035_), .B(micro_hash_ucr_2_Wx_35_), .C(_4901_), .Y(_5036_) );
AOI21X1 AOI21X1_896 ( .gnd(gnd), .vdd(vdd), .A(_5035_), .B(micro_hash_ucr_2_Wx_35_), .C(_5036_), .Y(_5037_) );
NOR2X1 NOR2X1_853 ( .gnd(gnd), .vdd(vdd), .A(_5037_), .B(_4594__bF_buf11), .Y(_4490__147_) );
INVX2 INVX2_209 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_76_), .Y(_5038_) );
OAI21X1 OAI21X1_1417 ( .gnd(gnd), .vdd(vdd), .A(_5038_), .B(micro_hash_ucr_2_Wx_36_), .C(_4768_), .Y(_5039_) );
AOI21X1 AOI21X1_897 ( .gnd(gnd), .vdd(vdd), .A(_5038_), .B(micro_hash_ucr_2_Wx_36_), .C(_5039_), .Y(_5040_) );
NOR2X1 NOR2X1_854 ( .gnd(gnd), .vdd(vdd), .A(_5040_), .B(_4594__bF_buf10), .Y(_4490__148_) );
INVX2 INVX2_210 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_77_), .Y(_5041_) );
OAI21X1 OAI21X1_1418 ( .gnd(gnd), .vdd(vdd), .A(_5041_), .B(micro_hash_ucr_2_Wx_37_), .C(_4906_), .Y(_5042_) );
AOI21X1 AOI21X1_898 ( .gnd(gnd), .vdd(vdd), .A(_5041_), .B(micro_hash_ucr_2_Wx_37_), .C(_5042_), .Y(_5043_) );
NOR2X1 NOR2X1_855 ( .gnd(gnd), .vdd(vdd), .A(_5043_), .B(_4594__bF_buf9), .Y(_4490__149_) );
INVX4 INVX4_96 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_78_), .Y(_5044_) );
OAI21X1 OAI21X1_1419 ( .gnd(gnd), .vdd(vdd), .A(_5044_), .B(micro_hash_ucr_2_Wx_38_), .C(_4909_), .Y(_5045_) );
AOI21X1 AOI21X1_899 ( .gnd(gnd), .vdd(vdd), .A(_5044_), .B(micro_hash_ucr_2_Wx_38_), .C(_5045_), .Y(_5046_) );
NOR2X1 NOR2X1_856 ( .gnd(gnd), .vdd(vdd), .A(_5046_), .B(_4594__bF_buf8), .Y(_4490__150_) );
INVX2 INVX2_211 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_79_), .Y(_5047_) );
AOI21X1 AOI21X1_900 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_39_), .B(_5047_), .C(micro_hash_ucr_2_Wx_127_), .Y(_5048_) );
OAI21X1 OAI21X1_1420 ( .gnd(gnd), .vdd(vdd), .A(_5047_), .B(micro_hash_ucr_2_Wx_39_), .C(_5048_), .Y(_5049_) );
AND2X2 AND2X2_290 ( .gnd(gnd), .vdd(vdd), .A(_5049_), .B(_4496__bF_buf1), .Y(_4490__151_) );
INVX2 INVX2_212 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_64_), .Y(_5050_) );
OAI21X1 OAI21X1_1421 ( .gnd(gnd), .vdd(vdd), .A(_5050_), .B(micro_hash_ucr_2_Wx_24_), .C(_4913_), .Y(_5051_) );
AOI21X1 AOI21X1_901 ( .gnd(gnd), .vdd(vdd), .A(_5050_), .B(micro_hash_ucr_2_Wx_24_), .C(_5051_), .Y(_5052_) );
NOR2X1 NOR2X1_857 ( .gnd(gnd), .vdd(vdd), .A(_5052_), .B(_4594__bF_buf7), .Y(_4490__136_) );
INVX2 INVX2_213 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_65_), .Y(_5053_) );
OAI21X1 OAI21X1_1422 ( .gnd(gnd), .vdd(vdd), .A(_5053_), .B(micro_hash_ucr_2_Wx_25_), .C(_4916_), .Y(_5054_) );
AOI21X1 AOI21X1_902 ( .gnd(gnd), .vdd(vdd), .A(_5053_), .B(micro_hash_ucr_2_Wx_25_), .C(_5054_), .Y(_5055_) );
NOR2X1 NOR2X1_858 ( .gnd(gnd), .vdd(vdd), .A(_5055_), .B(_4594__bF_buf6), .Y(_4490__137_) );
INVX4 INVX4_97 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_66_), .Y(_5056_) );
OAI21X1 OAI21X1_1423 ( .gnd(gnd), .vdd(vdd), .A(_5056_), .B(micro_hash_ucr_2_Wx_26_), .C(_4919_), .Y(_5057_) );
AOI21X1 AOI21X1_903 ( .gnd(gnd), .vdd(vdd), .A(_5056_), .B(micro_hash_ucr_2_Wx_26_), .C(_5057_), .Y(_5058_) );
NOR2X1 NOR2X1_859 ( .gnd(gnd), .vdd(vdd), .A(_5058_), .B(_4594__bF_buf5), .Y(_4490__138_) );
INVX2 INVX2_214 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_67_), .Y(_5059_) );
OAI21X1 OAI21X1_1424 ( .gnd(gnd), .vdd(vdd), .A(_5059_), .B(micro_hash_ucr_2_Wx_27_), .C(_4922_), .Y(_5060_) );
AOI21X1 AOI21X1_904 ( .gnd(gnd), .vdd(vdd), .A(_5059_), .B(micro_hash_ucr_2_Wx_27_), .C(_5060_), .Y(_5061_) );
NOR2X1 NOR2X1_860 ( .gnd(gnd), .vdd(vdd), .A(_5061_), .B(_4594__bF_buf4), .Y(_4490__139_) );
INVX2 INVX2_215 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_68_), .Y(_5062_) );
OAI21X1 OAI21X1_1425 ( .gnd(gnd), .vdd(vdd), .A(_5062_), .B(micro_hash_ucr_2_Wx_28_), .C(_4925_), .Y(_5063_) );
AOI21X1 AOI21X1_905 ( .gnd(gnd), .vdd(vdd), .A(_5062_), .B(micro_hash_ucr_2_Wx_28_), .C(_5063_), .Y(_5064_) );
NOR2X1 NOR2X1_861 ( .gnd(gnd), .vdd(vdd), .A(_5064_), .B(_4594__bF_buf3), .Y(_4490__140_) );
INVX2 INVX2_216 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_69_), .Y(_5065_) );
OAI21X1 OAI21X1_1426 ( .gnd(gnd), .vdd(vdd), .A(_5065_), .B(micro_hash_ucr_2_Wx_29_), .C(_4928_), .Y(_5066_) );
AOI21X1 AOI21X1_906 ( .gnd(gnd), .vdd(vdd), .A(_5065_), .B(micro_hash_ucr_2_Wx_29_), .C(_5066_), .Y(_5067_) );
NOR2X1 NOR2X1_862 ( .gnd(gnd), .vdd(vdd), .A(_5067_), .B(_4594__bF_buf2), .Y(_4490__141_) );
OAI21X1 OAI21X1_1427 ( .gnd(gnd), .vdd(vdd), .A(_4887_), .B(micro_hash_ucr_2_Wx_30_), .C(_4931_), .Y(_5068_) );
AOI21X1 AOI21X1_907 ( .gnd(gnd), .vdd(vdd), .A(_4887_), .B(micro_hash_ucr_2_Wx_30_), .C(_5068_), .Y(_5069_) );
NOR2X1 NOR2X1_863 ( .gnd(gnd), .vdd(vdd), .A(_5069_), .B(_4594__bF_buf1), .Y(_4490__142_) );
INVX1 INVX1_367 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_71_), .Y(_5070_) );
AOI21X1 AOI21X1_908 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_31_), .B(_5070_), .C(micro_hash_ucr_2_Wx_119_), .Y(_5071_) );
OAI21X1 OAI21X1_1428 ( .gnd(gnd), .vdd(vdd), .A(_5070_), .B(micro_hash_ucr_2_Wx_31_), .C(_5071_), .Y(_5072_) );
AND2X2 AND2X2_291 ( .gnd(gnd), .vdd(vdd), .A(_5072_), .B(_4496__bF_buf0), .Y(_4490__143_) );
AND2X2 AND2X2_292 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf13), .B(concatenador_2_data_out_104_), .Y(_4490__104_) );
AND2X2 AND2X2_293 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf12), .B(concatenador_2_data_out_105_), .Y(_4490__105_) );
AND2X2 AND2X2_294 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf11), .B(concatenador_2_data_out_106_), .Y(_4490__106_) );
AND2X2 AND2X2_295 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf10), .B(concatenador_2_data_out_107_), .Y(_4490__107_) );
AND2X2 AND2X2_296 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf9), .B(concatenador_2_data_out_108_), .Y(_4490__108_) );
AND2X2 AND2X2_297 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf8), .B(concatenador_2_data_out_109_), .Y(_4490__109_) );
AND2X2 AND2X2_298 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf7), .B(concatenador_2_data_out_110_), .Y(_4490__110_) );
AND2X2 AND2X2_299 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf6), .B(concatenador_2_data_out_111_), .Y(_4490__111_) );
AND2X2 AND2X2_300 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf5), .B(concatenador_2_data_out_120_), .Y(_4490__120_) );
AND2X2 AND2X2_301 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf4), .B(concatenador_2_data_out_121_), .Y(_4490__121_) );
AND2X2 AND2X2_302 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf3), .B(concatenador_2_data_out_122_), .Y(_4490__122_) );
AND2X2 AND2X2_303 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf2), .B(concatenador_2_data_out_123_), .Y(_4490__123_) );
AND2X2 AND2X2_304 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf1), .B(concatenador_2_data_out_124_), .Y(_4490__124_) );
AND2X2 AND2X2_305 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf0), .B(concatenador_2_data_out_125_), .Y(_4490__125_) );
AND2X2 AND2X2_306 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf13), .B(concatenador_2_data_out_126_), .Y(_4490__126_) );
AND2X2 AND2X2_307 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf12), .B(concatenador_2_data_out_127_), .Y(_4490__127_) );
AND2X2 AND2X2_308 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf11), .B(concatenador_2_data_out_112_), .Y(_4490__112_) );
AND2X2 AND2X2_309 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf10), .B(concatenador_2_data_out_113_), .Y(_4490__113_) );
AND2X2 AND2X2_310 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf9), .B(concatenador_2_data_out_114_), .Y(_4490__114_) );
AND2X2 AND2X2_311 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf8), .B(concatenador_2_data_out_115_), .Y(_4490__115_) );
AND2X2 AND2X2_312 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf7), .B(concatenador_2_data_out_116_), .Y(_4490__116_) );
AND2X2 AND2X2_313 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf6), .B(concatenador_2_data_out_117_), .Y(_4490__117_) );
AND2X2 AND2X2_314 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf5), .B(concatenador_2_data_out_118_), .Y(_4490__118_) );
AND2X2 AND2X2_315 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf4), .B(concatenador_2_data_out_119_), .Y(_4490__119_) );
AND2X2 AND2X2_316 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf3), .B(concatenador_2_data_out_80_), .Y(_4490__80_) );
AND2X2 AND2X2_317 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf2), .B(concatenador_2_data_out_81_), .Y(_4490__81_) );
AND2X2 AND2X2_318 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf1), .B(concatenador_2_data_out_82_), .Y(_4490__82_) );
AND2X2 AND2X2_319 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf0), .B(concatenador_2_data_out_83_), .Y(_4490__83_) );
AND2X2 AND2X2_320 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf13), .B(concatenador_2_data_out_84_), .Y(_4490__84_) );
AND2X2 AND2X2_321 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf12), .B(concatenador_2_data_out_85_), .Y(_4490__85_) );
AND2X2 AND2X2_322 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf11), .B(concatenador_2_data_out_86_), .Y(_4490__86_) );
AND2X2 AND2X2_323 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf10), .B(concatenador_2_data_out_87_), .Y(_4490__87_) );
AND2X2 AND2X2_324 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf9), .B(concatenador_2_data_out_96_), .Y(_4490__96_) );
AND2X2 AND2X2_325 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf8), .B(concatenador_2_data_out_97_), .Y(_4490__97_) );
AND2X2 AND2X2_326 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf7), .B(concatenador_2_data_out_98_), .Y(_4490__98_) );
AND2X2 AND2X2_327 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf6), .B(concatenador_2_data_out_99_), .Y(_4490__99_) );
AND2X2 AND2X2_328 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf5), .B(concatenador_2_data_out_100_), .Y(_4490__100_) );
AND2X2 AND2X2_329 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf4), .B(concatenador_2_data_out_101_), .Y(_4490__101_) );
AND2X2 AND2X2_330 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf3), .B(concatenador_2_data_out_102_), .Y(_4490__102_) );
AND2X2 AND2X2_331 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf2), .B(concatenador_2_data_out_103_), .Y(_4490__103_) );
AND2X2 AND2X2_332 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf1), .B(concatenador_2_data_out_88_), .Y(_4490__88_) );
AND2X2 AND2X2_333 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf0), .B(concatenador_2_data_out_89_), .Y(_4490__89_) );
AND2X2 AND2X2_334 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf13), .B(concatenador_2_data_out_90_), .Y(_4490__90_) );
AND2X2 AND2X2_335 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf12), .B(concatenador_2_data_out_91_), .Y(_4490__91_) );
AND2X2 AND2X2_336 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf11), .B(concatenador_2_data_out_92_), .Y(_4490__92_) );
AND2X2 AND2X2_337 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf10), .B(concatenador_2_data_out_93_), .Y(_4490__93_) );
AND2X2 AND2X2_338 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf9), .B(concatenador_2_data_out_94_), .Y(_4490__94_) );
AND2X2 AND2X2_339 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf8), .B(concatenador_2_data_out_95_), .Y(_4490__95_) );
AND2X2 AND2X2_340 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf7), .B(concatenador_2_data_out_56_), .Y(_4490__56_) );
AND2X2 AND2X2_341 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf6), .B(concatenador_2_data_out_57_), .Y(_4490__57_) );
AND2X2 AND2X2_342 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf5), .B(concatenador_2_data_out_58_), .Y(_4490__58_) );
AND2X2 AND2X2_343 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf4), .B(concatenador_2_data_out_59_), .Y(_4490__59_) );
AND2X2 AND2X2_344 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf3), .B(concatenador_2_data_out_60_), .Y(_4490__60_) );
AND2X2 AND2X2_345 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf2), .B(concatenador_2_data_out_61_), .Y(_4490__61_) );
AND2X2 AND2X2_346 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf1), .B(concatenador_2_data_out_62_), .Y(_4490__62_) );
AND2X2 AND2X2_347 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf0), .B(concatenador_2_data_out_63_), .Y(_4490__63_) );
AND2X2 AND2X2_348 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf13), .B(concatenador_2_data_out_72_), .Y(_4490__72_) );
AND2X2 AND2X2_349 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf12), .B(concatenador_2_data_out_73_), .Y(_4490__73_) );
AND2X2 AND2X2_350 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf11), .B(concatenador_2_data_out_74_), .Y(_4490__74_) );
AND2X2 AND2X2_351 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf10), .B(concatenador_2_data_out_75_), .Y(_4490__75_) );
AND2X2 AND2X2_352 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf9), .B(concatenador_2_data_out_76_), .Y(_4490__76_) );
AND2X2 AND2X2_353 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf8), .B(concatenador_2_data_out_77_), .Y(_4490__77_) );
AND2X2 AND2X2_354 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf7), .B(concatenador_2_data_out_78_), .Y(_4490__78_) );
AND2X2 AND2X2_355 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf6), .B(concatenador_2_data_out_79_), .Y(_4490__79_) );
AND2X2 AND2X2_356 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf5), .B(concatenador_2_data_out_64_), .Y(_4490__64_) );
AND2X2 AND2X2_357 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf4), .B(concatenador_2_data_out_65_), .Y(_4490__65_) );
AND2X2 AND2X2_358 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf3), .B(concatenador_2_data_out_66_), .Y(_4490__66_) );
AND2X2 AND2X2_359 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf2), .B(concatenador_2_data_out_67_), .Y(_4490__67_) );
AND2X2 AND2X2_360 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf1), .B(concatenador_2_data_out_68_), .Y(_4490__68_) );
AND2X2 AND2X2_361 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf0), .B(concatenador_2_data_out_69_), .Y(_4490__69_) );
AND2X2 AND2X2_362 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf13), .B(concatenador_2_data_out_70_), .Y(_4490__70_) );
AND2X2 AND2X2_363 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf12), .B(concatenador_2_data_out_71_), .Y(_4490__71_) );
AND2X2 AND2X2_364 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf11), .B(concatenador_2_data_out_32_), .Y(_4490__32_) );
AND2X2 AND2X2_365 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf10), .B(concatenador_2_data_out_33_), .Y(_4490__33_) );
AND2X2 AND2X2_366 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf9), .B(concatenador_2_data_out_34_), .Y(_4490__34_) );
AND2X2 AND2X2_367 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf8), .B(concatenador_2_data_out_35_), .Y(_4490__35_) );
AND2X2 AND2X2_368 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf7), .B(concatenador_2_data_out_36_), .Y(_4490__36_) );
AND2X2 AND2X2_369 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf6), .B(concatenador_2_data_out_37_), .Y(_4490__37_) );
AND2X2 AND2X2_370 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf5), .B(concatenador_2_data_out_38_), .Y(_4490__38_) );
AND2X2 AND2X2_371 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf4), .B(concatenador_2_data_out_39_), .Y(_4490__39_) );
AND2X2 AND2X2_372 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf3), .B(concatenador_2_data_out_48_), .Y(_4490__48_) );
AND2X2 AND2X2_373 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf2), .B(concatenador_2_data_out_49_), .Y(_4490__49_) );
AND2X2 AND2X2_374 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf1), .B(concatenador_2_data_out_50_), .Y(_4490__50_) );
AND2X2 AND2X2_375 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf0), .B(concatenador_2_data_out_51_), .Y(_4490__51_) );
AND2X2 AND2X2_376 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf13), .B(concatenador_2_data_out_52_), .Y(_4490__52_) );
AND2X2 AND2X2_377 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf12), .B(concatenador_2_data_out_53_), .Y(_4490__53_) );
AND2X2 AND2X2_378 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf11), .B(concatenador_2_data_out_54_), .Y(_4490__54_) );
AND2X2 AND2X2_379 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf10), .B(concatenador_2_data_out_55_), .Y(_4490__55_) );
AND2X2 AND2X2_380 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf9), .B(concatenador_2_data_out_40_), .Y(_4490__40_) );
AND2X2 AND2X2_381 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf8), .B(concatenador_2_data_out_41_), .Y(_4490__41_) );
AND2X2 AND2X2_382 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf7), .B(concatenador_2_data_out_42_), .Y(_4490__42_) );
AND2X2 AND2X2_383 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf6), .B(concatenador_2_data_out_43_), .Y(_4490__43_) );
AND2X2 AND2X2_384 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf5), .B(concatenador_2_data_out_44_), .Y(_4490__44_) );
AND2X2 AND2X2_385 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf4), .B(concatenador_2_data_out_45_), .Y(_4490__45_) );
AND2X2 AND2X2_386 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf3), .B(concatenador_2_data_out_46_), .Y(_4490__46_) );
AND2X2 AND2X2_387 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf2), .B(concatenador_2_data_out_47_), .Y(_4490__47_) );
AND2X2 AND2X2_388 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf1), .B(concatenador_2_data_out_8_), .Y(_4490__8_) );
AND2X2 AND2X2_389 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf0), .B(concatenador_2_data_out_9_), .Y(_4490__9_) );
AND2X2 AND2X2_390 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf13), .B(concatenador_2_data_out_10_), .Y(_4490__10_) );
AND2X2 AND2X2_391 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf12), .B(concatenador_2_data_out_11_), .Y(_4490__11_) );
AND2X2 AND2X2_392 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf11), .B(concatenador_2_data_out_12_), .Y(_4490__12_) );
AND2X2 AND2X2_393 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf10), .B(concatenador_2_data_out_13_), .Y(_4490__13_) );
AND2X2 AND2X2_394 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf9), .B(concatenador_2_data_out_14_), .Y(_4490__14_) );
AND2X2 AND2X2_395 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf8), .B(concatenador_2_data_out_15_), .Y(_4490__15_) );
AND2X2 AND2X2_396 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf7), .B(concatenador_2_data_out_24_), .Y(_4490__24_) );
AND2X2 AND2X2_397 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf6), .B(concatenador_2_data_out_25_), .Y(_4490__25_) );
AND2X2 AND2X2_398 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf5), .B(concatenador_2_data_out_26_), .Y(_4490__26_) );
AND2X2 AND2X2_399 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf4), .B(concatenador_2_data_out_27_), .Y(_4490__27_) );
AND2X2 AND2X2_400 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf3), .B(concatenador_2_data_out_28_), .Y(_4490__28_) );
AND2X2 AND2X2_401 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf2), .B(concatenador_2_data_out_29_), .Y(_4490__29_) );
AND2X2 AND2X2_402 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf1), .B(concatenador_2_data_out_30_), .Y(_4490__30_) );
AND2X2 AND2X2_403 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf0), .B(concatenador_2_data_out_31_), .Y(_4490__31_) );
AND2X2 AND2X2_404 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf13), .B(concatenador_2_data_out_16_), .Y(_4490__16_) );
AND2X2 AND2X2_405 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf12), .B(concatenador_2_data_out_17_), .Y(_4490__17_) );
AND2X2 AND2X2_406 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf11), .B(concatenador_2_data_out_18_), .Y(_4490__18_) );
AND2X2 AND2X2_407 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf10), .B(concatenador_2_data_out_19_), .Y(_4490__19_) );
AND2X2 AND2X2_408 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf9), .B(concatenador_2_data_out_20_), .Y(_4490__20_) );
AND2X2 AND2X2_409 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf8), .B(concatenador_2_data_out_21_), .Y(_4490__21_) );
AND2X2 AND2X2_410 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf7), .B(concatenador_2_data_out_22_), .Y(_4490__22_) );
AND2X2 AND2X2_411 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf6), .B(concatenador_2_data_out_23_), .Y(_4490__23_) );
INVX8 INVX8_113 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe69), .Y(_5073_) );
NOR2X1 NOR2X1_864 ( .gnd(gnd), .vdd(vdd), .A(_5073__bF_buf3), .B(_4594__bF_buf0), .Y(_4563_) );
AND2X2 AND2X2_412 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf5), .B(concatenador_2_data_out_0_), .Y(_4490__0_) );
AND2X2 AND2X2_413 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf4), .B(concatenador_2_data_out_1_), .Y(_4490__1_) );
AND2X2 AND2X2_414 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf3), .B(concatenador_2_data_out_2_), .Y(_4490__2_) );
AND2X2 AND2X2_415 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf2), .B(concatenador_2_data_out_3_), .Y(_4490__3_) );
AND2X2 AND2X2_416 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf1), .B(concatenador_2_data_out_4_), .Y(_4490__4_) );
AND2X2 AND2X2_417 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf0), .B(concatenador_2_data_out_5_), .Y(_4490__5_) );
AND2X2 AND2X2_418 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf13), .B(concatenador_2_data_out_6_), .Y(_4490__6_) );
AND2X2 AND2X2_419 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf12), .B(concatenador_2_data_out_7_), .Y(_4490__7_) );
NOR2X1 NOR2X1_865 ( .gnd(gnd), .vdd(vdd), .A(_8688__bF_buf1), .B(_4594__bF_buf12), .Y(_4564_) );
INVX8 INVX8_114 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe66_bF_buf4), .Y(_5074_) );
NOR2X1 NOR2X1_866 ( .gnd(gnd), .vdd(vdd), .A(_5074__bF_buf3), .B(_4594__bF_buf11), .Y(_4559_) );
INVX8 INVX8_115 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe68), .Y(_5075_) );
NOR2X1 NOR2X1_867 ( .gnd(gnd), .vdd(vdd), .A(_5075__bF_buf4), .B(_4594__bF_buf10), .Y(_4561_) );
INVX8 INVX8_116 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe67), .Y(_5076_) );
NOR2X1 NOR2X1_868 ( .gnd(gnd), .vdd(vdd), .A(_5076__bF_buf3), .B(_4594__bF_buf9), .Y(_4560_) );
INVX8 INVX8_117 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe63), .Y(_5077_) );
NOR2X1 NOR2X1_869 ( .gnd(gnd), .vdd(vdd), .A(_5077__bF_buf3), .B(_4594__bF_buf8), .Y(_4556_) );
INVX8 INVX8_118 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe65_bF_buf3), .Y(_5078_) );
NOR2X1 NOR2X1_870 ( .gnd(gnd), .vdd(vdd), .A(_5078_), .B(_4594__bF_buf7), .Y(_4558_) );
INVX8 INVX8_119 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe64_bF_buf4), .Y(_5079_) );
NOR2X1 NOR2X1_871 ( .gnd(gnd), .vdd(vdd), .A(_5079__bF_buf4), .B(_4594__bF_buf6), .Y(_4557_) );
INVX8 INVX8_120 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe60_bF_buf4), .Y(_5080_) );
NOR2X1 NOR2X1_872 ( .gnd(gnd), .vdd(vdd), .A(_5080__bF_buf3), .B(_4594__bF_buf5), .Y(_4553_) );
INVX8 INVX8_121 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe62_bF_buf4), .Y(_5081_) );
NOR2X1 NOR2X1_873 ( .gnd(gnd), .vdd(vdd), .A(_5081__bF_buf3), .B(_4594__bF_buf4), .Y(_4555_) );
INVX8 INVX8_122 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe61_bF_buf3), .Y(_5082_) );
NOR2X1 NOR2X1_874 ( .gnd(gnd), .vdd(vdd), .A(_5082_), .B(_4594__bF_buf3), .Y(_4554_) );
INVX8 INVX8_123 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe57_bF_buf3), .Y(_5083_) );
NOR2X1 NOR2X1_875 ( .gnd(gnd), .vdd(vdd), .A(_5083_), .B(_4594__bF_buf2), .Y(_4549_) );
INVX8 INVX8_124 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe59), .Y(_5084_) );
NOR2X1 NOR2X1_876 ( .gnd(gnd), .vdd(vdd), .A(_5084__bF_buf3), .B(_4594__bF_buf1), .Y(_4552_) );
INVX8 INVX8_125 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe58_bF_buf4), .Y(_5085_) );
NOR2X1 NOR2X1_877 ( .gnd(gnd), .vdd(vdd), .A(_5085__bF_buf3), .B(_4594__bF_buf0), .Y(_4550_) );
INVX8 INVX8_126 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe54_bF_buf4), .Y(_5086_) );
NOR2X1 NOR2X1_878 ( .gnd(gnd), .vdd(vdd), .A(_5086__bF_buf3), .B(_4594__bF_buf12), .Y(_4546_) );
INVX8 INVX8_127 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe56_bF_buf3), .Y(_5087_) );
NOR2X1 NOR2X1_879 ( .gnd(gnd), .vdd(vdd), .A(_5087__bF_buf4), .B(_4594__bF_buf11), .Y(_4548_) );
INVX8 INVX8_128 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe55), .Y(_5088_) );
NOR2X1 NOR2X1_880 ( .gnd(gnd), .vdd(vdd), .A(_5088_), .B(_4594__bF_buf10), .Y(_4547_) );
INVX8 INVX8_129 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe51), .Y(_5089_) );
NOR2X1 NOR2X1_881 ( .gnd(gnd), .vdd(vdd), .A(_5089__bF_buf3), .B(_4594__bF_buf9), .Y(_4543_) );
INVX8 INVX8_130 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe53_bF_buf3), .Y(_5090_) );
NOR2X1 NOR2X1_882 ( .gnd(gnd), .vdd(vdd), .A(_5090_), .B(_4594__bF_buf8), .Y(_4545_) );
INVX8 INVX8_131 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe52_bF_buf3), .Y(_5091_) );
NOR2X1 NOR2X1_883 ( .gnd(gnd), .vdd(vdd), .A(_5091__bF_buf4), .B(_4594__bF_buf7), .Y(_4544_) );
INVX8 INVX8_132 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe48_bF_buf4), .Y(_5092_) );
NOR2X1 NOR2X1_884 ( .gnd(gnd), .vdd(vdd), .A(_5092__bF_buf4), .B(_4594__bF_buf6), .Y(_4539_) );
INVX8 INVX8_133 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe50_bF_buf3), .Y(_5093_) );
NOR2X1 NOR2X1_885 ( .gnd(gnd), .vdd(vdd), .A(_5093__bF_buf4), .B(_4594__bF_buf5), .Y(_4542_) );
INVX8 INVX8_134 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe49_bF_buf3), .Y(_5094_) );
NOR2X1 NOR2X1_886 ( .gnd(gnd), .vdd(vdd), .A(_5094_), .B(_4594__bF_buf4), .Y(_4541_) );
INVX8 INVX8_135 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe45_bF_buf3), .Y(_5095_) );
NOR2X1 NOR2X1_887 ( .gnd(gnd), .vdd(vdd), .A(_5095_), .B(_4594__bF_buf3), .Y(_4536_) );
INVX8 INVX8_136 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe47), .Y(_5096_) );
NOR2X1 NOR2X1_888 ( .gnd(gnd), .vdd(vdd), .A(_5096__bF_buf3), .B(_4594__bF_buf2), .Y(_4538_) );
INVX8 INVX8_137 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe46_bF_buf4), .Y(_5097_) );
NOR2X1 NOR2X1_889 ( .gnd(gnd), .vdd(vdd), .A(_5097__bF_buf3), .B(_4594__bF_buf1), .Y(_4537_) );
INVX8 INVX8_138 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe42_bF_buf3), .Y(_5098_) );
NOR2X1 NOR2X1_890 ( .gnd(gnd), .vdd(vdd), .A(_5098__bF_buf4), .B(_4594__bF_buf0), .Y(_4533_) );
INVX8 INVX8_139 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe44_bF_buf3), .Y(_5099_) );
NOR2X1 NOR2X1_891 ( .gnd(gnd), .vdd(vdd), .A(_5099__bF_buf4), .B(_4594__bF_buf12), .Y(_4535_) );
INVX8 INVX8_140 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe43), .Y(_5100_) );
NOR2X1 NOR2X1_892 ( .gnd(gnd), .vdd(vdd), .A(_5100__bF_buf3), .B(_4594__bF_buf11), .Y(_4534_) );
INVX8 INVX8_141 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe39), .Y(_5101_) );
NOR2X1 NOR2X1_893 ( .gnd(gnd), .vdd(vdd), .A(_5101_), .B(_4594__bF_buf10), .Y(_4530_) );
INVX8 INVX8_142 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe41_bF_buf3), .Y(_5102_) );
NOR2X1 NOR2X1_894 ( .gnd(gnd), .vdd(vdd), .A(_5102_), .B(_4594__bF_buf9), .Y(_4532_) );
INVX8 INVX8_143 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe40_bF_buf4), .Y(_5103_) );
NOR2X1 NOR2X1_895 ( .gnd(gnd), .vdd(vdd), .A(_5103__bF_buf3), .B(_4594__bF_buf8), .Y(_4531_) );
INVX8 INVX8_144 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe36_bF_buf3), .Y(_5104_) );
NOR2X1 NOR2X1_896 ( .gnd(gnd), .vdd(vdd), .A(_5104__bF_buf4), .B(_4594__bF_buf7), .Y(_4526_) );
INVX8 INVX8_145 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe38_bF_buf3), .Y(_5105_) );
NOR2X1 NOR2X1_897 ( .gnd(gnd), .vdd(vdd), .A(_5105__bF_buf4), .B(_4594__bF_buf6), .Y(_4528_) );
INVX8 INVX8_146 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe37), .Y(_5106_) );
NOR2X1 NOR2X1_898 ( .gnd(gnd), .vdd(vdd), .A(_5106_), .B(_4594__bF_buf5), .Y(_4527_) );
INVX8 INVX8_147 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe33_bF_buf3), .Y(_5107_) );
NOR2X1 NOR2X1_899 ( .gnd(gnd), .vdd(vdd), .A(_5107_), .B(_4594__bF_buf4), .Y(_4523_) );
INVX8 INVX8_148 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe35), .Y(_5108_) );
NOR2X1 NOR2X1_900 ( .gnd(gnd), .vdd(vdd), .A(_5108__bF_buf3), .B(_4594__bF_buf3), .Y(_4525_) );
INVX8 INVX8_149 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe34_bF_buf3), .Y(_5109_) );
NOR2X1 NOR2X1_901 ( .gnd(gnd), .vdd(vdd), .A(_5109__bF_buf4), .B(_4594__bF_buf2), .Y(_4524_) );
INVX8 INVX8_150 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe30_bF_buf4), .Y(_5110_) );
NOR2X1 NOR2X1_902 ( .gnd(gnd), .vdd(vdd), .A(_5110__bF_buf3), .B(_4594__bF_buf1), .Y(_4520_) );
INVX8 INVX8_151 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe32_bF_buf3), .Y(_5111_) );
NOR2X1 NOR2X1_903 ( .gnd(gnd), .vdd(vdd), .A(_5111__bF_buf4), .B(_4594__bF_buf0), .Y(_4522_) );
INVX8 INVX8_152 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe31), .Y(_5112_) );
NOR2X1 NOR2X1_904 ( .gnd(gnd), .vdd(vdd), .A(_5112__bF_buf3), .B(_4594__bF_buf12), .Y(_4521_) );
INVX8 INVX8_153 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe27), .Y(_5113_) );
NOR2X1 NOR2X1_905 ( .gnd(gnd), .vdd(vdd), .A(_5113_), .B(_4594__bF_buf11), .Y(_4516_) );
INVX8 INVX8_154 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe29_bF_buf3), .Y(_5114_) );
NOR2X1 NOR2X1_906 ( .gnd(gnd), .vdd(vdd), .A(_5114_), .B(_4594__bF_buf10), .Y(_4519_) );
INVX8 INVX8_155 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe28_bF_buf3), .Y(_5115_) );
NOR2X1 NOR2X1_907 ( .gnd(gnd), .vdd(vdd), .A(_5115__bF_buf4), .B(_4594__bF_buf9), .Y(_4517_) );
INVX8 INVX8_156 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe24_bF_buf3), .Y(_5116_) );
NOR2X1 NOR2X1_908 ( .gnd(gnd), .vdd(vdd), .A(_5116__bF_buf4), .B(_4594__bF_buf8), .Y(_4513_) );
INVX8 INVX8_157 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe26_bF_buf3), .Y(_5117_) );
NOR2X1 NOR2X1_909 ( .gnd(gnd), .vdd(vdd), .A(_5117__bF_buf4), .B(_4594__bF_buf7), .Y(_4515_) );
INVX8 INVX8_158 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe25), .Y(_5118_) );
NOR2X1 NOR2X1_910 ( .gnd(gnd), .vdd(vdd), .A(_5118__bF_buf3), .B(_4594__bF_buf6), .Y(_4514_) );
INVX8 INVX8_159 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe21_bF_buf3), .Y(_5119_) );
NOR2X1 NOR2X1_911 ( .gnd(gnd), .vdd(vdd), .A(_5119_), .B(_4594__bF_buf5), .Y(_4510_) );
INVX8 INVX8_160 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe23), .Y(_5120_) );
NOR2X1 NOR2X1_912 ( .gnd(gnd), .vdd(vdd), .A(_5120__bF_buf3), .B(_4594__bF_buf4), .Y(_4512_) );
INVX8 INVX8_161 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe22_bF_buf4), .Y(_5121_) );
NOR2X1 NOR2X1_913 ( .gnd(gnd), .vdd(vdd), .A(_5121__bF_buf4), .B(_4594__bF_buf3), .Y(_4511_) );
INVX8 INVX8_162 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe18_bF_buf4), .Y(_5122_) );
NOR2X1 NOR2X1_914 ( .gnd(gnd), .vdd(vdd), .A(_5122__bF_buf4), .B(_4594__bF_buf2), .Y(_4506_) );
INVX8 INVX8_163 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe20_bF_buf3), .Y(_5123_) );
NOR2X1 NOR2X1_915 ( .gnd(gnd), .vdd(vdd), .A(_5123__bF_buf4), .B(_4594__bF_buf1), .Y(_4509_) );
INVX8 INVX8_164 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe19), .Y(_5124_) );
NOR2X1 NOR2X1_916 ( .gnd(gnd), .vdd(vdd), .A(_5124__bF_buf3), .B(_4594__bF_buf0), .Y(_4508_) );
INVX8 INVX8_165 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe15), .Y(_5125_) );
NOR2X1 NOR2X1_917 ( .gnd(gnd), .vdd(vdd), .A(_5125__bF_buf3), .B(_4594__bF_buf12), .Y(_4503_) );
INVX8 INVX8_166 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe17_bF_buf3), .Y(_5126_) );
NOR2X1 NOR2X1_918 ( .gnd(gnd), .vdd(vdd), .A(_5126_), .B(_4594__bF_buf11), .Y(_4505_) );
INVX8 INVX8_167 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe16_bF_buf4), .Y(_5127_) );
NOR2X1 NOR2X1_919 ( .gnd(gnd), .vdd(vdd), .A(_5127__bF_buf3), .B(_4594__bF_buf10), .Y(_4504_) );
INVX8 INVX8_168 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe12_bF_buf3), .Y(_5128_) );
NOR2X1 NOR2X1_920 ( .gnd(gnd), .vdd(vdd), .A(_5128_), .B(_4594__bF_buf9), .Y(_4500_) );
INVX8 INVX8_169 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe14_bF_buf4), .Y(_5129_) );
NOR2X1 NOR2X1_921 ( .gnd(gnd), .vdd(vdd), .A(_5129_), .B(_4594__bF_buf8), .Y(_4502_) );
INVX4 INVX4_98 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe13), .Y(_5130_) );
NOR2X1 NOR2X1_922 ( .gnd(gnd), .vdd(vdd), .A(_5130_), .B(_4594__bF_buf7), .Y(_4501_) );
INVX4 INVX4_99 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe9), .Y(_5131_) );
NOR2X1 NOR2X1_923 ( .gnd(gnd), .vdd(vdd), .A(_5131_), .B(_4594__bF_buf6), .Y(_4497_) );
INVX8 INVX8_170 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe11), .Y(_5132_) );
NOR2X1 NOR2X1_924 ( .gnd(gnd), .vdd(vdd), .A(_5132_), .B(_4594__bF_buf5), .Y(_4499_) );
INVX8 INVX8_171 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe10), .Y(_5133_) );
NOR2X1 NOR2X1_925 ( .gnd(gnd), .vdd(vdd), .A(_5133_), .B(_4594__bF_buf4), .Y(_4498_) );
INVX8 INVX8_172 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe6), .Y(_5134_) );
NOR2X1 NOR2X1_926 ( .gnd(gnd), .vdd(vdd), .A(_5134_), .B(_4594__bF_buf3), .Y(_4565_) );
INVX4 INVX4_100 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe8), .Y(_5135_) );
NOR2X1 NOR2X1_927 ( .gnd(gnd), .vdd(vdd), .A(_5135_), .B(_4594__bF_buf2), .Y(_4567_) );
INVX4 INVX4_101 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe7), .Y(_5136_) );
NOR2X1 NOR2X1_928 ( .gnd(gnd), .vdd(vdd), .A(_5136_), .B(_4594__bF_buf1), .Y(_4566_) );
AND2X2 AND2X2_420 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf11), .B(micro_hash_ucr_2_pipe3), .Y(_4540_) );
AND2X2 AND2X2_421 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf10), .B(micro_hash_ucr_2_pipe5), .Y(_4562_) );
AND2X2 AND2X2_422 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf9), .B(micro_hash_ucr_2_pipe4), .Y(_4551_) );
AND2X2 AND2X2_423 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf8), .B(micro_hash_ucr_2_pipe0), .Y(_4507_) );
AND2X2 AND2X2_424 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf7), .B(micro_hash_ucr_2_pipe2), .Y(_4529_) );
AND2X2 AND2X2_425 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf6), .B(micro_hash_ucr_2_pipe1), .Y(_4518_) );
NAND2X1 NAND2X1_592 ( .gnd(gnd), .vdd(vdd), .A(_8632__bF_buf1), .B(_8690_), .Y(_5137_) );
NAND2X1 NAND2X1_593 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_0_bF_buf1_), .B(micro_hash_ucr_2_b_0_bF_buf1_), .Y(_5138_) );
NAND2X1 NAND2X1_594 ( .gnd(gnd), .vdd(vdd), .A(_5138_), .B(_5137_), .Y(_5139_) );
NAND2X1 NAND2X1_595 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_0_), .B(micro_hash_ucr_2_pipe58_bF_buf3), .Y(_5140_) );
NAND2X1 NAND2X1_596 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_0_), .B(micro_hash_ucr_2_pipe56_bF_buf2), .Y(_5141_) );
NAND2X1 NAND2X1_597 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_0_), .B(micro_hash_ucr_2_pipe54_bF_buf3), .Y(_5142_) );
NAND2X1 NAND2X1_598 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_0_), .B(micro_hash_ucr_2_pipe52_bF_buf2), .Y(_5143_) );
NAND2X1 NAND2X1_599 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_0_), .B(micro_hash_ucr_2_pipe50_bF_buf2), .Y(_5144_) );
NAND2X1 NAND2X1_600 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_0_), .B(micro_hash_ucr_2_pipe48_bF_buf3), .Y(_5145_) );
NAND2X1 NAND2X1_601 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_0_), .B(micro_hash_ucr_2_pipe46_bF_buf3), .Y(_5146_) );
NAND2X1 NAND2X1_602 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_0_), .B(micro_hash_ucr_2_pipe44_bF_buf2), .Y(_5147_) );
INVX4 INVX4_102 ( .gnd(gnd), .vdd(vdd), .A(_5139__bF_buf3), .Y(_5148_) );
NOR2X1 NOR2X1_929 ( .gnd(gnd), .vdd(vdd), .A(_5114_), .B(_5148_), .Y(_5149_) );
NAND2X1 NAND2X1_603 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe27), .B(_5148_), .Y(_5150_) );
OAI21X1 OAI21X1_1429 ( .gnd(gnd), .vdd(vdd), .A(_5128_), .B(micro_hash_ucr_2_pipe13), .C(_5129_), .Y(_5151_) );
AOI21X1 AOI21X1_909 ( .gnd(gnd), .vdd(vdd), .A(_5125__bF_buf2), .B(_5151_), .C(micro_hash_ucr_2_pipe16_bF_buf3), .Y(_5152_) );
OAI21X1 OAI21X1_1430 ( .gnd(gnd), .vdd(vdd), .A(_5152_), .B(micro_hash_ucr_2_pipe17_bF_buf2), .C(_5122__bF_buf3), .Y(_5153_) );
AOI21X1 AOI21X1_910 ( .gnd(gnd), .vdd(vdd), .A(_5124__bF_buf2), .B(_5153_), .C(micro_hash_ucr_2_pipe20_bF_buf2), .Y(_5154_) );
OAI21X1 OAI21X1_1431 ( .gnd(gnd), .vdd(vdd), .A(_5154_), .B(micro_hash_ucr_2_pipe21_bF_buf2), .C(_5121__bF_buf3), .Y(_5155_) );
AOI21X1 AOI21X1_911 ( .gnd(gnd), .vdd(vdd), .A(_5120__bF_buf2), .B(_5155_), .C(micro_hash_ucr_2_pipe24_bF_buf2), .Y(_5156_) );
OAI21X1 OAI21X1_1432 ( .gnd(gnd), .vdd(vdd), .A(_5156_), .B(micro_hash_ucr_2_pipe25), .C(_5117__bF_buf3), .Y(_5157_) );
OAI21X1 OAI21X1_1433 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe6), .B(micro_hash_ucr_2_pipe7), .C(_5135_), .Y(_5158_) );
AOI21X1 AOI21X1_912 ( .gnd(gnd), .vdd(vdd), .A(_5131_), .B(_5158_), .C(micro_hash_ucr_2_pipe10), .Y(_5159_) );
OAI21X1 OAI21X1_1434 ( .gnd(gnd), .vdd(vdd), .A(_5159_), .B(micro_hash_ucr_2_pipe11), .C(_5128_), .Y(_5160_) );
NAND2X1 NAND2X1_604 ( .gnd(gnd), .vdd(vdd), .A(_5123__bF_buf3), .B(_5127__bF_buf2), .Y(_5161_) );
NOR2X1 NOR2X1_930 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe14_bF_buf3), .B(_5161_), .Y(_5162_) );
NOR2X1 NOR2X1_931 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe24_bF_buf1), .B(micro_hash_ucr_2_pipe26_bF_buf2), .Y(_5163_) );
NOR2X1 NOR2X1_932 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe22_bF_buf3), .B(micro_hash_ucr_2_pipe18_bF_buf3), .Y(_5164_) );
NAND3X1 NAND3X1_180 ( .gnd(gnd), .vdd(vdd), .A(_5163_), .B(_5164_), .C(_5162_), .Y(_5165_) );
OAI21X1 OAI21X1_1435 ( .gnd(gnd), .vdd(vdd), .A(_5160_), .B(_5165_), .C(_4630_), .Y(_5166_) );
NAND3X1 NAND3X1_181 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe6), .B(_5133_), .C(_5135_), .Y(_5167_) );
NOR2X1 NOR2X1_933 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe9), .B(micro_hash_ucr_2_pipe7), .Y(_5168_) );
NAND3X1 NAND3X1_182 ( .gnd(gnd), .vdd(vdd), .A(_4628_), .B(_5132_), .C(_5168_), .Y(_5169_) );
NOR2X1 NOR2X1_934 ( .gnd(gnd), .vdd(vdd), .A(_5167_), .B(_5169_), .Y(_5170_) );
OAI21X1 OAI21X1_1436 ( .gnd(gnd), .vdd(vdd), .A(_5136_), .B(micro_hash_ucr_2_pipe8), .C(_5131_), .Y(_5171_) );
AOI21X1 AOI21X1_913 ( .gnd(gnd), .vdd(vdd), .A(_5133_), .B(_5171_), .C(micro_hash_ucr_2_pipe11), .Y(_5172_) );
NAND3X1 NAND3X1_183 ( .gnd(gnd), .vdd(vdd), .A(_5119_), .B(_5124__bF_buf1), .C(_5130_), .Y(_5173_) );
NOR2X1 NOR2X1_935 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe15), .B(micro_hash_ucr_2_pipe17_bF_buf1), .Y(_5174_) );
NAND3X1 NAND3X1_184 ( .gnd(gnd), .vdd(vdd), .A(_5118__bF_buf2), .B(_5120__bF_buf1), .C(_5174_), .Y(_5175_) );
NOR2X1 NOR2X1_936 ( .gnd(gnd), .vdd(vdd), .A(_5173_), .B(_5175_), .Y(_5176_) );
NAND2X1 NAND2X1_605 ( .gnd(gnd), .vdd(vdd), .A(_5172_), .B(_5176_), .Y(_5177_) );
AOI21X1 AOI21X1_914 ( .gnd(gnd), .vdd(vdd), .A(_5139__bF_buf2), .B(_5177_), .C(_5170_), .Y(_5178_) );
NAND2X1 NAND2X1_606 ( .gnd(gnd), .vdd(vdd), .A(_5166_), .B(_5178_), .Y(_5179_) );
OAI21X1 OAI21X1_1437 ( .gnd(gnd), .vdd(vdd), .A(_5130_), .B(micro_hash_ucr_2_pipe14_bF_buf2), .C(_5125__bF_buf1), .Y(_5180_) );
AOI21X1 AOI21X1_915 ( .gnd(gnd), .vdd(vdd), .A(_5127__bF_buf1), .B(_5180_), .C(micro_hash_ucr_2_pipe17_bF_buf0), .Y(_5181_) );
OAI21X1 OAI21X1_1438 ( .gnd(gnd), .vdd(vdd), .A(_5181_), .B(micro_hash_ucr_2_pipe18_bF_buf2), .C(_5124__bF_buf0), .Y(_5182_) );
AOI21X1 AOI21X1_916 ( .gnd(gnd), .vdd(vdd), .A(_5123__bF_buf2), .B(_5182_), .C(micro_hash_ucr_2_pipe21_bF_buf1), .Y(_5183_) );
OAI21X1 OAI21X1_1439 ( .gnd(gnd), .vdd(vdd), .A(_5183_), .B(micro_hash_ucr_2_pipe22_bF_buf2), .C(_5120__bF_buf0), .Y(_5184_) );
AOI21X1 AOI21X1_917 ( .gnd(gnd), .vdd(vdd), .A(_5116__bF_buf3), .B(_5184_), .C(micro_hash_ucr_2_pipe25), .Y(_5185_) );
NAND2X1 NAND2X1_607 ( .gnd(gnd), .vdd(vdd), .A(_5117__bF_buf2), .B(_5148_), .Y(_5186_) );
OAI21X1 OAI21X1_1440 ( .gnd(gnd), .vdd(vdd), .A(_5185_), .B(_5186_), .C(_5179_), .Y(_5187_) );
AOI21X1 AOI21X1_918 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_0_), .B(_5157_), .C(_5187_), .Y(_5188_) );
OAI21X1 OAI21X1_1441 ( .gnd(gnd), .vdd(vdd), .A(_5188_), .B(micro_hash_ucr_2_pipe27), .C(_5150_), .Y(_5189_) );
OAI21X1 OAI21X1_1442 ( .gnd(gnd), .vdd(vdd), .A(_4630_), .B(_5115__bF_buf3), .C(_5114_), .Y(_5190_) );
AOI21X1 AOI21X1_919 ( .gnd(gnd), .vdd(vdd), .A(_5115__bF_buf2), .B(_5189_), .C(_5190_), .Y(_5191_) );
OAI21X1 OAI21X1_1443 ( .gnd(gnd), .vdd(vdd), .A(_5191_), .B(_5149_), .C(_5110__bF_buf2), .Y(_5192_) );
AOI21X1 AOI21X1_920 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe30_bF_buf3), .B(_4630_), .C(micro_hash_ucr_2_pipe31), .Y(_5193_) );
OAI21X1 OAI21X1_1444 ( .gnd(gnd), .vdd(vdd), .A(_5139__bF_buf1), .B(_5112__bF_buf2), .C(_5111__bF_buf3), .Y(_5194_) );
AOI21X1 AOI21X1_921 ( .gnd(gnd), .vdd(vdd), .A(_5193_), .B(_5192_), .C(_5194_), .Y(_5195_) );
NOR2X1 NOR2X1_937 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_0_), .B(_5111__bF_buf2), .Y(_5196_) );
OAI21X1 OAI21X1_1445 ( .gnd(gnd), .vdd(vdd), .A(_5195_), .B(_5196_), .C(_5107_), .Y(_5197_) );
OAI21X1 OAI21X1_1446 ( .gnd(gnd), .vdd(vdd), .A(_5107_), .B(_5148_), .C(_5197_), .Y(_5198_) );
NAND2X1 NAND2X1_608 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_0_), .B(micro_hash_ucr_2_pipe34_bF_buf2), .Y(_5199_) );
OAI21X1 OAI21X1_1447 ( .gnd(gnd), .vdd(vdd), .A(_5198_), .B(micro_hash_ucr_2_pipe34_bF_buf1), .C(_5199_), .Y(_5200_) );
NAND2X1 NAND2X1_609 ( .gnd(gnd), .vdd(vdd), .A(_5108__bF_buf2), .B(_5200_), .Y(_5201_) );
OAI21X1 OAI21X1_1448 ( .gnd(gnd), .vdd(vdd), .A(_5108__bF_buf1), .B(_5139__bF_buf0), .C(_5201_), .Y(_5202_) );
AOI21X1 AOI21X1_922 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe36_bF_buf2), .B(_4630_), .C(micro_hash_ucr_2_pipe37), .Y(_5203_) );
OAI21X1 OAI21X1_1449 ( .gnd(gnd), .vdd(vdd), .A(_5202_), .B(micro_hash_ucr_2_pipe36_bF_buf1), .C(_5203_), .Y(_5204_) );
AOI21X1 AOI21X1_923 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe37), .B(_5148_), .C(micro_hash_ucr_2_pipe38_bF_buf2), .Y(_5205_) );
AOI22X1 AOI22X1_40 ( .gnd(gnd), .vdd(vdd), .A(_4630_), .B(micro_hash_ucr_2_pipe38_bF_buf1), .C(_5204_), .D(_5205_), .Y(_5206_) );
NAND2X1 NAND2X1_610 ( .gnd(gnd), .vdd(vdd), .A(_5101_), .B(_5206_), .Y(_5207_) );
OAI21X1 OAI21X1_1450 ( .gnd(gnd), .vdd(vdd), .A(_5101_), .B(_5139__bF_buf3), .C(_5207_), .Y(_5208_) );
AOI21X1 AOI21X1_924 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe40_bF_buf3), .B(_4630_), .C(micro_hash_ucr_2_pipe41_bF_buf2), .Y(_5209_) );
OAI21X1 OAI21X1_1451 ( .gnd(gnd), .vdd(vdd), .A(_5208_), .B(micro_hash_ucr_2_pipe40_bF_buf2), .C(_5209_), .Y(_5210_) );
AOI21X1 AOI21X1_925 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe41_bF_buf1), .B(_5148_), .C(micro_hash_ucr_2_pipe42_bF_buf2), .Y(_5211_) );
AOI22X1 AOI22X1_41 ( .gnd(gnd), .vdd(vdd), .A(_4630_), .B(micro_hash_ucr_2_pipe42_bF_buf1), .C(_5210_), .D(_5211_), .Y(_5212_) );
NAND2X1 NAND2X1_611 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe43), .B(_5139__bF_buf2), .Y(_5213_) );
OAI21X1 OAI21X1_1452 ( .gnd(gnd), .vdd(vdd), .A(_5212_), .B(micro_hash_ucr_2_pipe43), .C(_5213_), .Y(_5214_) );
OAI21X1 OAI21X1_1453 ( .gnd(gnd), .vdd(vdd), .A(_5214_), .B(micro_hash_ucr_2_pipe44_bF_buf1), .C(_5147_), .Y(_5215_) );
NAND2X1 NAND2X1_612 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe45_bF_buf2), .B(_5139__bF_buf1), .Y(_5216_) );
OAI21X1 OAI21X1_1454 ( .gnd(gnd), .vdd(vdd), .A(_5215_), .B(micro_hash_ucr_2_pipe45_bF_buf1), .C(_5216_), .Y(_5217_) );
OAI21X1 OAI21X1_1455 ( .gnd(gnd), .vdd(vdd), .A(_5217_), .B(micro_hash_ucr_2_pipe46_bF_buf2), .C(_5146_), .Y(_5218_) );
NAND2X1 NAND2X1_613 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe47), .B(_5139__bF_buf0), .Y(_5219_) );
OAI21X1 OAI21X1_1456 ( .gnd(gnd), .vdd(vdd), .A(_5218_), .B(micro_hash_ucr_2_pipe47), .C(_5219_), .Y(_5220_) );
OAI21X1 OAI21X1_1457 ( .gnd(gnd), .vdd(vdd), .A(_5220_), .B(micro_hash_ucr_2_pipe48_bF_buf2), .C(_5145_), .Y(_5221_) );
NAND2X1 NAND2X1_614 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe49_bF_buf2), .B(_5139__bF_buf3), .Y(_5222_) );
OAI21X1 OAI21X1_1458 ( .gnd(gnd), .vdd(vdd), .A(_5221_), .B(micro_hash_ucr_2_pipe49_bF_buf1), .C(_5222_), .Y(_5223_) );
OAI21X1 OAI21X1_1459 ( .gnd(gnd), .vdd(vdd), .A(_5223_), .B(micro_hash_ucr_2_pipe50_bF_buf1), .C(_5144_), .Y(_5224_) );
NAND2X1 NAND2X1_615 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe51), .B(_5139__bF_buf2), .Y(_5225_) );
OAI21X1 OAI21X1_1460 ( .gnd(gnd), .vdd(vdd), .A(_5224_), .B(micro_hash_ucr_2_pipe51), .C(_5225_), .Y(_5226_) );
OAI21X1 OAI21X1_1461 ( .gnd(gnd), .vdd(vdd), .A(_5226_), .B(micro_hash_ucr_2_pipe52_bF_buf1), .C(_5143_), .Y(_5227_) );
NAND2X1 NAND2X1_616 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe53_bF_buf2), .B(_5139__bF_buf1), .Y(_5228_) );
OAI21X1 OAI21X1_1462 ( .gnd(gnd), .vdd(vdd), .A(_5227_), .B(micro_hash_ucr_2_pipe53_bF_buf1), .C(_5228_), .Y(_5229_) );
OAI21X1 OAI21X1_1463 ( .gnd(gnd), .vdd(vdd), .A(_5229_), .B(micro_hash_ucr_2_pipe54_bF_buf2), .C(_5142_), .Y(_5230_) );
NAND2X1 NAND2X1_617 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe55), .B(_5139__bF_buf0), .Y(_5231_) );
OAI21X1 OAI21X1_1464 ( .gnd(gnd), .vdd(vdd), .A(_5230_), .B(micro_hash_ucr_2_pipe55), .C(_5231_), .Y(_5232_) );
OAI21X1 OAI21X1_1465 ( .gnd(gnd), .vdd(vdd), .A(_5232_), .B(micro_hash_ucr_2_pipe56_bF_buf1), .C(_5141_), .Y(_5233_) );
NAND2X1 NAND2X1_618 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe57_bF_buf2), .B(_5139__bF_buf3), .Y(_5234_) );
OAI21X1 OAI21X1_1466 ( .gnd(gnd), .vdd(vdd), .A(_5233_), .B(micro_hash_ucr_2_pipe57_bF_buf1), .C(_5234_), .Y(_5235_) );
OAI21X1 OAI21X1_1467 ( .gnd(gnd), .vdd(vdd), .A(_5235_), .B(micro_hash_ucr_2_pipe58_bF_buf2), .C(_5140_), .Y(_5236_) );
NAND2X1 NAND2X1_619 ( .gnd(gnd), .vdd(vdd), .A(_5084__bF_buf2), .B(_5236_), .Y(_5237_) );
OAI21X1 OAI21X1_1468 ( .gnd(gnd), .vdd(vdd), .A(_5084__bF_buf1), .B(_5139__bF_buf2), .C(_5237_), .Y(_5238_) );
AOI21X1 AOI21X1_926 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe60_bF_buf3), .B(_4630_), .C(micro_hash_ucr_2_pipe61_bF_buf2), .Y(_5239_) );
OAI21X1 OAI21X1_1469 ( .gnd(gnd), .vdd(vdd), .A(_5238_), .B(micro_hash_ucr_2_pipe60_bF_buf2), .C(_5239_), .Y(_5240_) );
OAI21X1 OAI21X1_1470 ( .gnd(gnd), .vdd(vdd), .A(_5082_), .B(_5139__bF_buf1), .C(_5240_), .Y(_5241_) );
NAND2X1 NAND2X1_620 ( .gnd(gnd), .vdd(vdd), .A(_5081__bF_buf2), .B(_5241_), .Y(_5242_) );
OAI21X1 OAI21X1_1471 ( .gnd(gnd), .vdd(vdd), .A(_4630_), .B(_5081__bF_buf1), .C(_5242_), .Y(_5243_) );
NOR2X1 NOR2X1_938 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe63), .B(_5243_), .Y(_5244_) );
OAI21X1 OAI21X1_1472 ( .gnd(gnd), .vdd(vdd), .A(_5148_), .B(_5077__bF_buf2), .C(_5079__bF_buf3), .Y(_5245_) );
OAI22X1 OAI22X1_69 ( .gnd(gnd), .vdd(vdd), .A(_4630_), .B(_5079__bF_buf2), .C(_5244_), .D(_5245_), .Y(_5246_) );
NAND2X1 NAND2X1_621 ( .gnd(gnd), .vdd(vdd), .A(_5078_), .B(_5246_), .Y(_5247_) );
OAI21X1 OAI21X1_1473 ( .gnd(gnd), .vdd(vdd), .A(_5078_), .B(_5139__bF_buf0), .C(_5247_), .Y(_5248_) );
AOI21X1 AOI21X1_927 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe66_bF_buf3), .B(_4630_), .C(micro_hash_ucr_2_pipe67), .Y(_5249_) );
OAI21X1 OAI21X1_1474 ( .gnd(gnd), .vdd(vdd), .A(_5248_), .B(micro_hash_ucr_2_pipe66_bF_buf2), .C(_5249_), .Y(_5250_) );
OAI21X1 OAI21X1_1475 ( .gnd(gnd), .vdd(vdd), .A(_5076__bF_buf2), .B(_5139__bF_buf3), .C(_5250_), .Y(_5251_) );
MUX2X1 MUX2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_5251_), .B(micro_hash_ucr_2_a_0_), .S(_5075__bF_buf3), .Y(_5252_) );
OAI21X1 OAI21X1_1476 ( .gnd(gnd), .vdd(vdd), .A(_5148_), .B(_5073__bF_buf2), .C(_4496__bF_buf5), .Y(_5253_) );
AOI21X1 AOI21X1_928 ( .gnd(gnd), .vdd(vdd), .A(_5073__bF_buf1), .B(_5252_), .C(_5253_), .Y(_4491__0_) );
NOR2X1 NOR2X1_939 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_1_bF_buf1_), .B(micro_hash_ucr_2_b_1_bF_buf1_), .Y(_5254_) );
INVX8 INVX8_173 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_1_bF_buf0_), .Y(_5255_) );
NOR2X1 NOR2X1_940 ( .gnd(gnd), .vdd(vdd), .A(_5255_), .B(_8696_), .Y(_5256_) );
NOR2X1 NOR2X1_941 ( .gnd(gnd), .vdd(vdd), .A(_5254_), .B(_5256_), .Y(_5257_) );
NOR2X1 NOR2X1_942 ( .gnd(gnd), .vdd(vdd), .A(_4636_), .B(_5081__bF_buf0), .Y(_5258_) );
NAND2X1 NAND2X1_622 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_1_bF_buf1_), .B(micro_hash_ucr_2_pipe58_bF_buf1), .Y(_5259_) );
NAND2X1 NAND2X1_623 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_1_bF_buf0_), .B(micro_hash_ucr_2_pipe56_bF_buf0), .Y(_5260_) );
NAND2X1 NAND2X1_624 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_1_bF_buf3_), .B(micro_hash_ucr_2_pipe54_bF_buf1), .Y(_5261_) );
NAND2X1 NAND2X1_625 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_1_bF_buf2_), .B(micro_hash_ucr_2_pipe52_bF_buf0), .Y(_5262_) );
NOR2X1 NOR2X1_943 ( .gnd(gnd), .vdd(vdd), .A(_4636_), .B(_5097__bF_buf2), .Y(_5263_) );
NAND2X1 NAND2X1_626 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe38_bF_buf0), .B(_4636_), .Y(_5264_) );
INVX8 INVX8_174 ( .gnd(gnd), .vdd(vdd), .A(_5257_), .Y(_5265_) );
NAND2X1 NAND2X1_627 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_1_bF_buf1_), .B(micro_hash_ucr_2_pipe28_bF_buf2), .Y(_5266_) );
AOI21X1 AOI21X1_929 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe7), .B(_5135_), .C(micro_hash_ucr_2_pipe9), .Y(_5267_) );
OAI21X1 OAI21X1_1477 ( .gnd(gnd), .vdd(vdd), .A(_5267_), .B(micro_hash_ucr_2_pipe10), .C(_5132_), .Y(_5268_) );
AOI21X1 AOI21X1_930 ( .gnd(gnd), .vdd(vdd), .A(_5128_), .B(_5268_), .C(micro_hash_ucr_2_pipe13), .Y(_5269_) );
OAI21X1 OAI21X1_1478 ( .gnd(gnd), .vdd(vdd), .A(_5269_), .B(micro_hash_ucr_2_pipe14_bF_buf1), .C(_5125__bF_buf0), .Y(_5270_) );
NAND2X1 NAND2X1_628 ( .gnd(gnd), .vdd(vdd), .A(_5131_), .B(_5132_), .Y(_5271_) );
NOR2X1 NOR2X1_944 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe12_bF_buf2), .B(micro_hash_ucr_2_pipe14_bF_buf0), .Y(_5272_) );
NAND3X1 NAND3X1_185 ( .gnd(gnd), .vdd(vdd), .A(H_2_1_), .B(_5125__bF_buf3), .C(_5272_), .Y(_5273_) );
NOR2X1 NOR2X1_945 ( .gnd(gnd), .vdd(vdd), .A(_5271_), .B(_5273_), .Y(_5274_) );
NAND3X1 NAND3X1_186 ( .gnd(gnd), .vdd(vdd), .A(_5130_), .B(_5133_), .C(_5136_), .Y(_5275_) );
NOR2X1 NOR2X1_946 ( .gnd(gnd), .vdd(vdd), .A(_5158_), .B(_5275_), .Y(_5276_) );
AOI22X1 AOI22X1_42 ( .gnd(gnd), .vdd(vdd), .A(_5274_), .B(_5276_), .C(_5270_), .D(_5257_), .Y(_5277_) );
AOI21X1 AOI21X1_931 ( .gnd(gnd), .vdd(vdd), .A(_5130_), .B(_5160_), .C(micro_hash_ucr_2_pipe14_bF_buf4), .Y(_5278_) );
OAI21X1 OAI21X1_1479 ( .gnd(gnd), .vdd(vdd), .A(_5278_), .B(micro_hash_ucr_2_pipe15), .C(_5127__bF_buf0), .Y(_5279_) );
NAND2X1 NAND2X1_629 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_1_bF_buf0_), .B(_5279_), .Y(_5280_) );
OAI21X1 OAI21X1_1480 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe16_bF_buf2), .B(_5277_), .C(_5280_), .Y(_5281_) );
OAI21X1 OAI21X1_1481 ( .gnd(gnd), .vdd(vdd), .A(_5256_), .B(_5254_), .C(micro_hash_ucr_2_pipe17_bF_buf3), .Y(_5282_) );
OAI21X1 OAI21X1_1482 ( .gnd(gnd), .vdd(vdd), .A(_5281_), .B(micro_hash_ucr_2_pipe17_bF_buf2), .C(_5282_), .Y(_5283_) );
AOI21X1 AOI21X1_932 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_1_bF_buf3_), .B(micro_hash_ucr_2_pipe18_bF_buf1), .C(micro_hash_ucr_2_pipe19), .Y(_5284_) );
OAI21X1 OAI21X1_1483 ( .gnd(gnd), .vdd(vdd), .A(_5283_), .B(micro_hash_ucr_2_pipe18_bF_buf0), .C(_5284_), .Y(_5285_) );
OAI21X1 OAI21X1_1484 ( .gnd(gnd), .vdd(vdd), .A(_5124__bF_buf3), .B(_5257_), .C(_5285_), .Y(_5286_) );
NAND2X1 NAND2X1_630 ( .gnd(gnd), .vdd(vdd), .A(_5123__bF_buf1), .B(_5286_), .Y(_5287_) );
OAI21X1 OAI21X1_1485 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_1_bF_buf2_), .B(_5123__bF_buf0), .C(_5287_), .Y(_5288_) );
NAND2X1 NAND2X1_631 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe21_bF_buf0), .B(_5257_), .Y(_5289_) );
OAI21X1 OAI21X1_1486 ( .gnd(gnd), .vdd(vdd), .A(_5288_), .B(micro_hash_ucr_2_pipe21_bF_buf3), .C(_5289_), .Y(_5290_) );
NAND2X1 NAND2X1_632 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe22_bF_buf1), .B(_4636_), .Y(_5291_) );
OAI21X1 OAI21X1_1487 ( .gnd(gnd), .vdd(vdd), .A(_5290_), .B(micro_hash_ucr_2_pipe22_bF_buf0), .C(_5291_), .Y(_5292_) );
AOI21X1 AOI21X1_933 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe23), .B(_5257_), .C(micro_hash_ucr_2_pipe24_bF_buf0), .Y(_5293_) );
OAI21X1 OAI21X1_1488 ( .gnd(gnd), .vdd(vdd), .A(_5292_), .B(micro_hash_ucr_2_pipe23), .C(_5293_), .Y(_5294_) );
AOI21X1 AOI21X1_934 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe24_bF_buf3), .B(_4636_), .C(micro_hash_ucr_2_pipe25), .Y(_5295_) );
OAI21X1 OAI21X1_1489 ( .gnd(gnd), .vdd(vdd), .A(_5265_), .B(_5118__bF_buf1), .C(_5117__bF_buf1), .Y(_5296_) );
AOI21X1 AOI21X1_935 ( .gnd(gnd), .vdd(vdd), .A(_5295_), .B(_5294_), .C(_5296_), .Y(_5297_) );
NOR2X1 NOR2X1_947 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_1_bF_buf1_), .B(_5117__bF_buf0), .Y(_5298_) );
OAI21X1 OAI21X1_1490 ( .gnd(gnd), .vdd(vdd), .A(_5297_), .B(_5298_), .C(_5113_), .Y(_5299_) );
OAI21X1 OAI21X1_1491 ( .gnd(gnd), .vdd(vdd), .A(_5256_), .B(_5254_), .C(micro_hash_ucr_2_pipe27), .Y(_5300_) );
NAND3X1 NAND3X1_187 ( .gnd(gnd), .vdd(vdd), .A(_5115__bF_buf1), .B(_5300_), .C(_5299_), .Y(_5301_) );
AOI21X1 AOI21X1_936 ( .gnd(gnd), .vdd(vdd), .A(_5266_), .B(_5301_), .C(micro_hash_ucr_2_pipe29_bF_buf2), .Y(_5302_) );
OAI21X1 OAI21X1_1492 ( .gnd(gnd), .vdd(vdd), .A(_5265_), .B(_5114_), .C(_5110__bF_buf1), .Y(_5303_) );
AOI21X1 AOI21X1_937 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe30_bF_buf2), .B(_4636_), .C(micro_hash_ucr_2_pipe31), .Y(_5304_) );
OAI21X1 OAI21X1_1493 ( .gnd(gnd), .vdd(vdd), .A(_5302_), .B(_5303_), .C(_5304_), .Y(_5305_) );
OAI21X1 OAI21X1_1494 ( .gnd(gnd), .vdd(vdd), .A(_5112__bF_buf1), .B(_5265_), .C(_5305_), .Y(_5306_) );
NAND2X1 NAND2X1_633 ( .gnd(gnd), .vdd(vdd), .A(_5111__bF_buf1), .B(_5306_), .Y(_5307_) );
OAI21X1 OAI21X1_1495 ( .gnd(gnd), .vdd(vdd), .A(_4636_), .B(_5111__bF_buf0), .C(_5307_), .Y(_5308_) );
OAI21X1 OAI21X1_1496 ( .gnd(gnd), .vdd(vdd), .A(_5265_), .B(_5107_), .C(_5109__bF_buf3), .Y(_5309_) );
AOI21X1 AOI21X1_938 ( .gnd(gnd), .vdd(vdd), .A(_5107_), .B(_5308_), .C(_5309_), .Y(_5310_) );
OAI21X1 OAI21X1_1497 ( .gnd(gnd), .vdd(vdd), .A(_5109__bF_buf2), .B(micro_hash_ucr_2_a_1_bF_buf0_), .C(_5108__bF_buf0), .Y(_5311_) );
AOI21X1 AOI21X1_939 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe35), .B(_5257_), .C(micro_hash_ucr_2_pipe36_bF_buf0), .Y(_5312_) );
OAI21X1 OAI21X1_1498 ( .gnd(gnd), .vdd(vdd), .A(_5310_), .B(_5311_), .C(_5312_), .Y(_5313_) );
NAND2X1 NAND2X1_634 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe36_bF_buf3), .B(_4636_), .Y(_5314_) );
AOI21X1 AOI21X1_940 ( .gnd(gnd), .vdd(vdd), .A(_5314_), .B(_5313_), .C(micro_hash_ucr_2_pipe37), .Y(_5315_) );
NOR2X1 NOR2X1_948 ( .gnd(gnd), .vdd(vdd), .A(_5106_), .B(_5257_), .Y(_5316_) );
OAI21X1 OAI21X1_1499 ( .gnd(gnd), .vdd(vdd), .A(_5315_), .B(_5316_), .C(_5105__bF_buf3), .Y(_5317_) );
NAND3X1 NAND3X1_188 ( .gnd(gnd), .vdd(vdd), .A(_5101_), .B(_5264_), .C(_5317_), .Y(_5318_) );
AOI21X1 AOI21X1_941 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe39), .B(_5257_), .C(micro_hash_ucr_2_pipe40_bF_buf1), .Y(_5319_) );
OAI21X1 OAI21X1_1500 ( .gnd(gnd), .vdd(vdd), .A(_5103__bF_buf2), .B(micro_hash_ucr_2_a_1_bF_buf3_), .C(_5102_), .Y(_5320_) );
AOI21X1 AOI21X1_942 ( .gnd(gnd), .vdd(vdd), .A(_5319_), .B(_5318_), .C(_5320_), .Y(_5321_) );
OAI21X1 OAI21X1_1501 ( .gnd(gnd), .vdd(vdd), .A(_5265_), .B(_5102_), .C(_5098__bF_buf3), .Y(_5322_) );
OAI22X1 OAI22X1_70 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_1_bF_buf2_), .B(_5098__bF_buf2), .C(_5321_), .D(_5322_), .Y(_5323_) );
OAI21X1 OAI21X1_1502 ( .gnd(gnd), .vdd(vdd), .A(_5257_), .B(_5100__bF_buf2), .C(_5099__bF_buf3), .Y(_5324_) );
AOI21X1 AOI21X1_943 ( .gnd(gnd), .vdd(vdd), .A(_5100__bF_buf1), .B(_5323_), .C(_5324_), .Y(_5325_) );
NOR2X1 NOR2X1_949 ( .gnd(gnd), .vdd(vdd), .A(_4636_), .B(_5099__bF_buf2), .Y(_5326_) );
OAI21X1 OAI21X1_1503 ( .gnd(gnd), .vdd(vdd), .A(_5325_), .B(_5326_), .C(_5095_), .Y(_5327_) );
NAND2X1 NAND2X1_635 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe45_bF_buf0), .B(_5257_), .Y(_5328_) );
AOI21X1 AOI21X1_944 ( .gnd(gnd), .vdd(vdd), .A(_5328_), .B(_5327_), .C(micro_hash_ucr_2_pipe46_bF_buf1), .Y(_5329_) );
OAI21X1 OAI21X1_1504 ( .gnd(gnd), .vdd(vdd), .A(_5329_), .B(_5263_), .C(_5096__bF_buf2), .Y(_5330_) );
NAND2X1 NAND2X1_636 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe47), .B(_5257_), .Y(_5331_) );
AOI21X1 AOI21X1_945 ( .gnd(gnd), .vdd(vdd), .A(_5331_), .B(_5330_), .C(micro_hash_ucr_2_pipe48_bF_buf1), .Y(_5332_) );
OAI21X1 OAI21X1_1505 ( .gnd(gnd), .vdd(vdd), .A(_4636_), .B(_5092__bF_buf3), .C(_5094_), .Y(_5333_) );
AOI21X1 AOI21X1_946 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe49_bF_buf0), .B(_5265_), .C(micro_hash_ucr_2_pipe50_bF_buf0), .Y(_5334_) );
OAI21X1 OAI21X1_1506 ( .gnd(gnd), .vdd(vdd), .A(_5332_), .B(_5333_), .C(_5334_), .Y(_5335_) );
NAND2X1 NAND2X1_637 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_1_bF_buf1_), .B(micro_hash_ucr_2_pipe50_bF_buf3), .Y(_5336_) );
AOI21X1 AOI21X1_947 ( .gnd(gnd), .vdd(vdd), .A(_5336_), .B(_5335_), .C(micro_hash_ucr_2_pipe51), .Y(_5337_) );
NOR2X1 NOR2X1_950 ( .gnd(gnd), .vdd(vdd), .A(_5089__bF_buf2), .B(_5265_), .Y(_5338_) );
OAI21X1 OAI21X1_1507 ( .gnd(gnd), .vdd(vdd), .A(_5337_), .B(_5338_), .C(_5091__bF_buf3), .Y(_5339_) );
AOI21X1 AOI21X1_948 ( .gnd(gnd), .vdd(vdd), .A(_5262_), .B(_5339_), .C(micro_hash_ucr_2_pipe53_bF_buf0), .Y(_5340_) );
NOR2X1 NOR2X1_951 ( .gnd(gnd), .vdd(vdd), .A(_5090_), .B(_5265_), .Y(_5341_) );
OAI21X1 OAI21X1_1508 ( .gnd(gnd), .vdd(vdd), .A(_5340_), .B(_5341_), .C(_5086__bF_buf2), .Y(_5342_) );
AOI21X1 AOI21X1_949 ( .gnd(gnd), .vdd(vdd), .A(_5261_), .B(_5342_), .C(micro_hash_ucr_2_pipe55), .Y(_5343_) );
NOR2X1 NOR2X1_952 ( .gnd(gnd), .vdd(vdd), .A(_5088_), .B(_5265_), .Y(_5344_) );
OAI21X1 OAI21X1_1509 ( .gnd(gnd), .vdd(vdd), .A(_5343_), .B(_5344_), .C(_5087__bF_buf3), .Y(_5345_) );
AOI21X1 AOI21X1_950 ( .gnd(gnd), .vdd(vdd), .A(_5260_), .B(_5345_), .C(micro_hash_ucr_2_pipe57_bF_buf0), .Y(_5346_) );
NOR2X1 NOR2X1_953 ( .gnd(gnd), .vdd(vdd), .A(_5083_), .B(_5265_), .Y(_5347_) );
OAI21X1 OAI21X1_1510 ( .gnd(gnd), .vdd(vdd), .A(_5346_), .B(_5347_), .C(_5085__bF_buf2), .Y(_5348_) );
AOI21X1 AOI21X1_951 ( .gnd(gnd), .vdd(vdd), .A(_5259_), .B(_5348_), .C(micro_hash_ucr_2_pipe59), .Y(_5349_) );
OAI21X1 OAI21X1_1511 ( .gnd(gnd), .vdd(vdd), .A(_5265_), .B(_5084__bF_buf0), .C(_5080__bF_buf2), .Y(_5350_) );
AOI21X1 AOI21X1_952 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe60_bF_buf1), .B(_4636_), .C(micro_hash_ucr_2_pipe61_bF_buf1), .Y(_5351_) );
OAI21X1 OAI21X1_1512 ( .gnd(gnd), .vdd(vdd), .A(_5349_), .B(_5350_), .C(_5351_), .Y(_5352_) );
NAND2X1 NAND2X1_638 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe61_bF_buf0), .B(_5257_), .Y(_5353_) );
AOI21X1 AOI21X1_953 ( .gnd(gnd), .vdd(vdd), .A(_5353_), .B(_5352_), .C(micro_hash_ucr_2_pipe62_bF_buf3), .Y(_5354_) );
OAI21X1 OAI21X1_1513 ( .gnd(gnd), .vdd(vdd), .A(_5354_), .B(_5258_), .C(_5077__bF_buf1), .Y(_5355_) );
NAND2X1 NAND2X1_639 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe63), .B(_5257_), .Y(_5356_) );
AOI21X1 AOI21X1_954 ( .gnd(gnd), .vdd(vdd), .A(_5356_), .B(_5355_), .C(micro_hash_ucr_2_pipe64_bF_buf3), .Y(_5357_) );
OAI21X1 OAI21X1_1514 ( .gnd(gnd), .vdd(vdd), .A(_4636_), .B(_5079__bF_buf1), .C(_5078_), .Y(_5358_) );
OAI22X1 OAI22X1_71 ( .gnd(gnd), .vdd(vdd), .A(_5078_), .B(_5257_), .C(_5357_), .D(_5358_), .Y(_5359_) );
OAI21X1 OAI21X1_1515 ( .gnd(gnd), .vdd(vdd), .A(_5074__bF_buf2), .B(micro_hash_ucr_2_a_1_bF_buf0_), .C(_5076__bF_buf1), .Y(_5360_) );
AOI21X1 AOI21X1_955 ( .gnd(gnd), .vdd(vdd), .A(_5074__bF_buf1), .B(_5359_), .C(_5360_), .Y(_5361_) );
OAI21X1 OAI21X1_1516 ( .gnd(gnd), .vdd(vdd), .A(_5265_), .B(_5076__bF_buf0), .C(_5075__bF_buf2), .Y(_5362_) );
OAI22X1 OAI22X1_72 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_1_bF_buf3_), .B(_5075__bF_buf1), .C(_5361_), .D(_5362_), .Y(_5363_) );
OAI21X1 OAI21X1_1517 ( .gnd(gnd), .vdd(vdd), .A(_5257_), .B(_5073__bF_buf0), .C(_4496__bF_buf4), .Y(_5364_) );
AOI21X1 AOI21X1_956 ( .gnd(gnd), .vdd(vdd), .A(_5073__bF_buf3), .B(_5363_), .C(_5364_), .Y(_4491__1_) );
INVX8 INVX8_175 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_2_), .Y(_5365_) );
NAND2X1 NAND2X1_640 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_2_), .B(micro_hash_ucr_2_pipe62_bF_buf2), .Y(_5366_) );
NAND2X1 NAND2X1_641 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_2_), .B(micro_hash_ucr_2_pipe60_bF_buf0), .Y(_5367_) );
NAND2X1 NAND2X1_642 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe54_bF_buf0), .B(_5365__bF_buf3), .Y(_5368_) );
NAND2X1 NAND2X1_643 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe52_bF_buf3), .B(_5365__bF_buf2), .Y(_5369_) );
NAND2X1 NAND2X1_644 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe50_bF_buf2), .B(_5365__bF_buf1), .Y(_5370_) );
NAND2X1 NAND2X1_645 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe48_bF_buf0), .B(_5365__bF_buf0), .Y(_5371_) );
INVX8 INVX8_176 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_2_bF_buf1_), .Y(_5372_) );
NAND2X1 NAND2X1_646 ( .gnd(gnd), .vdd(vdd), .A(_5372_), .B(_4583_), .Y(_5373_) );
NAND2X1 NAND2X1_647 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_2_bF_buf0_), .B(micro_hash_ucr_2_b_2_bF_buf1_), .Y(_5374_) );
NAND2X1 NAND2X1_648 ( .gnd(gnd), .vdd(vdd), .A(_5374_), .B(_5373_), .Y(_5375_) );
NOR2X1 NOR2X1_954 ( .gnd(gnd), .vdd(vdd), .A(_5365__bF_buf3), .B(_5115__bF_buf0), .Y(_5376_) );
NOR2X1 NOR2X1_955 ( .gnd(gnd), .vdd(vdd), .A(_5365__bF_buf2), .B(_5117__bF_buf4), .Y(_5377_) );
NOR2X1 NOR2X1_956 ( .gnd(gnd), .vdd(vdd), .A(_5365__bF_buf1), .B(_5116__bF_buf2), .Y(_5378_) );
NOR2X1 NOR2X1_957 ( .gnd(gnd), .vdd(vdd), .A(_5365__bF_buf0), .B(_5121__bF_buf2), .Y(_5379_) );
INVX8 INVX8_177 ( .gnd(gnd), .vdd(vdd), .A(_5375_), .Y(_5380_) );
NAND2X1 NAND2X1_649 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe17_bF_buf1), .B(_5380__bF_buf3), .Y(_5381_) );
NAND2X1 NAND2X1_650 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe15), .B(_5380__bF_buf2), .Y(_5382_) );
AOI21X1 AOI21X1_957 ( .gnd(gnd), .vdd(vdd), .A(_5134_), .B(_5136_), .C(micro_hash_ucr_2_pipe8), .Y(_5383_) );
OAI21X1 OAI21X1_1518 ( .gnd(gnd), .vdd(vdd), .A(_5383_), .B(micro_hash_ucr_2_pipe9), .C(_5133_), .Y(_5384_) );
AOI21X1 AOI21X1_958 ( .gnd(gnd), .vdd(vdd), .A(_5132_), .B(_5384_), .C(micro_hash_ucr_2_pipe12_bF_buf1), .Y(_5385_) );
OR2X2 OR2X2_46 ( .gnd(gnd), .vdd(vdd), .A(_5158_), .B(_5271_), .Y(_5386_) );
NOR2X1 NOR2X1_958 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe12_bF_buf0), .B(micro_hash_ucr_2_pipe10), .Y(_5387_) );
NOR2X1 NOR2X1_959 ( .gnd(gnd), .vdd(vdd), .A(H_2_2_), .B(micro_hash_ucr_2_pipe7), .Y(_5388_) );
NAND2X1 NAND2X1_651 ( .gnd(gnd), .vdd(vdd), .A(_5387_), .B(_5388_), .Y(_5389_) );
OAI22X1 OAI22X1_73 ( .gnd(gnd), .vdd(vdd), .A(_5386_), .B(_5389_), .C(_5385_), .D(micro_hash_ucr_2_a_2_), .Y(_5390_) );
NAND2X1 NAND2X1_652 ( .gnd(gnd), .vdd(vdd), .A(_5130_), .B(_5390_), .Y(_5391_) );
OAI21X1 OAI21X1_1519 ( .gnd(gnd), .vdd(vdd), .A(_5172_), .B(micro_hash_ucr_2_pipe12_bF_buf3), .C(_5130_), .Y(_5392_) );
AOI21X1 AOI21X1_959 ( .gnd(gnd), .vdd(vdd), .A(_5375_), .B(_5392_), .C(micro_hash_ucr_2_pipe14_bF_buf3), .Y(_5393_) );
AOI22X1 AOI22X1_43 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_2_), .B(micro_hash_ucr_2_pipe14_bF_buf2), .C(_5391_), .D(_5393_), .Y(_5394_) );
OAI21X1 OAI21X1_1520 ( .gnd(gnd), .vdd(vdd), .A(_5394_), .B(micro_hash_ucr_2_pipe15), .C(_5382_), .Y(_5395_) );
NAND2X1 NAND2X1_653 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe16_bF_buf1), .B(_5365__bF_buf3), .Y(_5396_) );
OAI21X1 OAI21X1_1521 ( .gnd(gnd), .vdd(vdd), .A(_5395_), .B(micro_hash_ucr_2_pipe16_bF_buf0), .C(_5396_), .Y(_5397_) );
OAI21X1 OAI21X1_1522 ( .gnd(gnd), .vdd(vdd), .A(_5397_), .B(micro_hash_ucr_2_pipe17_bF_buf0), .C(_5381_), .Y(_5398_) );
NAND2X1 NAND2X1_654 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe18_bF_buf4), .B(_5365__bF_buf2), .Y(_5399_) );
OAI21X1 OAI21X1_1523 ( .gnd(gnd), .vdd(vdd), .A(_5398_), .B(micro_hash_ucr_2_pipe18_bF_buf3), .C(_5399_), .Y(_5400_) );
OAI21X1 OAI21X1_1524 ( .gnd(gnd), .vdd(vdd), .A(_5380__bF_buf1), .B(_5124__bF_buf2), .C(_5123__bF_buf4), .Y(_5401_) );
AOI21X1 AOI21X1_960 ( .gnd(gnd), .vdd(vdd), .A(_5124__bF_buf1), .B(_5400_), .C(_5401_), .Y(_5402_) );
NOR2X1 NOR2X1_960 ( .gnd(gnd), .vdd(vdd), .A(_5365__bF_buf1), .B(_5123__bF_buf3), .Y(_5403_) );
OAI21X1 OAI21X1_1525 ( .gnd(gnd), .vdd(vdd), .A(_5402_), .B(_5403_), .C(_5119_), .Y(_5404_) );
NAND2X1 NAND2X1_655 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe21_bF_buf2), .B(_5380__bF_buf0), .Y(_5405_) );
AOI21X1 AOI21X1_961 ( .gnd(gnd), .vdd(vdd), .A(_5405_), .B(_5404_), .C(micro_hash_ucr_2_pipe22_bF_buf4), .Y(_5406_) );
OAI21X1 OAI21X1_1526 ( .gnd(gnd), .vdd(vdd), .A(_5406_), .B(_5379_), .C(_5120__bF_buf3), .Y(_5407_) );
NAND2X1 NAND2X1_656 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe23), .B(_5380__bF_buf3), .Y(_5408_) );
AOI21X1 AOI21X1_962 ( .gnd(gnd), .vdd(vdd), .A(_5408_), .B(_5407_), .C(micro_hash_ucr_2_pipe24_bF_buf2), .Y(_5409_) );
OAI21X1 OAI21X1_1527 ( .gnd(gnd), .vdd(vdd), .A(_5409_), .B(_5378_), .C(_5118__bF_buf0), .Y(_5410_) );
NAND2X1 NAND2X1_657 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe25), .B(_5380__bF_buf2), .Y(_5411_) );
AOI21X1 AOI21X1_963 ( .gnd(gnd), .vdd(vdd), .A(_5411_), .B(_5410_), .C(micro_hash_ucr_2_pipe26_bF_buf1), .Y(_5412_) );
OAI21X1 OAI21X1_1528 ( .gnd(gnd), .vdd(vdd), .A(_5412_), .B(_5377_), .C(_5113_), .Y(_5413_) );
NAND2X1 NAND2X1_658 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe27), .B(_5380__bF_buf1), .Y(_5414_) );
AOI21X1 AOI21X1_964 ( .gnd(gnd), .vdd(vdd), .A(_5414_), .B(_5413_), .C(micro_hash_ucr_2_pipe28_bF_buf1), .Y(_5415_) );
OAI21X1 OAI21X1_1529 ( .gnd(gnd), .vdd(vdd), .A(_5415_), .B(_5376_), .C(_5114_), .Y(_5416_) );
AOI21X1 AOI21X1_965 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe29_bF_buf1), .B(_5380__bF_buf0), .C(micro_hash_ucr_2_pipe30_bF_buf1), .Y(_5417_) );
OAI21X1 OAI21X1_1530 ( .gnd(gnd), .vdd(vdd), .A(_5110__bF_buf0), .B(micro_hash_ucr_2_a_2_), .C(_5112__bF_buf0), .Y(_5418_) );
AOI21X1 AOI21X1_966 ( .gnd(gnd), .vdd(vdd), .A(_5417_), .B(_5416_), .C(_5418_), .Y(_5419_) );
OAI21X1 OAI21X1_1531 ( .gnd(gnd), .vdd(vdd), .A(_5375_), .B(_5112__bF_buf3), .C(_5111__bF_buf4), .Y(_5420_) );
OAI22X1 OAI22X1_74 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_2_), .B(_5111__bF_buf3), .C(_5419_), .D(_5420_), .Y(_5421_) );
AOI21X1 AOI21X1_967 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe33_bF_buf2), .B(_5380__bF_buf3), .C(micro_hash_ucr_2_pipe34_bF_buf0), .Y(_5422_) );
OAI21X1 OAI21X1_1532 ( .gnd(gnd), .vdd(vdd), .A(_5421_), .B(micro_hash_ucr_2_pipe33_bF_buf1), .C(_5422_), .Y(_5423_) );
AOI21X1 AOI21X1_968 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe34_bF_buf3), .B(_5365__bF_buf0), .C(micro_hash_ucr_2_pipe35), .Y(_5424_) );
OAI21X1 OAI21X1_1533 ( .gnd(gnd), .vdd(vdd), .A(_5375_), .B(_5108__bF_buf3), .C(_5104__bF_buf3), .Y(_5425_) );
AOI21X1 AOI21X1_969 ( .gnd(gnd), .vdd(vdd), .A(_5424_), .B(_5423_), .C(_5425_), .Y(_5426_) );
NOR2X1 NOR2X1_961 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_2_), .B(_5104__bF_buf2), .Y(_5427_) );
OAI21X1 OAI21X1_1534 ( .gnd(gnd), .vdd(vdd), .A(_5426_), .B(_5427_), .C(_5106_), .Y(_5428_) );
NAND2X1 NAND2X1_659 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe37), .B(_5375_), .Y(_5429_) );
NAND3X1 NAND3X1_189 ( .gnd(gnd), .vdd(vdd), .A(_5105__bF_buf2), .B(_5429_), .C(_5428_), .Y(_5430_) );
AOI21X1 AOI21X1_970 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_2_), .B(micro_hash_ucr_2_pipe38_bF_buf3), .C(micro_hash_ucr_2_pipe39), .Y(_5431_) );
AOI22X1 AOI22X1_44 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe39), .B(_5375_), .C(_5430_), .D(_5431_), .Y(_5432_) );
AOI21X1 AOI21X1_971 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe40_bF_buf0), .B(_5365__bF_buf3), .C(micro_hash_ucr_2_pipe41_bF_buf0), .Y(_5433_) );
OAI21X1 OAI21X1_1535 ( .gnd(gnd), .vdd(vdd), .A(_5432_), .B(micro_hash_ucr_2_pipe40_bF_buf4), .C(_5433_), .Y(_5434_) );
AOI21X1 AOI21X1_972 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe41_bF_buf3), .B(_5380__bF_buf2), .C(micro_hash_ucr_2_pipe42_bF_buf0), .Y(_5435_) );
AOI22X1 AOI22X1_45 ( .gnd(gnd), .vdd(vdd), .A(_5365__bF_buf2), .B(micro_hash_ucr_2_pipe42_bF_buf3), .C(_5434_), .D(_5435_), .Y(_5436_) );
OAI21X1 OAI21X1_1536 ( .gnd(gnd), .vdd(vdd), .A(_5375_), .B(_5100__bF_buf0), .C(_5099__bF_buf1), .Y(_5437_) );
AOI21X1 AOI21X1_973 ( .gnd(gnd), .vdd(vdd), .A(_5100__bF_buf3), .B(_5436_), .C(_5437_), .Y(_5438_) );
OAI21X1 OAI21X1_1537 ( .gnd(gnd), .vdd(vdd), .A(_5099__bF_buf0), .B(micro_hash_ucr_2_a_2_), .C(_5095_), .Y(_5439_) );
AOI21X1 AOI21X1_974 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe45_bF_buf3), .B(_5380__bF_buf1), .C(micro_hash_ucr_2_pipe46_bF_buf0), .Y(_5440_) );
OAI21X1 OAI21X1_1538 ( .gnd(gnd), .vdd(vdd), .A(_5438_), .B(_5439_), .C(_5440_), .Y(_5441_) );
NAND2X1 NAND2X1_660 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe46_bF_buf4), .B(_5365__bF_buf1), .Y(_5442_) );
AOI21X1 AOI21X1_975 ( .gnd(gnd), .vdd(vdd), .A(_5442_), .B(_5441_), .C(micro_hash_ucr_2_pipe47), .Y(_5443_) );
NOR2X1 NOR2X1_962 ( .gnd(gnd), .vdd(vdd), .A(_5096__bF_buf1), .B(_5380__bF_buf0), .Y(_5444_) );
OAI21X1 OAI21X1_1539 ( .gnd(gnd), .vdd(vdd), .A(_5443_), .B(_5444_), .C(_5092__bF_buf2), .Y(_5445_) );
AOI21X1 AOI21X1_976 ( .gnd(gnd), .vdd(vdd), .A(_5371_), .B(_5445_), .C(micro_hash_ucr_2_pipe49_bF_buf3), .Y(_5446_) );
NOR2X1 NOR2X1_963 ( .gnd(gnd), .vdd(vdd), .A(_5094_), .B(_5380__bF_buf3), .Y(_5447_) );
OAI21X1 OAI21X1_1540 ( .gnd(gnd), .vdd(vdd), .A(_5446_), .B(_5447_), .C(_5093__bF_buf3), .Y(_5448_) );
AOI21X1 AOI21X1_977 ( .gnd(gnd), .vdd(vdd), .A(_5370_), .B(_5448_), .C(micro_hash_ucr_2_pipe51), .Y(_5449_) );
NOR2X1 NOR2X1_964 ( .gnd(gnd), .vdd(vdd), .A(_5089__bF_buf1), .B(_5380__bF_buf2), .Y(_5450_) );
OAI21X1 OAI21X1_1541 ( .gnd(gnd), .vdd(vdd), .A(_5449_), .B(_5450_), .C(_5091__bF_buf2), .Y(_5451_) );
AOI21X1 AOI21X1_978 ( .gnd(gnd), .vdd(vdd), .A(_5369_), .B(_5451_), .C(micro_hash_ucr_2_pipe53_bF_buf3), .Y(_5452_) );
NOR2X1 NOR2X1_965 ( .gnd(gnd), .vdd(vdd), .A(_5090_), .B(_5380__bF_buf1), .Y(_5453_) );
OAI21X1 OAI21X1_1542 ( .gnd(gnd), .vdd(vdd), .A(_5452_), .B(_5453_), .C(_5086__bF_buf1), .Y(_5454_) );
NAND3X1 NAND3X1_190 ( .gnd(gnd), .vdd(vdd), .A(_5088_), .B(_5368_), .C(_5454_), .Y(_5455_) );
NAND2X1 NAND2X1_661 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe55), .B(_5380__bF_buf0), .Y(_5456_) );
AOI21X1 AOI21X1_979 ( .gnd(gnd), .vdd(vdd), .A(_5456_), .B(_5455_), .C(micro_hash_ucr_2_pipe56_bF_buf3), .Y(_5457_) );
OAI21X1 OAI21X1_1543 ( .gnd(gnd), .vdd(vdd), .A(_5365__bF_buf0), .B(_5087__bF_buf2), .C(_5083_), .Y(_5458_) );
AOI21X1 AOI21X1_980 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe57_bF_buf3), .B(_5375_), .C(micro_hash_ucr_2_pipe58_bF_buf0), .Y(_5459_) );
OAI21X1 OAI21X1_1544 ( .gnd(gnd), .vdd(vdd), .A(_5457_), .B(_5458_), .C(_5459_), .Y(_5460_) );
NAND2X1 NAND2X1_662 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_2_), .B(micro_hash_ucr_2_pipe58_bF_buf4), .Y(_5461_) );
AOI21X1 AOI21X1_981 ( .gnd(gnd), .vdd(vdd), .A(_5461_), .B(_5460_), .C(micro_hash_ucr_2_pipe59), .Y(_5462_) );
NOR2X1 NOR2X1_966 ( .gnd(gnd), .vdd(vdd), .A(_5084__bF_buf3), .B(_5375_), .Y(_5463_) );
OAI21X1 OAI21X1_1545 ( .gnd(gnd), .vdd(vdd), .A(_5462_), .B(_5463_), .C(_5080__bF_buf1), .Y(_5464_) );
AOI21X1 AOI21X1_982 ( .gnd(gnd), .vdd(vdd), .A(_5367_), .B(_5464_), .C(micro_hash_ucr_2_pipe61_bF_buf3), .Y(_5465_) );
NOR2X1 NOR2X1_967 ( .gnd(gnd), .vdd(vdd), .A(_5082_), .B(_5375_), .Y(_5466_) );
OAI21X1 OAI21X1_1546 ( .gnd(gnd), .vdd(vdd), .A(_5465_), .B(_5466_), .C(_5081__bF_buf3), .Y(_5467_) );
AOI21X1 AOI21X1_983 ( .gnd(gnd), .vdd(vdd), .A(_5366_), .B(_5467_), .C(micro_hash_ucr_2_pipe63), .Y(_5468_) );
OAI21X1 OAI21X1_1547 ( .gnd(gnd), .vdd(vdd), .A(_5375_), .B(_5077__bF_buf0), .C(_5079__bF_buf0), .Y(_5469_) );
AOI21X1 AOI21X1_984 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe64_bF_buf2), .B(_5365__bF_buf3), .C(micro_hash_ucr_2_pipe65_bF_buf2), .Y(_5470_) );
OAI21X1 OAI21X1_1548 ( .gnd(gnd), .vdd(vdd), .A(_5468_), .B(_5469_), .C(_5470_), .Y(_5471_) );
AOI21X1 AOI21X1_985 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe65_bF_buf1), .B(_5380__bF_buf3), .C(micro_hash_ucr_2_pipe66_bF_buf1), .Y(_5472_) );
AOI22X1 AOI22X1_46 ( .gnd(gnd), .vdd(vdd), .A(_5365__bF_buf2), .B(micro_hash_ucr_2_pipe66_bF_buf0), .C(_5471_), .D(_5472_), .Y(_5473_) );
AOI21X1 AOI21X1_986 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe67), .B(_5375_), .C(micro_hash_ucr_2_pipe68), .Y(_5474_) );
OAI21X1 OAI21X1_1549 ( .gnd(gnd), .vdd(vdd), .A(_5473_), .B(micro_hash_ucr_2_pipe67), .C(_5474_), .Y(_5475_) );
AOI21X1 AOI21X1_987 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_2_), .B(micro_hash_ucr_2_pipe68), .C(micro_hash_ucr_2_pipe69), .Y(_5476_) );
OAI21X1 OAI21X1_1550 ( .gnd(gnd), .vdd(vdd), .A(_5380__bF_buf2), .B(_5073__bF_buf2), .C(_4496__bF_buf3), .Y(_5477_) );
AOI21X1 AOI21X1_988 ( .gnd(gnd), .vdd(vdd), .A(_5476_), .B(_5475_), .C(_5477_), .Y(_4491__2_) );
NAND2X1 NAND2X1_663 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe64_bF_buf1), .B(_4654__bF_buf2), .Y(_5478_) );
NAND2X1 NAND2X1_664 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe54_bF_buf4), .B(_4654__bF_buf1), .Y(_5479_) );
NAND2X1 NAND2X1_665 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe52_bF_buf2), .B(_4654__bF_buf0), .Y(_5480_) );
NAND2X1 NAND2X1_666 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe50_bF_buf1), .B(_4654__bF_buf3), .Y(_5481_) );
NAND2X1 NAND2X1_667 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe48_bF_buf4), .B(_4654__bF_buf2), .Y(_5482_) );
NAND2X1 NAND2X1_668 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe46_bF_buf3), .B(_4654__bF_buf1), .Y(_5483_) );
NAND2X1 NAND2X1_669 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe44_bF_buf0), .B(_4654__bF_buf0), .Y(_5484_) );
NAND2X1 NAND2X1_670 ( .gnd(gnd), .vdd(vdd), .A(_8654_), .B(_4588_), .Y(_5485_) );
NAND2X1 NAND2X1_671 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_3_bF_buf1_), .B(micro_hash_ucr_2_b_3_bF_buf1_), .Y(_5486_) );
AND2X2 AND2X2_426 ( .gnd(gnd), .vdd(vdd), .A(_5485_), .B(_5486_), .Y(_5487_) );
NAND2X1 NAND2X1_672 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe26_bF_buf0), .B(_4654__bF_buf3), .Y(_5488_) );
NAND2X1 NAND2X1_673 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe17_bF_buf3), .B(_5487__bF_buf3), .Y(_5489_) );
NOR2X1 NOR2X1_968 ( .gnd(gnd), .vdd(vdd), .A(_4654__bF_buf2), .B(_5127__bF_buf3), .Y(_5490_) );
NAND2X1 NAND2X1_674 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe15), .B(_5487__bF_buf2), .Y(_5491_) );
NAND3X1 NAND3X1_191 ( .gnd(gnd), .vdd(vdd), .A(_4653_), .B(_5131_), .C(_5136_), .Y(_5492_) );
NOR2X1 NOR2X1_969 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe8), .B(_5134_), .Y(_5493_) );
NOR2X1 NOR2X1_970 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe13), .B(micro_hash_ucr_2_pipe11), .Y(_5494_) );
NAND3X1 NAND3X1_192 ( .gnd(gnd), .vdd(vdd), .A(_5387_), .B(_5494_), .C(_5493_), .Y(_5495_) );
OAI22X1 OAI22X1_75 ( .gnd(gnd), .vdd(vdd), .A(_5492_), .B(_5495_), .C(_5269_), .D(_5487__bF_buf1), .Y(_5496_) );
AOI21X1 AOI21X1_989 ( .gnd(gnd), .vdd(vdd), .A(_5129_), .B(_5496_), .C(micro_hash_ucr_2_pipe15), .Y(_5497_) );
OAI21X1 OAI21X1_1551 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_3_), .B(_5278_), .C(_5497_), .Y(_5498_) );
AOI21X1 AOI21X1_990 ( .gnd(gnd), .vdd(vdd), .A(_5491_), .B(_5498_), .C(micro_hash_ucr_2_pipe16_bF_buf4), .Y(_5499_) );
OAI21X1 OAI21X1_1552 ( .gnd(gnd), .vdd(vdd), .A(_5499_), .B(_5490_), .C(_5126_), .Y(_5500_) );
AOI21X1 AOI21X1_991 ( .gnd(gnd), .vdd(vdd), .A(_5489_), .B(_5500_), .C(micro_hash_ucr_2_pipe18_bF_buf2), .Y(_5501_) );
OAI21X1 OAI21X1_1553 ( .gnd(gnd), .vdd(vdd), .A(_4654__bF_buf1), .B(_5122__bF_buf2), .C(_5124__bF_buf0), .Y(_5502_) );
INVX4 INVX4_103 ( .gnd(gnd), .vdd(vdd), .A(_5487__bF_buf0), .Y(_5503_) );
AOI21X1 AOI21X1_992 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe19), .B(_5503_), .C(micro_hash_ucr_2_pipe20_bF_buf1), .Y(_5504_) );
OAI21X1 OAI21X1_1554 ( .gnd(gnd), .vdd(vdd), .A(_5501_), .B(_5502_), .C(_5504_), .Y(_5505_) );
NAND2X1 NAND2X1_675 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_3_), .B(micro_hash_ucr_2_pipe20_bF_buf0), .Y(_5506_) );
AOI21X1 AOI21X1_993 ( .gnd(gnd), .vdd(vdd), .A(_5506_), .B(_5505_), .C(micro_hash_ucr_2_pipe21_bF_buf1), .Y(_5507_) );
NOR2X1 NOR2X1_971 ( .gnd(gnd), .vdd(vdd), .A(_5119_), .B(_5503_), .Y(_5508_) );
OAI21X1 OAI21X1_1555 ( .gnd(gnd), .vdd(vdd), .A(_5507_), .B(_5508_), .C(_5121__bF_buf1), .Y(_5509_) );
AOI21X1 AOI21X1_994 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_3_), .B(micro_hash_ucr_2_pipe22_bF_buf3), .C(micro_hash_ucr_2_pipe23), .Y(_5510_) );
OAI21X1 OAI21X1_1556 ( .gnd(gnd), .vdd(vdd), .A(_5487__bF_buf3), .B(_5120__bF_buf2), .C(_5116__bF_buf1), .Y(_5511_) );
AOI21X1 AOI21X1_995 ( .gnd(gnd), .vdd(vdd), .A(_5510_), .B(_5509_), .C(_5511_), .Y(_5512_) );
NOR2X1 NOR2X1_972 ( .gnd(gnd), .vdd(vdd), .A(_4654__bF_buf0), .B(_5116__bF_buf0), .Y(_5513_) );
OAI21X1 OAI21X1_1557 ( .gnd(gnd), .vdd(vdd), .A(_5512_), .B(_5513_), .C(_5118__bF_buf3), .Y(_5514_) );
NAND2X1 NAND2X1_676 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe25), .B(_5487__bF_buf2), .Y(_5515_) );
NAND3X1 NAND3X1_193 ( .gnd(gnd), .vdd(vdd), .A(_5117__bF_buf3), .B(_5515_), .C(_5514_), .Y(_5516_) );
NAND3X1 NAND3X1_194 ( .gnd(gnd), .vdd(vdd), .A(_5113_), .B(_5488_), .C(_5516_), .Y(_5517_) );
NAND2X1 NAND2X1_677 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe27), .B(_5487__bF_buf1), .Y(_5518_) );
AOI21X1 AOI21X1_996 ( .gnd(gnd), .vdd(vdd), .A(_5518_), .B(_5517_), .C(micro_hash_ucr_2_pipe28_bF_buf0), .Y(_5519_) );
OAI21X1 OAI21X1_1558 ( .gnd(gnd), .vdd(vdd), .A(_4654__bF_buf3), .B(_5115__bF_buf4), .C(_5114_), .Y(_5520_) );
OAI22X1 OAI22X1_76 ( .gnd(gnd), .vdd(vdd), .A(_5114_), .B(_5487__bF_buf0), .C(_5519_), .D(_5520_), .Y(_5521_) );
OAI21X1 OAI21X1_1559 ( .gnd(gnd), .vdd(vdd), .A(_5110__bF_buf3), .B(micro_hash_ucr_2_a_3_), .C(_5112__bF_buf2), .Y(_5522_) );
AOI21X1 AOI21X1_997 ( .gnd(gnd), .vdd(vdd), .A(_5110__bF_buf2), .B(_5521_), .C(_5522_), .Y(_5523_) );
OAI21X1 OAI21X1_1560 ( .gnd(gnd), .vdd(vdd), .A(_5503_), .B(_5112__bF_buf1), .C(_5111__bF_buf2), .Y(_5524_) );
OAI22X1 OAI22X1_77 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_3_), .B(_5111__bF_buf1), .C(_5523_), .D(_5524_), .Y(_5525_) );
NAND2X1 NAND2X1_678 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe33_bF_buf0), .B(_5487__bF_buf3), .Y(_5526_) );
OAI21X1 OAI21X1_1561 ( .gnd(gnd), .vdd(vdd), .A(_5525_), .B(micro_hash_ucr_2_pipe33_bF_buf3), .C(_5526_), .Y(_5527_) );
NAND2X1 NAND2X1_679 ( .gnd(gnd), .vdd(vdd), .A(_5109__bF_buf1), .B(_5527_), .Y(_5528_) );
OAI21X1 OAI21X1_1562 ( .gnd(gnd), .vdd(vdd), .A(_4654__bF_buf2), .B(_5109__bF_buf0), .C(_5528_), .Y(_5529_) );
NAND2X1 NAND2X1_680 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe35), .B(_5503_), .Y(_5530_) );
OAI21X1 OAI21X1_1563 ( .gnd(gnd), .vdd(vdd), .A(_5529_), .B(micro_hash_ucr_2_pipe35), .C(_5530_), .Y(_5531_) );
OAI21X1 OAI21X1_1564 ( .gnd(gnd), .vdd(vdd), .A(_5104__bF_buf1), .B(micro_hash_ucr_2_a_3_), .C(_5106_), .Y(_5532_) );
AOI21X1 AOI21X1_998 ( .gnd(gnd), .vdd(vdd), .A(_5104__bF_buf0), .B(_5531_), .C(_5532_), .Y(_5533_) );
OAI21X1 OAI21X1_1565 ( .gnd(gnd), .vdd(vdd), .A(_5503_), .B(_5106_), .C(_5105__bF_buf1), .Y(_5534_) );
OAI22X1 OAI22X1_78 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_3_), .B(_5105__bF_buf0), .C(_5533_), .D(_5534_), .Y(_5535_) );
NAND2X1 NAND2X1_681 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe39), .B(_5487__bF_buf2), .Y(_5536_) );
OAI21X1 OAI21X1_1566 ( .gnd(gnd), .vdd(vdd), .A(_5535_), .B(micro_hash_ucr_2_pipe39), .C(_5536_), .Y(_5537_) );
NAND2X1 NAND2X1_682 ( .gnd(gnd), .vdd(vdd), .A(_5103__bF_buf1), .B(_5537_), .Y(_5538_) );
AOI21X1 AOI21X1_999 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_3_), .B(micro_hash_ucr_2_pipe40_bF_buf3), .C(micro_hash_ucr_2_pipe41_bF_buf2), .Y(_5539_) );
OAI21X1 OAI21X1_1567 ( .gnd(gnd), .vdd(vdd), .A(_5487__bF_buf1), .B(_5102_), .C(_5098__bF_buf1), .Y(_5540_) );
AOI21X1 AOI21X1_1000 ( .gnd(gnd), .vdd(vdd), .A(_5539_), .B(_5538_), .C(_5540_), .Y(_5541_) );
NOR2X1 NOR2X1_973 ( .gnd(gnd), .vdd(vdd), .A(_4654__bF_buf1), .B(_5098__bF_buf0), .Y(_5542_) );
OAI21X1 OAI21X1_1568 ( .gnd(gnd), .vdd(vdd), .A(_5541_), .B(_5542_), .C(_5100__bF_buf2), .Y(_5543_) );
NAND2X1 NAND2X1_683 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe43), .B(_5487__bF_buf0), .Y(_5544_) );
NAND3X1 NAND3X1_195 ( .gnd(gnd), .vdd(vdd), .A(_5099__bF_buf4), .B(_5544_), .C(_5543_), .Y(_5545_) );
NAND3X1 NAND3X1_196 ( .gnd(gnd), .vdd(vdd), .A(_5095_), .B(_5484_), .C(_5545_), .Y(_5546_) );
NAND2X1 NAND2X1_684 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe45_bF_buf2), .B(_5487__bF_buf3), .Y(_5547_) );
NAND3X1 NAND3X1_197 ( .gnd(gnd), .vdd(vdd), .A(_5097__bF_buf1), .B(_5547_), .C(_5546_), .Y(_5548_) );
NAND3X1 NAND3X1_198 ( .gnd(gnd), .vdd(vdd), .A(_5096__bF_buf0), .B(_5483_), .C(_5548_), .Y(_5549_) );
NAND2X1 NAND2X1_685 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe47), .B(_5487__bF_buf2), .Y(_5550_) );
NAND3X1 NAND3X1_199 ( .gnd(gnd), .vdd(vdd), .A(_5092__bF_buf1), .B(_5550_), .C(_5549_), .Y(_5551_) );
NAND3X1 NAND3X1_200 ( .gnd(gnd), .vdd(vdd), .A(_5094_), .B(_5482_), .C(_5551_), .Y(_5552_) );
NAND2X1 NAND2X1_686 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe49_bF_buf2), .B(_5487__bF_buf1), .Y(_5553_) );
NAND3X1 NAND3X1_201 ( .gnd(gnd), .vdd(vdd), .A(_5093__bF_buf2), .B(_5553_), .C(_5552_), .Y(_5554_) );
NAND3X1 NAND3X1_202 ( .gnd(gnd), .vdd(vdd), .A(_5089__bF_buf0), .B(_5481_), .C(_5554_), .Y(_5555_) );
NAND2X1 NAND2X1_687 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe51), .B(_5487__bF_buf0), .Y(_5556_) );
NAND3X1 NAND3X1_203 ( .gnd(gnd), .vdd(vdd), .A(_5091__bF_buf1), .B(_5556_), .C(_5555_), .Y(_5557_) );
NAND3X1 NAND3X1_204 ( .gnd(gnd), .vdd(vdd), .A(_5090_), .B(_5480_), .C(_5557_), .Y(_5558_) );
NAND2X1 NAND2X1_688 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe53_bF_buf2), .B(_5487__bF_buf3), .Y(_5559_) );
NAND3X1 NAND3X1_205 ( .gnd(gnd), .vdd(vdd), .A(_5086__bF_buf0), .B(_5559_), .C(_5558_), .Y(_5560_) );
NAND3X1 NAND3X1_206 ( .gnd(gnd), .vdd(vdd), .A(_5088_), .B(_5479_), .C(_5560_), .Y(_5561_) );
NAND2X1 NAND2X1_689 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe55), .B(_5487__bF_buf2), .Y(_5562_) );
AOI21X1 AOI21X1_1001 ( .gnd(gnd), .vdd(vdd), .A(_5562_), .B(_5561_), .C(micro_hash_ucr_2_pipe56_bF_buf2), .Y(_5563_) );
OAI21X1 OAI21X1_1569 ( .gnd(gnd), .vdd(vdd), .A(_4654__bF_buf0), .B(_5087__bF_buf1), .C(_5083_), .Y(_5564_) );
AOI21X1 AOI21X1_1002 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe57_bF_buf2), .B(_5503_), .C(micro_hash_ucr_2_pipe58_bF_buf3), .Y(_5565_) );
OAI21X1 OAI21X1_1570 ( .gnd(gnd), .vdd(vdd), .A(_5563_), .B(_5564_), .C(_5565_), .Y(_5566_) );
OAI21X1 OAI21X1_1571 ( .gnd(gnd), .vdd(vdd), .A(_4654__bF_buf3), .B(_5085__bF_buf1), .C(_5566_), .Y(_5567_) );
OAI21X1 OAI21X1_1572 ( .gnd(gnd), .vdd(vdd), .A(_5503_), .B(_5084__bF_buf2), .C(_5080__bF_buf0), .Y(_5568_) );
AOI21X1 AOI21X1_1003 ( .gnd(gnd), .vdd(vdd), .A(_5084__bF_buf1), .B(_5567_), .C(_5568_), .Y(_5569_) );
OAI21X1 OAI21X1_1573 ( .gnd(gnd), .vdd(vdd), .A(_5080__bF_buf3), .B(micro_hash_ucr_2_a_3_), .C(_5082_), .Y(_5570_) );
AOI21X1 AOI21X1_1004 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe61_bF_buf2), .B(_5487__bF_buf1), .C(micro_hash_ucr_2_pipe62_bF_buf1), .Y(_5571_) );
OAI21X1 OAI21X1_1574 ( .gnd(gnd), .vdd(vdd), .A(_5569_), .B(_5570_), .C(_5571_), .Y(_5572_) );
NAND2X1 NAND2X1_690 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe62_bF_buf0), .B(_4654__bF_buf2), .Y(_5573_) );
AOI21X1 AOI21X1_1005 ( .gnd(gnd), .vdd(vdd), .A(_5573_), .B(_5572_), .C(micro_hash_ucr_2_pipe63), .Y(_5574_) );
NOR2X1 NOR2X1_974 ( .gnd(gnd), .vdd(vdd), .A(_5077__bF_buf3), .B(_5487__bF_buf0), .Y(_5575_) );
OAI21X1 OAI21X1_1575 ( .gnd(gnd), .vdd(vdd), .A(_5574_), .B(_5575_), .C(_5079__bF_buf4), .Y(_5576_) );
NAND3X1 NAND3X1_207 ( .gnd(gnd), .vdd(vdd), .A(_5078_), .B(_5478_), .C(_5576_), .Y(_5577_) );
AOI21X1 AOI21X1_1006 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe65_bF_buf0), .B(_5487__bF_buf3), .C(micro_hash_ucr_2_pipe66_bF_buf4), .Y(_5578_) );
OAI21X1 OAI21X1_1576 ( .gnd(gnd), .vdd(vdd), .A(_5074__bF_buf0), .B(micro_hash_ucr_2_a_3_), .C(_5076__bF_buf3), .Y(_5579_) );
AOI21X1 AOI21X1_1007 ( .gnd(gnd), .vdd(vdd), .A(_5578_), .B(_5577_), .C(_5579_), .Y(_5580_) );
OAI21X1 OAI21X1_1577 ( .gnd(gnd), .vdd(vdd), .A(_5503_), .B(_5076__bF_buf2), .C(_5075__bF_buf0), .Y(_5581_) );
OAI22X1 OAI22X1_79 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_3_), .B(_5075__bF_buf4), .C(_5580_), .D(_5581_), .Y(_5582_) );
OAI21X1 OAI21X1_1578 ( .gnd(gnd), .vdd(vdd), .A(_5487__bF_buf2), .B(_5073__bF_buf1), .C(_4496__bF_buf2), .Y(_5583_) );
AOI21X1 AOI21X1_1008 ( .gnd(gnd), .vdd(vdd), .A(_5073__bF_buf0), .B(_5582_), .C(_5583_), .Y(_4491__3_) );
NAND2X1 NAND2X1_691 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe64_bF_buf0), .B(_4668__bF_buf2), .Y(_5584_) );
NAND2X1 NAND2X1_692 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe48_bF_buf3), .B(_4668__bF_buf1), .Y(_5585_) );
NOR2X1 NOR2X1_975 ( .gnd(gnd), .vdd(vdd), .A(_4668__bF_buf0), .B(_5097__bF_buf0), .Y(_5586_) );
NAND2X1 NAND2X1_693 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe36_bF_buf2), .B(_4668__bF_buf3), .Y(_5587_) );
NAND2X1 NAND2X1_694 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe34_bF_buf2), .B(_4668__bF_buf2), .Y(_5588_) );
NAND2X1 NAND2X1_695 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe32_bF_buf2), .B(_4668__bF_buf1), .Y(_5589_) );
NAND2X1 NAND2X1_696 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_4_), .B(micro_hash_ucr_2_pipe22_bF_buf2), .Y(_5590_) );
NAND2X1 NAND2X1_697 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_4_), .B(micro_hash_ucr_2_pipe20_bF_buf3), .Y(_5591_) );
INVX1 INVX1_368 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_4_), .Y(_5592_) );
INVX8 INVX8_178 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_4_bF_buf1_), .Y(_5593_) );
NAND2X1 NAND2X1_698 ( .gnd(gnd), .vdd(vdd), .A(_5592_), .B(_5593_), .Y(_5594_) );
NAND2X1 NAND2X1_699 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_4_), .B(micro_hash_ucr_2_b_4_bF_buf0_), .Y(_5595_) );
NAND2X1 NAND2X1_700 ( .gnd(gnd), .vdd(vdd), .A(_5595_), .B(_5594_), .Y(_5596_) );
NOR2X1 NOR2X1_976 ( .gnd(gnd), .vdd(vdd), .A(_5126_), .B(_5596_), .Y(_5597_) );
INVX8 INVX8_179 ( .gnd(gnd), .vdd(vdd), .A(_5596_), .Y(_5598_) );
NAND3X1 NAND3X1_208 ( .gnd(gnd), .vdd(vdd), .A(_4665_), .B(_5131_), .C(_5136_), .Y(_5599_) );
OAI22X1 OAI22X1_80 ( .gnd(gnd), .vdd(vdd), .A(_5495_), .B(_5599_), .C(_5269_), .D(_5598__bF_buf3), .Y(_5600_) );
AND2X2 AND2X2_427 ( .gnd(gnd), .vdd(vdd), .A(_5600_), .B(_5129_), .Y(_5601_) );
OAI21X1 OAI21X1_1579 ( .gnd(gnd), .vdd(vdd), .A(_5278_), .B(micro_hash_ucr_2_a_4_), .C(_5125__bF_buf2), .Y(_5602_) );
OAI22X1 OAI22X1_81 ( .gnd(gnd), .vdd(vdd), .A(_5125__bF_buf1), .B(_5596_), .C(_5601_), .D(_5602_), .Y(_5603_) );
NAND2X1 NAND2X1_701 ( .gnd(gnd), .vdd(vdd), .A(_5127__bF_buf2), .B(_5603_), .Y(_5604_) );
OAI21X1 OAI21X1_1580 ( .gnd(gnd), .vdd(vdd), .A(_4668__bF_buf0), .B(_5127__bF_buf1), .C(_5604_), .Y(_5605_) );
AND2X2 AND2X2_428 ( .gnd(gnd), .vdd(vdd), .A(_5605_), .B(_5126_), .Y(_5606_) );
OAI21X1 OAI21X1_1581 ( .gnd(gnd), .vdd(vdd), .A(_5606_), .B(_5597_), .C(_5122__bF_buf1), .Y(_5607_) );
OAI21X1 OAI21X1_1582 ( .gnd(gnd), .vdd(vdd), .A(_4668__bF_buf3), .B(_5122__bF_buf0), .C(_5607_), .Y(_5608_) );
AND2X2 AND2X2_429 ( .gnd(gnd), .vdd(vdd), .A(_5608_), .B(_5124__bF_buf3), .Y(_5609_) );
NOR2X1 NOR2X1_977 ( .gnd(gnd), .vdd(vdd), .A(_5124__bF_buf2), .B(_5596_), .Y(_5610_) );
OAI21X1 OAI21X1_1583 ( .gnd(gnd), .vdd(vdd), .A(_5609_), .B(_5610_), .C(_5123__bF_buf2), .Y(_5611_) );
AOI21X1 AOI21X1_1009 ( .gnd(gnd), .vdd(vdd), .A(_5591_), .B(_5611_), .C(micro_hash_ucr_2_pipe21_bF_buf0), .Y(_5612_) );
NOR2X1 NOR2X1_978 ( .gnd(gnd), .vdd(vdd), .A(_5119_), .B(_5596_), .Y(_5613_) );
OAI21X1 OAI21X1_1584 ( .gnd(gnd), .vdd(vdd), .A(_5612_), .B(_5613_), .C(_5121__bF_buf0), .Y(_5614_) );
AOI21X1 AOI21X1_1010 ( .gnd(gnd), .vdd(vdd), .A(_5590_), .B(_5614_), .C(micro_hash_ucr_2_pipe23), .Y(_5615_) );
OAI21X1 OAI21X1_1585 ( .gnd(gnd), .vdd(vdd), .A(_5596_), .B(_5120__bF_buf1), .C(_5116__bF_buf4), .Y(_5616_) );
AOI21X1 AOI21X1_1011 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe24_bF_buf1), .B(_4668__bF_buf2), .C(micro_hash_ucr_2_pipe25), .Y(_5617_) );
OAI21X1 OAI21X1_1586 ( .gnd(gnd), .vdd(vdd), .A(_5615_), .B(_5616_), .C(_5617_), .Y(_5618_) );
AOI21X1 AOI21X1_1012 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe25), .B(_5598__bF_buf2), .C(micro_hash_ucr_2_pipe26_bF_buf3), .Y(_5619_) );
AOI22X1 AOI22X1_47 ( .gnd(gnd), .vdd(vdd), .A(_4668__bF_buf1), .B(micro_hash_ucr_2_pipe26_bF_buf2), .C(_5618_), .D(_5619_), .Y(_5620_) );
OAI21X1 OAI21X1_1587 ( .gnd(gnd), .vdd(vdd), .A(_5596_), .B(_5113_), .C(_5115__bF_buf3), .Y(_5621_) );
AOI21X1 AOI21X1_1013 ( .gnd(gnd), .vdd(vdd), .A(_5113_), .B(_5620_), .C(_5621_), .Y(_5622_) );
OAI21X1 OAI21X1_1588 ( .gnd(gnd), .vdd(vdd), .A(_5115__bF_buf2), .B(micro_hash_ucr_2_a_4_), .C(_5114_), .Y(_5623_) );
AOI21X1 AOI21X1_1014 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe29_bF_buf0), .B(_5598__bF_buf1), .C(micro_hash_ucr_2_pipe30_bF_buf0), .Y(_5624_) );
OAI21X1 OAI21X1_1589 ( .gnd(gnd), .vdd(vdd), .A(_5622_), .B(_5623_), .C(_5624_), .Y(_5625_) );
NAND2X1 NAND2X1_702 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe30_bF_buf4), .B(_4668__bF_buf0), .Y(_5626_) );
AOI21X1 AOI21X1_1015 ( .gnd(gnd), .vdd(vdd), .A(_5626_), .B(_5625_), .C(micro_hash_ucr_2_pipe31), .Y(_5627_) );
NOR2X1 NOR2X1_979 ( .gnd(gnd), .vdd(vdd), .A(_5112__bF_buf0), .B(_5598__bF_buf0), .Y(_5628_) );
OAI21X1 OAI21X1_1590 ( .gnd(gnd), .vdd(vdd), .A(_5627_), .B(_5628_), .C(_5111__bF_buf0), .Y(_5629_) );
AOI21X1 AOI21X1_1016 ( .gnd(gnd), .vdd(vdd), .A(_5589_), .B(_5629_), .C(micro_hash_ucr_2_pipe33_bF_buf2), .Y(_5630_) );
NOR2X1 NOR2X1_980 ( .gnd(gnd), .vdd(vdd), .A(_5107_), .B(_5598__bF_buf3), .Y(_5631_) );
OAI21X1 OAI21X1_1591 ( .gnd(gnd), .vdd(vdd), .A(_5630_), .B(_5631_), .C(_5109__bF_buf4), .Y(_5632_) );
AOI21X1 AOI21X1_1017 ( .gnd(gnd), .vdd(vdd), .A(_5588_), .B(_5632_), .C(micro_hash_ucr_2_pipe35), .Y(_5633_) );
NOR2X1 NOR2X1_981 ( .gnd(gnd), .vdd(vdd), .A(_5108__bF_buf2), .B(_5598__bF_buf2), .Y(_5634_) );
OAI21X1 OAI21X1_1592 ( .gnd(gnd), .vdd(vdd), .A(_5633_), .B(_5634_), .C(_5104__bF_buf4), .Y(_5635_) );
NAND3X1 NAND3X1_209 ( .gnd(gnd), .vdd(vdd), .A(_5106_), .B(_5587_), .C(_5635_), .Y(_5636_) );
AOI21X1 AOI21X1_1018 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe37), .B(_5598__bF_buf1), .C(micro_hash_ucr_2_pipe38_bF_buf2), .Y(_5637_) );
OAI21X1 OAI21X1_1593 ( .gnd(gnd), .vdd(vdd), .A(_5105__bF_buf4), .B(micro_hash_ucr_2_a_4_), .C(_5101_), .Y(_5638_) );
AOI21X1 AOI21X1_1019 ( .gnd(gnd), .vdd(vdd), .A(_5637_), .B(_5636_), .C(_5638_), .Y(_5639_) );
OAI21X1 OAI21X1_1594 ( .gnd(gnd), .vdd(vdd), .A(_5596_), .B(_5101_), .C(_5103__bF_buf0), .Y(_5640_) );
OAI22X1 OAI22X1_82 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_4_), .B(_5103__bF_buf3), .C(_5639_), .D(_5640_), .Y(_5641_) );
NAND2X1 NAND2X1_703 ( .gnd(gnd), .vdd(vdd), .A(_5102_), .B(_5641_), .Y(_5642_) );
NAND2X1 NAND2X1_704 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe41_bF_buf1), .B(_5596_), .Y(_5643_) );
NAND3X1 NAND3X1_210 ( .gnd(gnd), .vdd(vdd), .A(_5098__bF_buf4), .B(_5643_), .C(_5642_), .Y(_5644_) );
AOI21X1 AOI21X1_1020 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_4_), .B(micro_hash_ucr_2_pipe42_bF_buf2), .C(micro_hash_ucr_2_pipe43), .Y(_5645_) );
OAI21X1 OAI21X1_1595 ( .gnd(gnd), .vdd(vdd), .A(_5598__bF_buf0), .B(_5100__bF_buf1), .C(_5099__bF_buf3), .Y(_5646_) );
AOI21X1 AOI21X1_1021 ( .gnd(gnd), .vdd(vdd), .A(_5645_), .B(_5644_), .C(_5646_), .Y(_5647_) );
NOR2X1 NOR2X1_982 ( .gnd(gnd), .vdd(vdd), .A(_4668__bF_buf3), .B(_5099__bF_buf2), .Y(_5648_) );
OAI21X1 OAI21X1_1596 ( .gnd(gnd), .vdd(vdd), .A(_5647_), .B(_5648_), .C(_5095_), .Y(_5649_) );
NAND2X1 NAND2X1_705 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe45_bF_buf1), .B(_5598__bF_buf3), .Y(_5650_) );
AOI21X1 AOI21X1_1022 ( .gnd(gnd), .vdd(vdd), .A(_5650_), .B(_5649_), .C(micro_hash_ucr_2_pipe46_bF_buf2), .Y(_5651_) );
OAI21X1 OAI21X1_1597 ( .gnd(gnd), .vdd(vdd), .A(_5651_), .B(_5586_), .C(_5096__bF_buf3), .Y(_5652_) );
NAND2X1 NAND2X1_706 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe47), .B(_5598__bF_buf2), .Y(_5653_) );
NAND3X1 NAND3X1_211 ( .gnd(gnd), .vdd(vdd), .A(_5092__bF_buf0), .B(_5653_), .C(_5652_), .Y(_5654_) );
NAND3X1 NAND3X1_212 ( .gnd(gnd), .vdd(vdd), .A(_5094_), .B(_5585_), .C(_5654_), .Y(_5655_) );
AOI21X1 AOI21X1_1023 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe49_bF_buf1), .B(_5598__bF_buf1), .C(micro_hash_ucr_2_pipe50_bF_buf0), .Y(_5656_) );
OAI21X1 OAI21X1_1598 ( .gnd(gnd), .vdd(vdd), .A(_5093__bF_buf1), .B(micro_hash_ucr_2_a_4_), .C(_5089__bF_buf3), .Y(_5657_) );
AOI21X1 AOI21X1_1024 ( .gnd(gnd), .vdd(vdd), .A(_5656_), .B(_5655_), .C(_5657_), .Y(_5658_) );
OAI21X1 OAI21X1_1599 ( .gnd(gnd), .vdd(vdd), .A(_5596_), .B(_5089__bF_buf2), .C(_5091__bF_buf0), .Y(_5659_) );
OAI22X1 OAI22X1_83 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_4_), .B(_5091__bF_buf4), .C(_5658_), .D(_5659_), .Y(_5660_) );
NAND2X1 NAND2X1_707 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe53_bF_buf1), .B(_5598__bF_buf0), .Y(_5661_) );
OAI21X1 OAI21X1_1600 ( .gnd(gnd), .vdd(vdd), .A(_5660_), .B(micro_hash_ucr_2_pipe53_bF_buf0), .C(_5661_), .Y(_5662_) );
NAND2X1 NAND2X1_708 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe54_bF_buf3), .B(_4668__bF_buf2), .Y(_5663_) );
OAI21X1 OAI21X1_1601 ( .gnd(gnd), .vdd(vdd), .A(_5662_), .B(micro_hash_ucr_2_pipe54_bF_buf2), .C(_5663_), .Y(_5664_) );
NAND2X1 NAND2X1_709 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe55), .B(_5598__bF_buf3), .Y(_5665_) );
OAI21X1 OAI21X1_1602 ( .gnd(gnd), .vdd(vdd), .A(_5664_), .B(micro_hash_ucr_2_pipe55), .C(_5665_), .Y(_5666_) );
OAI21X1 OAI21X1_1603 ( .gnd(gnd), .vdd(vdd), .A(_4668__bF_buf1), .B(_5087__bF_buf0), .C(_5083_), .Y(_5667_) );
AOI21X1 AOI21X1_1025 ( .gnd(gnd), .vdd(vdd), .A(_5087__bF_buf4), .B(_5666_), .C(_5667_), .Y(_5668_) );
OAI21X1 OAI21X1_1604 ( .gnd(gnd), .vdd(vdd), .A(_5598__bF_buf2), .B(_5083_), .C(_5085__bF_buf0), .Y(_5669_) );
OAI22X1 OAI22X1_84 ( .gnd(gnd), .vdd(vdd), .A(_4668__bF_buf0), .B(_5085__bF_buf3), .C(_5668_), .D(_5669_), .Y(_5670_) );
OAI21X1 OAI21X1_1605 ( .gnd(gnd), .vdd(vdd), .A(_5596_), .B(_5084__bF_buf0), .C(_5080__bF_buf2), .Y(_5671_) );
AOI21X1 AOI21X1_1026 ( .gnd(gnd), .vdd(vdd), .A(_5084__bF_buf3), .B(_5670_), .C(_5671_), .Y(_5672_) );
OAI21X1 OAI21X1_1606 ( .gnd(gnd), .vdd(vdd), .A(_5080__bF_buf1), .B(micro_hash_ucr_2_a_4_), .C(_5082_), .Y(_5673_) );
AOI21X1 AOI21X1_1027 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe61_bF_buf1), .B(_5598__bF_buf1), .C(micro_hash_ucr_2_pipe62_bF_buf4), .Y(_5674_) );
OAI21X1 OAI21X1_1607 ( .gnd(gnd), .vdd(vdd), .A(_5672_), .B(_5673_), .C(_5674_), .Y(_5675_) );
NAND2X1 NAND2X1_710 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe62_bF_buf3), .B(_4668__bF_buf3), .Y(_5676_) );
AOI21X1 AOI21X1_1028 ( .gnd(gnd), .vdd(vdd), .A(_5676_), .B(_5675_), .C(micro_hash_ucr_2_pipe63), .Y(_5677_) );
NOR2X1 NOR2X1_983 ( .gnd(gnd), .vdd(vdd), .A(_5077__bF_buf2), .B(_5598__bF_buf0), .Y(_5678_) );
OAI21X1 OAI21X1_1608 ( .gnd(gnd), .vdd(vdd), .A(_5677_), .B(_5678_), .C(_5079__bF_buf3), .Y(_5679_) );
NAND3X1 NAND3X1_213 ( .gnd(gnd), .vdd(vdd), .A(_5078_), .B(_5584_), .C(_5679_), .Y(_5680_) );
NAND2X1 NAND2X1_711 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe65_bF_buf3), .B(_5598__bF_buf3), .Y(_5681_) );
AOI21X1 AOI21X1_1029 ( .gnd(gnd), .vdd(vdd), .A(_5681_), .B(_5680_), .C(micro_hash_ucr_2_pipe66_bF_buf3), .Y(_5682_) );
OAI21X1 OAI21X1_1609 ( .gnd(gnd), .vdd(vdd), .A(_4668__bF_buf2), .B(_5074__bF_buf3), .C(_5076__bF_buf1), .Y(_5683_) );
AOI21X1 AOI21X1_1030 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe67), .B(_5596_), .C(micro_hash_ucr_2_pipe68), .Y(_5684_) );
OAI21X1 OAI21X1_1610 ( .gnd(gnd), .vdd(vdd), .A(_5682_), .B(_5683_), .C(_5684_), .Y(_5685_) );
AOI21X1 AOI21X1_1031 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_4_), .B(micro_hash_ucr_2_pipe68), .C(micro_hash_ucr_2_pipe69), .Y(_5686_) );
OAI21X1 OAI21X1_1611 ( .gnd(gnd), .vdd(vdd), .A(_5598__bF_buf2), .B(_5073__bF_buf3), .C(_4496__bF_buf1), .Y(_5687_) );
AOI21X1 AOI21X1_1032 ( .gnd(gnd), .vdd(vdd), .A(_5686_), .B(_5685_), .C(_5687_), .Y(_4491__4_) );
NAND2X1 NAND2X1_712 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_5_bF_buf1_), .B(micro_hash_ucr_2_pipe66_bF_buf2), .Y(_5688_) );
NAND2X1 NAND2X1_713 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_5_bF_buf0_), .B(micro_hash_ucr_2_pipe64_bF_buf4), .Y(_5689_) );
NAND2X1 NAND2X1_714 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_5_bF_buf3_), .B(micro_hash_ucr_2_pipe62_bF_buf2), .Y(_5690_) );
NAND2X1 NAND2X1_715 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_5_bF_buf2_), .B(micro_hash_ucr_2_pipe54_bF_buf1), .Y(_5691_) );
NAND2X1 NAND2X1_716 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_5_bF_buf1_), .B(micro_hash_ucr_2_pipe42_bF_buf1), .Y(_5692_) );
NAND2X1 NAND2X1_717 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_5_bF_buf0_), .B(micro_hash_ucr_2_pipe40_bF_buf2), .Y(_5693_) );
NAND2X1 NAND2X1_718 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe34_bF_buf1), .B(_4674__bF_buf2), .Y(_5694_) );
NAND2X1 NAND2X1_719 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe32_bF_buf1), .B(_4674__bF_buf1), .Y(_5695_) );
NAND2X1 NAND2X1_720 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe30_bF_buf3), .B(_4674__bF_buf0), .Y(_5696_) );
NAND2X1 NAND2X1_721 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe22_bF_buf1), .B(_4674__bF_buf3), .Y(_5697_) );
NAND2X1 NAND2X1_722 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe20_bF_buf2), .B(_4674__bF_buf2), .Y(_5698_) );
NAND2X1 NAND2X1_723 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe18_bF_buf1), .B(_4674__bF_buf1), .Y(_5699_) );
NAND2X1 NAND2X1_724 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe16_bF_buf3), .B(_4674__bF_buf0), .Y(_5700_) );
NAND2X1 NAND2X1_725 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe14_bF_buf1), .B(_4674__bF_buf3), .Y(_5701_) );
NOR2X1 NOR2X1_984 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_5_), .B(micro_hash_ucr_2_b_5_bF_buf1_), .Y(_5702_) );
NAND2X1 NAND2X1_726 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_5_), .B(micro_hash_ucr_2_b_5_bF_buf0_), .Y(_5703_) );
INVX4 INVX4_104 ( .gnd(gnd), .vdd(vdd), .A(_5703_), .Y(_5704_) );
NOR2X1 NOR2X1_985 ( .gnd(gnd), .vdd(vdd), .A(_5702_), .B(_5704_), .Y(_5705_) );
NAND2X1 NAND2X1_727 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe13), .B(_5705__bF_buf3), .Y(_5706_) );
NOR2X1 NOR2X1_986 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe13), .B(_5128_), .Y(_5707_) );
NAND2X1 NAND2X1_728 ( .gnd(gnd), .vdd(vdd), .A(_4674__bF_buf2), .B(_5160_), .Y(_5708_) );
INVX4 INVX4_105 ( .gnd(gnd), .vdd(vdd), .A(_5705__bF_buf2), .Y(_5709_) );
NOR2X1 NOR2X1_987 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe9), .B(micro_hash_ucr_2_pipe10), .Y(_5710_) );
INVX1 INVX1_369 ( .gnd(gnd), .vdd(vdd), .A(_5710_), .Y(_5711_) );
NAND3X1 NAND3X1_214 ( .gnd(gnd), .vdd(vdd), .A(_4673_), .B(_5132_), .C(_5136_), .Y(_5712_) );
NOR3X1 NOR3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_5711_), .B(_5158_), .C(_5712_), .Y(_5713_) );
NAND2X1 NAND2X1_729 ( .gnd(gnd), .vdd(vdd), .A(_5133_), .B(_5171_), .Y(_5714_) );
NAND3X1 NAND3X1_215 ( .gnd(gnd), .vdd(vdd), .A(_5130_), .B(_5132_), .C(_5714_), .Y(_5715_) );
AOI21X1 AOI21X1_1033 ( .gnd(gnd), .vdd(vdd), .A(_5709_), .B(_5715_), .C(_5713_), .Y(_5716_) );
OAI21X1 OAI21X1_1612 ( .gnd(gnd), .vdd(vdd), .A(_5716_), .B(_5707_), .C(_5708_), .Y(_5717_) );
NAND3X1 NAND3X1_216 ( .gnd(gnd), .vdd(vdd), .A(_5129_), .B(_5706_), .C(_5717_), .Y(_5718_) );
NAND3X1 NAND3X1_217 ( .gnd(gnd), .vdd(vdd), .A(_5125__bF_buf0), .B(_5701_), .C(_5718_), .Y(_5719_) );
NAND2X1 NAND2X1_730 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe15), .B(_5705__bF_buf1), .Y(_5720_) );
NAND3X1 NAND3X1_218 ( .gnd(gnd), .vdd(vdd), .A(_5127__bF_buf0), .B(_5720_), .C(_5719_), .Y(_5721_) );
NAND3X1 NAND3X1_219 ( .gnd(gnd), .vdd(vdd), .A(_5126_), .B(_5700_), .C(_5721_), .Y(_5722_) );
NAND2X1 NAND2X1_731 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe17_bF_buf2), .B(_5705__bF_buf0), .Y(_5723_) );
NAND3X1 NAND3X1_220 ( .gnd(gnd), .vdd(vdd), .A(_5122__bF_buf4), .B(_5723_), .C(_5722_), .Y(_5724_) );
NAND3X1 NAND3X1_221 ( .gnd(gnd), .vdd(vdd), .A(_5124__bF_buf1), .B(_5699_), .C(_5724_), .Y(_5725_) );
NAND2X1 NAND2X1_732 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe19), .B(_5705__bF_buf3), .Y(_5726_) );
NAND3X1 NAND3X1_222 ( .gnd(gnd), .vdd(vdd), .A(_5123__bF_buf1), .B(_5726_), .C(_5725_), .Y(_5727_) );
NAND3X1 NAND3X1_223 ( .gnd(gnd), .vdd(vdd), .A(_5119_), .B(_5698_), .C(_5727_), .Y(_5728_) );
NAND2X1 NAND2X1_733 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe21_bF_buf3), .B(_5705__bF_buf2), .Y(_5729_) );
NAND3X1 NAND3X1_224 ( .gnd(gnd), .vdd(vdd), .A(_5121__bF_buf4), .B(_5729_), .C(_5728_), .Y(_5730_) );
NAND3X1 NAND3X1_225 ( .gnd(gnd), .vdd(vdd), .A(_5120__bF_buf0), .B(_5697_), .C(_5730_), .Y(_5731_) );
AOI21X1 AOI21X1_1034 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe23), .B(_5705__bF_buf1), .C(micro_hash_ucr_2_pipe24_bF_buf0), .Y(_5732_) );
OAI21X1 OAI21X1_1613 ( .gnd(gnd), .vdd(vdd), .A(_5116__bF_buf3), .B(micro_hash_ucr_2_a_5_bF_buf3_), .C(_5118__bF_buf2), .Y(_5733_) );
AOI21X1 AOI21X1_1035 ( .gnd(gnd), .vdd(vdd), .A(_5732_), .B(_5731_), .C(_5733_), .Y(_5734_) );
OAI21X1 OAI21X1_1614 ( .gnd(gnd), .vdd(vdd), .A(_5709_), .B(_5118__bF_buf1), .C(_5117__bF_buf2), .Y(_5735_) );
NAND2X1 NAND2X1_734 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe26_bF_buf1), .B(_4674__bF_buf1), .Y(_5736_) );
OAI21X1 OAI21X1_1615 ( .gnd(gnd), .vdd(vdd), .A(_5734_), .B(_5735_), .C(_5736_), .Y(_5737_) );
OAI21X1 OAI21X1_1616 ( .gnd(gnd), .vdd(vdd), .A(_5705__bF_buf0), .B(_5113_), .C(_5115__bF_buf1), .Y(_5738_) );
AOI21X1 AOI21X1_1036 ( .gnd(gnd), .vdd(vdd), .A(_5113_), .B(_5737_), .C(_5738_), .Y(_5739_) );
NOR2X1 NOR2X1_988 ( .gnd(gnd), .vdd(vdd), .A(_4674__bF_buf0), .B(_5115__bF_buf0), .Y(_5740_) );
OAI21X1 OAI21X1_1617 ( .gnd(gnd), .vdd(vdd), .A(_5739_), .B(_5740_), .C(_5114_), .Y(_5741_) );
NAND2X1 NAND2X1_735 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe29_bF_buf3), .B(_5705__bF_buf3), .Y(_5742_) );
NAND3X1 NAND3X1_226 ( .gnd(gnd), .vdd(vdd), .A(_5110__bF_buf1), .B(_5742_), .C(_5741_), .Y(_5743_) );
NAND3X1 NAND3X1_227 ( .gnd(gnd), .vdd(vdd), .A(_5112__bF_buf3), .B(_5696_), .C(_5743_), .Y(_5744_) );
NAND2X1 NAND2X1_736 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe31), .B(_5705__bF_buf2), .Y(_5745_) );
NAND3X1 NAND3X1_228 ( .gnd(gnd), .vdd(vdd), .A(_5111__bF_buf4), .B(_5745_), .C(_5744_), .Y(_5746_) );
NAND3X1 NAND3X1_229 ( .gnd(gnd), .vdd(vdd), .A(_5107_), .B(_5695_), .C(_5746_), .Y(_5747_) );
NAND2X1 NAND2X1_737 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe33_bF_buf1), .B(_5705__bF_buf1), .Y(_5748_) );
NAND3X1 NAND3X1_230 ( .gnd(gnd), .vdd(vdd), .A(_5109__bF_buf3), .B(_5748_), .C(_5747_), .Y(_5749_) );
NAND3X1 NAND3X1_231 ( .gnd(gnd), .vdd(vdd), .A(_5108__bF_buf1), .B(_5694_), .C(_5749_), .Y(_5750_) );
NAND2X1 NAND2X1_738 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe35), .B(_5705__bF_buf0), .Y(_5751_) );
AOI21X1 AOI21X1_1037 ( .gnd(gnd), .vdd(vdd), .A(_5751_), .B(_5750_), .C(micro_hash_ucr_2_pipe36_bF_buf1), .Y(_5752_) );
OAI21X1 OAI21X1_1618 ( .gnd(gnd), .vdd(vdd), .A(_4674__bF_buf3), .B(_5104__bF_buf3), .C(_5106_), .Y(_5753_) );
AOI21X1 AOI21X1_1038 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe37), .B(_5709_), .C(micro_hash_ucr_2_pipe38_bF_buf1), .Y(_5754_) );
OAI21X1 OAI21X1_1619 ( .gnd(gnd), .vdd(vdd), .A(_5752_), .B(_5753_), .C(_5754_), .Y(_5755_) );
NAND2X1 NAND2X1_739 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_5_bF_buf2_), .B(micro_hash_ucr_2_pipe38_bF_buf0), .Y(_5756_) );
NAND3X1 NAND3X1_232 ( .gnd(gnd), .vdd(vdd), .A(_5101_), .B(_5756_), .C(_5755_), .Y(_5757_) );
OAI21X1 OAI21X1_1620 ( .gnd(gnd), .vdd(vdd), .A(_5704_), .B(_5702_), .C(micro_hash_ucr_2_pipe39), .Y(_5758_) );
NAND3X1 NAND3X1_233 ( .gnd(gnd), .vdd(vdd), .A(_5103__bF_buf2), .B(_5758_), .C(_5757_), .Y(_5759_) );
NAND3X1 NAND3X1_234 ( .gnd(gnd), .vdd(vdd), .A(_5102_), .B(_5693_), .C(_5759_), .Y(_5760_) );
OAI21X1 OAI21X1_1621 ( .gnd(gnd), .vdd(vdd), .A(_5704_), .B(_5702_), .C(micro_hash_ucr_2_pipe41_bF_buf0), .Y(_5761_) );
NAND3X1 NAND3X1_235 ( .gnd(gnd), .vdd(vdd), .A(_5098__bF_buf3), .B(_5761_), .C(_5760_), .Y(_5762_) );
NAND3X1 NAND3X1_236 ( .gnd(gnd), .vdd(vdd), .A(_5100__bF_buf0), .B(_5692_), .C(_5762_), .Y(_5763_) );
OAI21X1 OAI21X1_1622 ( .gnd(gnd), .vdd(vdd), .A(_5704_), .B(_5702_), .C(micro_hash_ucr_2_pipe43), .Y(_5764_) );
NAND3X1 NAND3X1_237 ( .gnd(gnd), .vdd(vdd), .A(_5099__bF_buf1), .B(_5764_), .C(_5763_), .Y(_5765_) );
AOI21X1 AOI21X1_1039 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_5_bF_buf1_), .B(micro_hash_ucr_2_pipe44_bF_buf3), .C(micro_hash_ucr_2_pipe45_bF_buf0), .Y(_5766_) );
NOR2X1 NOR2X1_989 ( .gnd(gnd), .vdd(vdd), .A(_5095_), .B(_5705__bF_buf3), .Y(_5767_) );
AOI21X1 AOI21X1_1040 ( .gnd(gnd), .vdd(vdd), .A(_5766_), .B(_5765_), .C(_5767_), .Y(_5768_) );
AOI21X1 AOI21X1_1041 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe46_bF_buf1), .B(_4674__bF_buf2), .C(micro_hash_ucr_2_pipe47), .Y(_5769_) );
OAI21X1 OAI21X1_1623 ( .gnd(gnd), .vdd(vdd), .A(_5768_), .B(micro_hash_ucr_2_pipe46_bF_buf0), .C(_5769_), .Y(_5770_) );
AOI21X1 AOI21X1_1042 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe47), .B(_5705__bF_buf2), .C(micro_hash_ucr_2_pipe48_bF_buf2), .Y(_5771_) );
NAND2X1 NAND2X1_740 ( .gnd(gnd), .vdd(vdd), .A(_5771_), .B(_5770_), .Y(_5772_) );
NAND2X1 NAND2X1_741 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe48_bF_buf1), .B(_4674__bF_buf1), .Y(_5773_) );
NAND3X1 NAND3X1_238 ( .gnd(gnd), .vdd(vdd), .A(_5094_), .B(_5773_), .C(_5772_), .Y(_5774_) );
NAND2X1 NAND2X1_742 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe49_bF_buf0), .B(_5705__bF_buf1), .Y(_5775_) );
AOI21X1 AOI21X1_1043 ( .gnd(gnd), .vdd(vdd), .A(_5775_), .B(_5774_), .C(micro_hash_ucr_2_pipe50_bF_buf3), .Y(_5776_) );
OAI21X1 OAI21X1_1624 ( .gnd(gnd), .vdd(vdd), .A(_4674__bF_buf0), .B(_5093__bF_buf0), .C(_5089__bF_buf1), .Y(_5777_) );
AOI21X1 AOI21X1_1044 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe51), .B(_5709_), .C(micro_hash_ucr_2_pipe52_bF_buf1), .Y(_5778_) );
OAI21X1 OAI21X1_1625 ( .gnd(gnd), .vdd(vdd), .A(_5776_), .B(_5777_), .C(_5778_), .Y(_5779_) );
NAND2X1 NAND2X1_743 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_5_bF_buf0_), .B(micro_hash_ucr_2_pipe52_bF_buf0), .Y(_5780_) );
NAND3X1 NAND3X1_239 ( .gnd(gnd), .vdd(vdd), .A(_5090_), .B(_5780_), .C(_5779_), .Y(_5781_) );
OAI21X1 OAI21X1_1626 ( .gnd(gnd), .vdd(vdd), .A(_5704_), .B(_5702_), .C(micro_hash_ucr_2_pipe53_bF_buf3), .Y(_5782_) );
NAND3X1 NAND3X1_240 ( .gnd(gnd), .vdd(vdd), .A(_5086__bF_buf3), .B(_5782_), .C(_5781_), .Y(_5783_) );
AOI21X1 AOI21X1_1045 ( .gnd(gnd), .vdd(vdd), .A(_5691_), .B(_5783_), .C(micro_hash_ucr_2_pipe55), .Y(_5784_) );
OAI21X1 OAI21X1_1627 ( .gnd(gnd), .vdd(vdd), .A(_5709_), .B(_5088_), .C(_5087__bF_buf3), .Y(_5785_) );
AOI21X1 AOI21X1_1046 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe56_bF_buf1), .B(_4674__bF_buf3), .C(micro_hash_ucr_2_pipe57_bF_buf1), .Y(_5786_) );
OAI21X1 OAI21X1_1628 ( .gnd(gnd), .vdd(vdd), .A(_5784_), .B(_5785_), .C(_5786_), .Y(_5787_) );
AOI21X1 AOI21X1_1047 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe57_bF_buf0), .B(_5705__bF_buf0), .C(micro_hash_ucr_2_pipe58_bF_buf2), .Y(_5788_) );
NOR2X1 NOR2X1_990 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_5_bF_buf3_), .B(_5085__bF_buf2), .Y(_5789_) );
AOI21X1 AOI21X1_1048 ( .gnd(gnd), .vdd(vdd), .A(_5788_), .B(_5787_), .C(_5789_), .Y(_5790_) );
AOI21X1 AOI21X1_1049 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe59), .B(_5709_), .C(micro_hash_ucr_2_pipe60_bF_buf4), .Y(_5791_) );
OAI21X1 OAI21X1_1629 ( .gnd(gnd), .vdd(vdd), .A(_5790_), .B(micro_hash_ucr_2_pipe59), .C(_5791_), .Y(_5792_) );
NAND2X1 NAND2X1_744 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_5_bF_buf2_), .B(micro_hash_ucr_2_pipe60_bF_buf3), .Y(_5793_) );
NAND3X1 NAND3X1_241 ( .gnd(gnd), .vdd(vdd), .A(_5082_), .B(_5793_), .C(_5792_), .Y(_5794_) );
OAI21X1 OAI21X1_1630 ( .gnd(gnd), .vdd(vdd), .A(_5704_), .B(_5702_), .C(micro_hash_ucr_2_pipe61_bF_buf0), .Y(_5795_) );
NAND3X1 NAND3X1_242 ( .gnd(gnd), .vdd(vdd), .A(_5081__bF_buf2), .B(_5795_), .C(_5794_), .Y(_5796_) );
NAND3X1 NAND3X1_243 ( .gnd(gnd), .vdd(vdd), .A(_5077__bF_buf1), .B(_5690_), .C(_5796_), .Y(_5797_) );
OAI21X1 OAI21X1_1631 ( .gnd(gnd), .vdd(vdd), .A(_5704_), .B(_5702_), .C(micro_hash_ucr_2_pipe63), .Y(_5798_) );
NAND3X1 NAND3X1_244 ( .gnd(gnd), .vdd(vdd), .A(_5079__bF_buf2), .B(_5798_), .C(_5797_), .Y(_5799_) );
NAND3X1 NAND3X1_245 ( .gnd(gnd), .vdd(vdd), .A(_5078_), .B(_5689_), .C(_5799_), .Y(_5800_) );
OAI21X1 OAI21X1_1632 ( .gnd(gnd), .vdd(vdd), .A(_5704_), .B(_5702_), .C(micro_hash_ucr_2_pipe65_bF_buf2), .Y(_5801_) );
NAND3X1 NAND3X1_246 ( .gnd(gnd), .vdd(vdd), .A(_5074__bF_buf2), .B(_5801_), .C(_5800_), .Y(_5802_) );
NAND3X1 NAND3X1_247 ( .gnd(gnd), .vdd(vdd), .A(_5076__bF_buf0), .B(_5688_), .C(_5802_), .Y(_5803_) );
OAI21X1 OAI21X1_1633 ( .gnd(gnd), .vdd(vdd), .A(_5704_), .B(_5702_), .C(micro_hash_ucr_2_pipe67), .Y(_5804_) );
NAND3X1 NAND3X1_248 ( .gnd(gnd), .vdd(vdd), .A(_5075__bF_buf3), .B(_5804_), .C(_5803_), .Y(_5805_) );
AOI21X1 AOI21X1_1050 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_5_bF_buf1_), .B(micro_hash_ucr_2_pipe68), .C(micro_hash_ucr_2_pipe69), .Y(_5806_) );
OAI21X1 OAI21X1_1634 ( .gnd(gnd), .vdd(vdd), .A(_5705__bF_buf3), .B(_5073__bF_buf2), .C(_4496__bF_buf0), .Y(_5807_) );
AOI21X1 AOI21X1_1051 ( .gnd(gnd), .vdd(vdd), .A(_5806_), .B(_5805_), .C(_5807_), .Y(_4491__5_) );
NAND2X1 NAND2X1_745 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_6_bF_buf1_), .B(micro_hash_ucr_2_pipe66_bF_buf1), .Y(_5808_) );
NAND2X1 NAND2X1_746 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_6_bF_buf0_), .B(micro_hash_ucr_2_pipe64_bF_buf3), .Y(_5809_) );
NAND2X1 NAND2X1_747 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_6_bF_buf3_), .B(micro_hash_ucr_2_pipe62_bF_buf1), .Y(_5810_) );
NAND2X1 NAND2X1_748 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_6_bF_buf2_), .B(micro_hash_ucr_2_pipe50_bF_buf2), .Y(_5811_) );
NAND2X1 NAND2X1_749 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_6_bF_buf1_), .B(micro_hash_ucr_2_pipe48_bF_buf0), .Y(_5812_) );
NAND2X1 NAND2X1_750 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_6_bF_buf0_), .B(micro_hash_ucr_2_pipe46_bF_buf4), .Y(_5813_) );
NAND2X1 NAND2X1_751 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_6_bF_buf3_), .B(micro_hash_ucr_2_pipe44_bF_buf2), .Y(_5814_) );
NAND2X1 NAND2X1_752 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_6_bF_buf2_), .B(micro_hash_ucr_2_pipe32_bF_buf0), .Y(_5815_) );
NAND2X1 NAND2X1_753 ( .gnd(gnd), .vdd(vdd), .A(_8681_), .B(_4622__bF_buf2), .Y(_5816_) );
NAND2X1 NAND2X1_754 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_6_), .B(micro_hash_ucr_2_b_6_), .Y(_5817_) );
NAND2X1 NAND2X1_755 ( .gnd(gnd), .vdd(vdd), .A(_5817_), .B(_5816_), .Y(_5818_) );
INVX8 INVX8_180 ( .gnd(gnd), .vdd(vdd), .A(_5818__bF_buf3), .Y(_5819_) );
NAND2X1 NAND2X1_756 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe20_bF_buf1), .B(_4688_), .Y(_5820_) );
NOR2X1 NOR2X1_991 ( .gnd(gnd), .vdd(vdd), .A(_4688_), .B(_5122__bF_buf3), .Y(_5821_) );
NAND2X1 NAND2X1_757 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_6_bF_buf1_), .B(micro_hash_ucr_2_pipe14_bF_buf0), .Y(_5822_) );
NOR3X1 NOR3X1_6 ( .gnd(gnd), .vdd(vdd), .A(H_2_6_), .B(micro_hash_ucr_2_pipe12_bF_buf2), .C(micro_hash_ucr_2_pipe7), .Y(_5823_) );
NAND3X1 NAND3X1_249 ( .gnd(gnd), .vdd(vdd), .A(_5710_), .B(_5823_), .C(_5383_), .Y(_5824_) );
OAI21X1 OAI21X1_1635 ( .gnd(gnd), .vdd(vdd), .A(_5159_), .B(micro_hash_ucr_2_a_6_bF_buf0_), .C(_5824_), .Y(_5825_) );
AOI22X1 AOI22X1_48 ( .gnd(gnd), .vdd(vdd), .A(_4688_), .B(micro_hash_ucr_2_pipe12_bF_buf1), .C(_5825_), .D(_5132_), .Y(_5826_) );
AOI21X1 AOI21X1_1052 ( .gnd(gnd), .vdd(vdd), .A(_5818__bF_buf2), .B(_5392_), .C(micro_hash_ucr_2_pipe14_bF_buf4), .Y(_5827_) );
OAI21X1 OAI21X1_1636 ( .gnd(gnd), .vdd(vdd), .A(_5826_), .B(micro_hash_ucr_2_pipe13), .C(_5827_), .Y(_5828_) );
NAND3X1 NAND3X1_250 ( .gnd(gnd), .vdd(vdd), .A(_5125__bF_buf3), .B(_5822_), .C(_5828_), .Y(_5829_) );
NAND2X1 NAND2X1_758 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe15), .B(_5818__bF_buf1), .Y(_5830_) );
NAND3X1 NAND3X1_251 ( .gnd(gnd), .vdd(vdd), .A(_5127__bF_buf3), .B(_5830_), .C(_5829_), .Y(_5831_) );
AOI21X1 AOI21X1_1053 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_6_bF_buf3_), .B(micro_hash_ucr_2_pipe16_bF_buf2), .C(micro_hash_ucr_2_pipe17_bF_buf1), .Y(_5832_) );
OAI21X1 OAI21X1_1637 ( .gnd(gnd), .vdd(vdd), .A(_5819_), .B(_5126_), .C(_5122__bF_buf2), .Y(_5833_) );
AOI21X1 AOI21X1_1054 ( .gnd(gnd), .vdd(vdd), .A(_5832_), .B(_5831_), .C(_5833_), .Y(_5834_) );
OAI21X1 OAI21X1_1638 ( .gnd(gnd), .vdd(vdd), .A(_5834_), .B(_5821_), .C(_5124__bF_buf0), .Y(_5835_) );
NAND2X1 NAND2X1_759 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe19), .B(_5819_), .Y(_5836_) );
NAND3X1 NAND3X1_252 ( .gnd(gnd), .vdd(vdd), .A(_5123__bF_buf0), .B(_5836_), .C(_5835_), .Y(_5837_) );
NAND3X1 NAND3X1_253 ( .gnd(gnd), .vdd(vdd), .A(_5119_), .B(_5820_), .C(_5837_), .Y(_5838_) );
NAND2X1 NAND2X1_760 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe21_bF_buf2), .B(_5819_), .Y(_5839_) );
AOI21X1 AOI21X1_1055 ( .gnd(gnd), .vdd(vdd), .A(_5839_), .B(_5838_), .C(micro_hash_ucr_2_pipe22_bF_buf0), .Y(_5840_) );
OAI21X1 OAI21X1_1639 ( .gnd(gnd), .vdd(vdd), .A(_4688_), .B(_5121__bF_buf3), .C(_5120__bF_buf3), .Y(_5841_) );
OAI22X1 OAI22X1_85 ( .gnd(gnd), .vdd(vdd), .A(_5120__bF_buf2), .B(_5819_), .C(_5840_), .D(_5841_), .Y(_5842_) );
OAI21X1 OAI21X1_1640 ( .gnd(gnd), .vdd(vdd), .A(_5116__bF_buf2), .B(micro_hash_ucr_2_a_6_bF_buf2_), .C(_5118__bF_buf0), .Y(_5843_) );
AOI21X1 AOI21X1_1056 ( .gnd(gnd), .vdd(vdd), .A(_5116__bF_buf1), .B(_5842_), .C(_5843_), .Y(_5844_) );
OAI21X1 OAI21X1_1641 ( .gnd(gnd), .vdd(vdd), .A(_5818__bF_buf0), .B(_5118__bF_buf3), .C(_5117__bF_buf1), .Y(_5845_) );
OAI22X1 OAI22X1_86 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_6_bF_buf1_), .B(_5117__bF_buf0), .C(_5844_), .D(_5845_), .Y(_5846_) );
NAND2X1 NAND2X1_761 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe27), .B(_5819_), .Y(_5847_) );
OAI21X1 OAI21X1_1642 ( .gnd(gnd), .vdd(vdd), .A(_5846_), .B(micro_hash_ucr_2_pipe27), .C(_5847_), .Y(_5848_) );
AOI21X1 AOI21X1_1057 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe28_bF_buf3), .B(_4688_), .C(micro_hash_ucr_2_pipe29_bF_buf2), .Y(_5849_) );
OAI21X1 OAI21X1_1643 ( .gnd(gnd), .vdd(vdd), .A(_5848_), .B(micro_hash_ucr_2_pipe28_bF_buf2), .C(_5849_), .Y(_5850_) );
AOI21X1 AOI21X1_1058 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe29_bF_buf1), .B(_5819_), .C(micro_hash_ucr_2_pipe30_bF_buf2), .Y(_5851_) );
AOI22X1 AOI22X1_49 ( .gnd(gnd), .vdd(vdd), .A(_4688_), .B(micro_hash_ucr_2_pipe30_bF_buf1), .C(_5850_), .D(_5851_), .Y(_5852_) );
NAND2X1 NAND2X1_762 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe31), .B(_5818__bF_buf3), .Y(_5853_) );
OAI21X1 OAI21X1_1644 ( .gnd(gnd), .vdd(vdd), .A(_5852_), .B(micro_hash_ucr_2_pipe31), .C(_5853_), .Y(_5854_) );
OAI21X1 OAI21X1_1645 ( .gnd(gnd), .vdd(vdd), .A(_5854_), .B(micro_hash_ucr_2_pipe32_bF_buf3), .C(_5815_), .Y(_5855_) );
NAND2X1 NAND2X1_763 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe33_bF_buf0), .B(_5818__bF_buf2), .Y(_5856_) );
OAI21X1 OAI21X1_1646 ( .gnd(gnd), .vdd(vdd), .A(_5855_), .B(micro_hash_ucr_2_pipe33_bF_buf3), .C(_5856_), .Y(_5857_) );
OAI21X1 OAI21X1_1647 ( .gnd(gnd), .vdd(vdd), .A(_5109__bF_buf2), .B(micro_hash_ucr_2_a_6_bF_buf0_), .C(_5108__bF_buf0), .Y(_5858_) );
AOI21X1 AOI21X1_1059 ( .gnd(gnd), .vdd(vdd), .A(_5109__bF_buf1), .B(_5857_), .C(_5858_), .Y(_5859_) );
OAI21X1 OAI21X1_1648 ( .gnd(gnd), .vdd(vdd), .A(_5818__bF_buf1), .B(_5108__bF_buf3), .C(_5104__bF_buf2), .Y(_5860_) );
OAI22X1 OAI22X1_87 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_6_bF_buf3_), .B(_5104__bF_buf1), .C(_5859_), .D(_5860_), .Y(_5861_) );
OAI21X1 OAI21X1_1649 ( .gnd(gnd), .vdd(vdd), .A(_5819_), .B(_5106_), .C(_5105__bF_buf3), .Y(_5862_) );
AOI21X1 AOI21X1_1060 ( .gnd(gnd), .vdd(vdd), .A(_5106_), .B(_5861_), .C(_5862_), .Y(_5863_) );
NOR2X1 NOR2X1_992 ( .gnd(gnd), .vdd(vdd), .A(_4688_), .B(_5105__bF_buf2), .Y(_5864_) );
OAI21X1 OAI21X1_1650 ( .gnd(gnd), .vdd(vdd), .A(_5863_), .B(_5864_), .C(_5101_), .Y(_5865_) );
NAND2X1 NAND2X1_764 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe39), .B(_5819_), .Y(_5866_) );
AOI21X1 AOI21X1_1061 ( .gnd(gnd), .vdd(vdd), .A(_5866_), .B(_5865_), .C(micro_hash_ucr_2_pipe40_bF_buf1), .Y(_5867_) );
OAI21X1 OAI21X1_1651 ( .gnd(gnd), .vdd(vdd), .A(_4688_), .B(_5103__bF_buf1), .C(_5102_), .Y(_5868_) );
AOI21X1 AOI21X1_1062 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe41_bF_buf3), .B(_5818__bF_buf0), .C(micro_hash_ucr_2_pipe42_bF_buf0), .Y(_5869_) );
OAI21X1 OAI21X1_1652 ( .gnd(gnd), .vdd(vdd), .A(_5867_), .B(_5868_), .C(_5869_), .Y(_5870_) );
NAND2X1 NAND2X1_765 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_6_bF_buf2_), .B(micro_hash_ucr_2_pipe42_bF_buf3), .Y(_5871_) );
AOI21X1 AOI21X1_1063 ( .gnd(gnd), .vdd(vdd), .A(_5871_), .B(_5870_), .C(micro_hash_ucr_2_pipe43), .Y(_5872_) );
NOR2X1 NOR2X1_993 ( .gnd(gnd), .vdd(vdd), .A(_5100__bF_buf3), .B(_5818__bF_buf3), .Y(_5873_) );
OAI21X1 OAI21X1_1653 ( .gnd(gnd), .vdd(vdd), .A(_5872_), .B(_5873_), .C(_5099__bF_buf0), .Y(_5874_) );
AOI21X1 AOI21X1_1064 ( .gnd(gnd), .vdd(vdd), .A(_5814_), .B(_5874_), .C(micro_hash_ucr_2_pipe45_bF_buf3), .Y(_5875_) );
NOR2X1 NOR2X1_994 ( .gnd(gnd), .vdd(vdd), .A(_5095_), .B(_5818__bF_buf2), .Y(_5876_) );
OAI21X1 OAI21X1_1654 ( .gnd(gnd), .vdd(vdd), .A(_5875_), .B(_5876_), .C(_5097__bF_buf3), .Y(_5877_) );
AOI21X1 AOI21X1_1065 ( .gnd(gnd), .vdd(vdd), .A(_5813_), .B(_5877_), .C(micro_hash_ucr_2_pipe47), .Y(_5878_) );
NOR2X1 NOR2X1_995 ( .gnd(gnd), .vdd(vdd), .A(_5096__bF_buf2), .B(_5818__bF_buf1), .Y(_5879_) );
OAI21X1 OAI21X1_1655 ( .gnd(gnd), .vdd(vdd), .A(_5878_), .B(_5879_), .C(_5092__bF_buf4), .Y(_5880_) );
AOI21X1 AOI21X1_1066 ( .gnd(gnd), .vdd(vdd), .A(_5812_), .B(_5880_), .C(micro_hash_ucr_2_pipe49_bF_buf3), .Y(_5881_) );
NOR2X1 NOR2X1_996 ( .gnd(gnd), .vdd(vdd), .A(_5094_), .B(_5818__bF_buf0), .Y(_5882_) );
OAI21X1 OAI21X1_1656 ( .gnd(gnd), .vdd(vdd), .A(_5881_), .B(_5882_), .C(_5093__bF_buf4), .Y(_5883_) );
AOI21X1 AOI21X1_1067 ( .gnd(gnd), .vdd(vdd), .A(_5811_), .B(_5883_), .C(micro_hash_ucr_2_pipe51), .Y(_5884_) );
NOR2X1 NOR2X1_997 ( .gnd(gnd), .vdd(vdd), .A(_5089__bF_buf0), .B(_5818__bF_buf3), .Y(_5885_) );
OAI21X1 OAI21X1_1657 ( .gnd(gnd), .vdd(vdd), .A(_5884_), .B(_5885_), .C(_5091__bF_buf3), .Y(_5886_) );
OAI21X1 OAI21X1_1658 ( .gnd(gnd), .vdd(vdd), .A(_4688_), .B(_5091__bF_buf2), .C(_5886_), .Y(_5887_) );
OAI21X1 OAI21X1_1659 ( .gnd(gnd), .vdd(vdd), .A(_5818__bF_buf2), .B(_5090_), .C(_5086__bF_buf2), .Y(_5888_) );
AOI21X1 AOI21X1_1068 ( .gnd(gnd), .vdd(vdd), .A(_5090_), .B(_5887_), .C(_5888_), .Y(_5889_) );
OAI21X1 OAI21X1_1660 ( .gnd(gnd), .vdd(vdd), .A(_5086__bF_buf1), .B(micro_hash_ucr_2_a_6_bF_buf1_), .C(_5088_), .Y(_5890_) );
AOI21X1 AOI21X1_1069 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe55), .B(_5819_), .C(micro_hash_ucr_2_pipe56_bF_buf0), .Y(_5891_) );
OAI21X1 OAI21X1_1661 ( .gnd(gnd), .vdd(vdd), .A(_5889_), .B(_5890_), .C(_5891_), .Y(_5892_) );
NAND2X1 NAND2X1_766 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe56_bF_buf3), .B(_4688_), .Y(_5893_) );
NAND3X1 NAND3X1_254 ( .gnd(gnd), .vdd(vdd), .A(_5083_), .B(_5893_), .C(_5892_), .Y(_5894_) );
NAND2X1 NAND2X1_767 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe57_bF_buf3), .B(_5819_), .Y(_5895_) );
AOI21X1 AOI21X1_1070 ( .gnd(gnd), .vdd(vdd), .A(_5895_), .B(_5894_), .C(micro_hash_ucr_2_pipe58_bF_buf1), .Y(_5896_) );
OAI21X1 OAI21X1_1662 ( .gnd(gnd), .vdd(vdd), .A(_4688_), .B(_5085__bF_buf1), .C(_5084__bF_buf2), .Y(_5897_) );
AOI21X1 AOI21X1_1071 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe59), .B(_5818__bF_buf1), .C(micro_hash_ucr_2_pipe60_bF_buf2), .Y(_5898_) );
OAI21X1 OAI21X1_1663 ( .gnd(gnd), .vdd(vdd), .A(_5896_), .B(_5897_), .C(_5898_), .Y(_5899_) );
NAND2X1 NAND2X1_768 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_6_bF_buf0_), .B(micro_hash_ucr_2_pipe60_bF_buf1), .Y(_5900_) );
AOI21X1 AOI21X1_1072 ( .gnd(gnd), .vdd(vdd), .A(_5900_), .B(_5899_), .C(micro_hash_ucr_2_pipe61_bF_buf3), .Y(_5901_) );
NOR2X1 NOR2X1_998 ( .gnd(gnd), .vdd(vdd), .A(_5082_), .B(_5818__bF_buf0), .Y(_5902_) );
OAI21X1 OAI21X1_1664 ( .gnd(gnd), .vdd(vdd), .A(_5901_), .B(_5902_), .C(_5081__bF_buf1), .Y(_5903_) );
NAND3X1 NAND3X1_255 ( .gnd(gnd), .vdd(vdd), .A(_5077__bF_buf0), .B(_5810_), .C(_5903_), .Y(_5904_) );
NAND2X1 NAND2X1_769 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe63), .B(_5818__bF_buf3), .Y(_5905_) );
NAND3X1 NAND3X1_256 ( .gnd(gnd), .vdd(vdd), .A(_5079__bF_buf1), .B(_5905_), .C(_5904_), .Y(_5906_) );
NAND3X1 NAND3X1_257 ( .gnd(gnd), .vdd(vdd), .A(_5078_), .B(_5809_), .C(_5906_), .Y(_5907_) );
NAND2X1 NAND2X1_770 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe65_bF_buf1), .B(_5818__bF_buf2), .Y(_5908_) );
NAND3X1 NAND3X1_258 ( .gnd(gnd), .vdd(vdd), .A(_5074__bF_buf1), .B(_5908_), .C(_5907_), .Y(_5909_) );
NAND3X1 NAND3X1_259 ( .gnd(gnd), .vdd(vdd), .A(_5076__bF_buf3), .B(_5808_), .C(_5909_), .Y(_5910_) );
NAND2X1 NAND2X1_771 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe67), .B(_5818__bF_buf1), .Y(_5911_) );
NAND3X1 NAND3X1_260 ( .gnd(gnd), .vdd(vdd), .A(_5075__bF_buf2), .B(_5911_), .C(_5910_), .Y(_5912_) );
AOI21X1 AOI21X1_1073 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_6_bF_buf3_), .B(micro_hash_ucr_2_pipe68), .C(micro_hash_ucr_2_pipe69), .Y(_5913_) );
OAI21X1 OAI21X1_1665 ( .gnd(gnd), .vdd(vdd), .A(_5819_), .B(_5073__bF_buf1), .C(_4496__bF_buf13), .Y(_5914_) );
AOI21X1 AOI21X1_1074 ( .gnd(gnd), .vdd(vdd), .A(_5913_), .B(_5912_), .C(_5914_), .Y(_4491__6_) );
INVX8 INVX8_181 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_7_), .Y(_5915_) );
NAND2X1 NAND2X1_772 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe62_bF_buf0), .B(_5915__bF_buf3), .Y(_5916_) );
NAND2X1 NAND2X1_773 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe60_bF_buf0), .B(_5915__bF_buf2), .Y(_5917_) );
OR2X2 OR2X2_47 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_7_), .B(micro_hash_ucr_2_b_7_bF_buf2_), .Y(_5918_) );
NAND2X1 NAND2X1_774 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_7_), .B(micro_hash_ucr_2_b_7_bF_buf1_), .Y(_5919_) );
NAND2X1 NAND2X1_775 ( .gnd(gnd), .vdd(vdd), .A(_5919_), .B(_5918_), .Y(_5920_) );
INVX8 INVX8_182 ( .gnd(gnd), .vdd(vdd), .A(_5920_), .Y(_5921_) );
NAND2X1 NAND2X1_776 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe44_bF_buf1), .B(_5915__bF_buf1), .Y(_5922_) );
NAND2X1 NAND2X1_777 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe42_bF_buf2), .B(_5915__bF_buf0), .Y(_5923_) );
NAND2X1 NAND2X1_778 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe40_bF_buf0), .B(_5915__bF_buf3), .Y(_5924_) );
NAND2X1 NAND2X1_779 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe38_bF_buf3), .B(_5915__bF_buf2), .Y(_5925_) );
NAND2X1 NAND2X1_780 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe36_bF_buf0), .B(_5915__bF_buf1), .Y(_5926_) );
NAND2X1 NAND2X1_781 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe34_bF_buf0), .B(_5915__bF_buf0), .Y(_5927_) );
NAND2X1 NAND2X1_782 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe28_bF_buf1), .B(_5915__bF_buf3), .Y(_5928_) );
NOR2X1 NOR2X1_999 ( .gnd(gnd), .vdd(vdd), .A(_5126_), .B(_5920_), .Y(_5929_) );
NAND2X1 NAND2X1_783 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_7_), .B(micro_hash_ucr_2_pipe16_bF_buf1), .Y(_5930_) );
NOR2X1 NOR2X1_1000 ( .gnd(gnd), .vdd(vdd), .A(_5125__bF_buf2), .B(_5920_), .Y(_5931_) );
NAND2X1 NAND2X1_784 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_7_), .B(micro_hash_ucr_2_pipe14_bF_buf3), .Y(_5932_) );
NAND3X1 NAND3X1_261 ( .gnd(gnd), .vdd(vdd), .A(_4694_), .B(_5136_), .C(_5387_), .Y(_5933_) );
NOR2X1 NOR2X1_1001 ( .gnd(gnd), .vdd(vdd), .A(_5933_), .B(_5386_), .Y(_5934_) );
AOI21X1 AOI21X1_1075 ( .gnd(gnd), .vdd(vdd), .A(_5915__bF_buf2), .B(_5160_), .C(_5934_), .Y(_5935_) );
AOI21X1 AOI21X1_1076 ( .gnd(gnd), .vdd(vdd), .A(_5920_), .B(_5392_), .C(micro_hash_ucr_2_pipe14_bF_buf2), .Y(_5936_) );
OAI21X1 OAI21X1_1666 ( .gnd(gnd), .vdd(vdd), .A(_5935_), .B(micro_hash_ucr_2_pipe13), .C(_5936_), .Y(_5937_) );
AOI21X1 AOI21X1_1077 ( .gnd(gnd), .vdd(vdd), .A(_5932_), .B(_5937_), .C(micro_hash_ucr_2_pipe15), .Y(_5938_) );
OAI21X1 OAI21X1_1667 ( .gnd(gnd), .vdd(vdd), .A(_5938_), .B(_5931_), .C(_5127__bF_buf2), .Y(_5939_) );
AOI21X1 AOI21X1_1078 ( .gnd(gnd), .vdd(vdd), .A(_5930_), .B(_5939_), .C(micro_hash_ucr_2_pipe17_bF_buf0), .Y(_5940_) );
OAI21X1 OAI21X1_1668 ( .gnd(gnd), .vdd(vdd), .A(_5940_), .B(_5929_), .C(_5122__bF_buf1), .Y(_5941_) );
AOI21X1 AOI21X1_1079 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_7_), .B(micro_hash_ucr_2_pipe18_bF_buf0), .C(micro_hash_ucr_2_pipe19), .Y(_5942_) );
OAI21X1 OAI21X1_1669 ( .gnd(gnd), .vdd(vdd), .A(_5921__bF_buf3), .B(_5124__bF_buf3), .C(_5123__bF_buf4), .Y(_5943_) );
AOI21X1 AOI21X1_1080 ( .gnd(gnd), .vdd(vdd), .A(_5942_), .B(_5941_), .C(_5943_), .Y(_5944_) );
NOR2X1 NOR2X1_1002 ( .gnd(gnd), .vdd(vdd), .A(_5915__bF_buf1), .B(_5123__bF_buf3), .Y(_5945_) );
OAI21X1 OAI21X1_1670 ( .gnd(gnd), .vdd(vdd), .A(_5944_), .B(_5945_), .C(_5119_), .Y(_5946_) );
AOI21X1 AOI21X1_1081 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe21_bF_buf1), .B(_5921__bF_buf2), .C(micro_hash_ucr_2_pipe22_bF_buf4), .Y(_5947_) );
OAI21X1 OAI21X1_1671 ( .gnd(gnd), .vdd(vdd), .A(_5121__bF_buf2), .B(micro_hash_ucr_2_a_7_), .C(_5120__bF_buf1), .Y(_5948_) );
AOI21X1 AOI21X1_1082 ( .gnd(gnd), .vdd(vdd), .A(_5947_), .B(_5946_), .C(_5948_), .Y(_5949_) );
OAI21X1 OAI21X1_1672 ( .gnd(gnd), .vdd(vdd), .A(_5920_), .B(_5120__bF_buf0), .C(_5116__bF_buf0), .Y(_5950_) );
OAI22X1 OAI22X1_88 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_7_), .B(_5116__bF_buf4), .C(_5949_), .D(_5950_), .Y(_5951_) );
OAI21X1 OAI21X1_1673 ( .gnd(gnd), .vdd(vdd), .A(_5921__bF_buf1), .B(_5118__bF_buf2), .C(_5117__bF_buf4), .Y(_5952_) );
AOI21X1 AOI21X1_1083 ( .gnd(gnd), .vdd(vdd), .A(_5118__bF_buf1), .B(_5951_), .C(_5952_), .Y(_5953_) );
NOR2X1 NOR2X1_1003 ( .gnd(gnd), .vdd(vdd), .A(_5915__bF_buf0), .B(_5117__bF_buf3), .Y(_5954_) );
OAI21X1 OAI21X1_1674 ( .gnd(gnd), .vdd(vdd), .A(_5953_), .B(_5954_), .C(_5113_), .Y(_5955_) );
NAND2X1 NAND2X1_785 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe27), .B(_5921__bF_buf0), .Y(_5956_) );
NAND3X1 NAND3X1_262 ( .gnd(gnd), .vdd(vdd), .A(_5115__bF_buf4), .B(_5956_), .C(_5955_), .Y(_5957_) );
NAND3X1 NAND3X1_263 ( .gnd(gnd), .vdd(vdd), .A(_5114_), .B(_5928_), .C(_5957_), .Y(_5958_) );
AOI21X1 AOI21X1_1084 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe29_bF_buf0), .B(_5921__bF_buf3), .C(micro_hash_ucr_2_pipe30_bF_buf0), .Y(_5959_) );
AND2X2 AND2X2_430 ( .gnd(gnd), .vdd(vdd), .A(_5958_), .B(_5959_), .Y(_5960_) );
OAI21X1 OAI21X1_1675 ( .gnd(gnd), .vdd(vdd), .A(_5110__bF_buf0), .B(micro_hash_ucr_2_a_7_), .C(_5112__bF_buf2), .Y(_5961_) );
AOI21X1 AOI21X1_1085 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe31), .B(_5921__bF_buf2), .C(micro_hash_ucr_2_pipe32_bF_buf2), .Y(_5962_) );
OAI21X1 OAI21X1_1676 ( .gnd(gnd), .vdd(vdd), .A(_5960_), .B(_5961_), .C(_5962_), .Y(_5963_) );
NAND2X1 NAND2X1_786 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe32_bF_buf1), .B(_5915__bF_buf3), .Y(_5964_) );
NAND3X1 NAND3X1_264 ( .gnd(gnd), .vdd(vdd), .A(_5107_), .B(_5964_), .C(_5963_), .Y(_5965_) );
NAND2X1 NAND2X1_787 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe33_bF_buf2), .B(_5921__bF_buf1), .Y(_5966_) );
NAND3X1 NAND3X1_265 ( .gnd(gnd), .vdd(vdd), .A(_5109__bF_buf0), .B(_5966_), .C(_5965_), .Y(_5967_) );
NAND3X1 NAND3X1_266 ( .gnd(gnd), .vdd(vdd), .A(_5108__bF_buf2), .B(_5927_), .C(_5967_), .Y(_5968_) );
NAND2X1 NAND2X1_788 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe35), .B(_5921__bF_buf0), .Y(_5969_) );
NAND3X1 NAND3X1_267 ( .gnd(gnd), .vdd(vdd), .A(_5104__bF_buf0), .B(_5969_), .C(_5968_), .Y(_5970_) );
NAND3X1 NAND3X1_268 ( .gnd(gnd), .vdd(vdd), .A(_5106_), .B(_5926_), .C(_5970_), .Y(_5971_) );
NAND2X1 NAND2X1_789 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe37), .B(_5921__bF_buf3), .Y(_5972_) );
NAND3X1 NAND3X1_269 ( .gnd(gnd), .vdd(vdd), .A(_5105__bF_buf1), .B(_5972_), .C(_5971_), .Y(_5973_) );
NAND3X1 NAND3X1_270 ( .gnd(gnd), .vdd(vdd), .A(_5101_), .B(_5925_), .C(_5973_), .Y(_5974_) );
NAND2X1 NAND2X1_790 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe39), .B(_5921__bF_buf2), .Y(_5975_) );
NAND3X1 NAND3X1_271 ( .gnd(gnd), .vdd(vdd), .A(_5103__bF_buf0), .B(_5975_), .C(_5974_), .Y(_5976_) );
NAND3X1 NAND3X1_272 ( .gnd(gnd), .vdd(vdd), .A(_5102_), .B(_5924_), .C(_5976_), .Y(_5977_) );
NAND2X1 NAND2X1_791 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe41_bF_buf2), .B(_5921__bF_buf1), .Y(_5978_) );
NAND3X1 NAND3X1_273 ( .gnd(gnd), .vdd(vdd), .A(_5098__bF_buf2), .B(_5978_), .C(_5977_), .Y(_5979_) );
NAND3X1 NAND3X1_274 ( .gnd(gnd), .vdd(vdd), .A(_5100__bF_buf2), .B(_5923_), .C(_5979_), .Y(_5980_) );
NAND2X1 NAND2X1_792 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe43), .B(_5921__bF_buf0), .Y(_5981_) );
NAND3X1 NAND3X1_275 ( .gnd(gnd), .vdd(vdd), .A(_5099__bF_buf4), .B(_5981_), .C(_5980_), .Y(_5982_) );
NAND3X1 NAND3X1_276 ( .gnd(gnd), .vdd(vdd), .A(_5095_), .B(_5922_), .C(_5982_), .Y(_5983_) );
AOI21X1 AOI21X1_1086 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe45_bF_buf2), .B(_5921__bF_buf3), .C(micro_hash_ucr_2_pipe46_bF_buf3), .Y(_5984_) );
OAI21X1 OAI21X1_1677 ( .gnd(gnd), .vdd(vdd), .A(_5097__bF_buf2), .B(micro_hash_ucr_2_a_7_), .C(_5096__bF_buf1), .Y(_5985_) );
AOI21X1 AOI21X1_1087 ( .gnd(gnd), .vdd(vdd), .A(_5984_), .B(_5983_), .C(_5985_), .Y(_5986_) );
OAI21X1 OAI21X1_1678 ( .gnd(gnd), .vdd(vdd), .A(_5920_), .B(_5096__bF_buf0), .C(_5092__bF_buf3), .Y(_5987_) );
OAI22X1 OAI22X1_89 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_7_), .B(_5092__bF_buf2), .C(_5986_), .D(_5987_), .Y(_5988_) );
NAND2X1 NAND2X1_793 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe49_bF_buf2), .B(_5921__bF_buf2), .Y(_5989_) );
OAI21X1 OAI21X1_1679 ( .gnd(gnd), .vdd(vdd), .A(_5988_), .B(micro_hash_ucr_2_pipe49_bF_buf1), .C(_5989_), .Y(_5990_) );
NAND2X1 NAND2X1_794 ( .gnd(gnd), .vdd(vdd), .A(_5093__bF_buf3), .B(_5990_), .Y(_5991_) );
OAI21X1 OAI21X1_1680 ( .gnd(gnd), .vdd(vdd), .A(_5915__bF_buf2), .B(_5093__bF_buf2), .C(_5991_), .Y(_5992_) );
NAND2X1 NAND2X1_795 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe51), .B(_5920_), .Y(_5993_) );
OAI21X1 OAI21X1_1681 ( .gnd(gnd), .vdd(vdd), .A(_5992_), .B(micro_hash_ucr_2_pipe51), .C(_5993_), .Y(_5994_) );
OAI21X1 OAI21X1_1682 ( .gnd(gnd), .vdd(vdd), .A(_5091__bF_buf1), .B(micro_hash_ucr_2_a_7_), .C(_5090_), .Y(_5995_) );
AOI21X1 AOI21X1_1088 ( .gnd(gnd), .vdd(vdd), .A(_5091__bF_buf0), .B(_5994_), .C(_5995_), .Y(_5996_) );
AOI21X1 AOI21X1_1089 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe53_bF_buf2), .B(_5921__bF_buf1), .C(_5996_), .Y(_5997_) );
AOI21X1 AOI21X1_1090 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_7_), .B(micro_hash_ucr_2_pipe54_bF_buf0), .C(micro_hash_ucr_2_pipe55), .Y(_5998_) );
OAI21X1 OAI21X1_1683 ( .gnd(gnd), .vdd(vdd), .A(_5997_), .B(micro_hash_ucr_2_pipe54_bF_buf4), .C(_5998_), .Y(_5999_) );
NAND2X1 NAND2X1_796 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe55), .B(_5920_), .Y(_6000_) );
AOI21X1 AOI21X1_1091 ( .gnd(gnd), .vdd(vdd), .A(_6000_), .B(_5999_), .C(micro_hash_ucr_2_pipe56_bF_buf2), .Y(_6001_) );
OAI21X1 OAI21X1_1684 ( .gnd(gnd), .vdd(vdd), .A(_5087__bF_buf2), .B(micro_hash_ucr_2_a_7_), .C(_5083_), .Y(_6002_) );
AOI21X1 AOI21X1_1092 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe57_bF_buf2), .B(_5921__bF_buf0), .C(micro_hash_ucr_2_pipe58_bF_buf0), .Y(_6003_) );
OAI21X1 OAI21X1_1685 ( .gnd(gnd), .vdd(vdd), .A(_6001_), .B(_6002_), .C(_6003_), .Y(_6004_) );
NAND2X1 NAND2X1_797 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe58_bF_buf4), .B(_5915__bF_buf1), .Y(_6005_) );
AOI21X1 AOI21X1_1093 ( .gnd(gnd), .vdd(vdd), .A(_6005_), .B(_6004_), .C(micro_hash_ucr_2_pipe59), .Y(_6006_) );
NOR2X1 NOR2X1_1004 ( .gnd(gnd), .vdd(vdd), .A(_5084__bF_buf1), .B(_5921__bF_buf3), .Y(_6007_) );
OAI21X1 OAI21X1_1686 ( .gnd(gnd), .vdd(vdd), .A(_6006_), .B(_6007_), .C(_5080__bF_buf0), .Y(_6008_) );
AOI21X1 AOI21X1_1094 ( .gnd(gnd), .vdd(vdd), .A(_5917_), .B(_6008_), .C(micro_hash_ucr_2_pipe61_bF_buf2), .Y(_6009_) );
NOR2X1 NOR2X1_1005 ( .gnd(gnd), .vdd(vdd), .A(_5082_), .B(_5921__bF_buf2), .Y(_6010_) );
OAI21X1 OAI21X1_1687 ( .gnd(gnd), .vdd(vdd), .A(_6009_), .B(_6010_), .C(_5081__bF_buf0), .Y(_6011_) );
NAND3X1 NAND3X1_277 ( .gnd(gnd), .vdd(vdd), .A(_5077__bF_buf3), .B(_5916_), .C(_6011_), .Y(_6012_) );
NAND2X1 NAND2X1_798 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe63), .B(_5921__bF_buf1), .Y(_6013_) );
AOI21X1 AOI21X1_1095 ( .gnd(gnd), .vdd(vdd), .A(_6013_), .B(_6012_), .C(micro_hash_ucr_2_pipe64_bF_buf2), .Y(_6014_) );
OAI21X1 OAI21X1_1688 ( .gnd(gnd), .vdd(vdd), .A(_5915__bF_buf0), .B(_5079__bF_buf0), .C(_5078_), .Y(_6015_) );
AOI21X1 AOI21X1_1096 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe65_bF_buf0), .B(_5920_), .C(micro_hash_ucr_2_pipe66_bF_buf0), .Y(_6016_) );
OAI21X1 OAI21X1_1689 ( .gnd(gnd), .vdd(vdd), .A(_6014_), .B(_6015_), .C(_6016_), .Y(_6017_) );
NAND2X1 NAND2X1_799 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_7_), .B(micro_hash_ucr_2_pipe66_bF_buf4), .Y(_6018_) );
NAND3X1 NAND3X1_278 ( .gnd(gnd), .vdd(vdd), .A(_5076__bF_buf2), .B(_6018_), .C(_6017_), .Y(_6019_) );
NAND2X1 NAND2X1_800 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe67), .B(_5920_), .Y(_6020_) );
NAND3X1 NAND3X1_279 ( .gnd(gnd), .vdd(vdd), .A(_5075__bF_buf1), .B(_6020_), .C(_6019_), .Y(_6021_) );
AOI21X1 AOI21X1_1097 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_a_7_), .B(micro_hash_ucr_2_pipe68), .C(micro_hash_ucr_2_pipe69), .Y(_6022_) );
OAI21X1 OAI21X1_1690 ( .gnd(gnd), .vdd(vdd), .A(_5921__bF_buf0), .B(_5073__bF_buf0), .C(_4496__bF_buf12), .Y(_6023_) );
AOI21X1 AOI21X1_1098 ( .gnd(gnd), .vdd(vdd), .A(_6022_), .B(_6021_), .C(_6023_), .Y(_4491__7_) );
INVX1 INVX1_370 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_k_0_), .Y(_6024_) );
NOR2X1 NOR2X1_1006 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe40_bF_buf4), .B(micro_hash_ucr_2_pipe7), .Y(_6025_) );
AOI21X1 AOI21X1_1099 ( .gnd(gnd), .vdd(vdd), .A(_6024_), .B(_6025_), .C(_4594__bF_buf0), .Y(_4495__0_) );
NAND2X1 NAND2X1_801 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_k_1_), .B(_6025_), .Y(_6026_) );
NOR2X1 NOR2X1_1007 ( .gnd(gnd), .vdd(vdd), .A(_6026_), .B(_4594__bF_buf12), .Y(_4495__1_) );
NAND2X1 NAND2X1_802 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_k_2_), .B(_6025_), .Y(_6027_) );
NOR2X1 NOR2X1_1008 ( .gnd(gnd), .vdd(vdd), .A(_6027_), .B(_4594__bF_buf11), .Y(_4495__2_) );
OAI21X1 OAI21X1_1691 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe7), .B(micro_hash_ucr_2_k_3_), .C(_5103__bF_buf3), .Y(_6028_) );
NOR2X1 NOR2X1_1009 ( .gnd(gnd), .vdd(vdd), .A(_6028_), .B(_4594__bF_buf10), .Y(_4495__3_) );
OAI21X1 OAI21X1_1692 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe7), .B(micro_hash_ucr_2_k_4_), .C(_5103__bF_buf2), .Y(_6029_) );
NOR2X1 NOR2X1_1010 ( .gnd(gnd), .vdd(vdd), .A(_6029_), .B(_4594__bF_buf9), .Y(_4495__4_) );
INVX2 INVX2_217 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_k_5_), .Y(_6030_) );
OAI21X1 OAI21X1_1693 ( .gnd(gnd), .vdd(vdd), .A(_6030_), .B(micro_hash_ucr_2_pipe7), .C(_5103__bF_buf1), .Y(_6031_) );
AND2X2 AND2X2_431 ( .gnd(gnd), .vdd(vdd), .A(_4496__bF_buf11), .B(_6031_), .Y(_4495__5_) );
NAND2X1 NAND2X1_803 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_k_6_), .B(_6025_), .Y(_6032_) );
NOR2X1 NOR2X1_1011 ( .gnd(gnd), .vdd(vdd), .A(_6032_), .B(_4594__bF_buf8), .Y(_4495__6_) );
INVX1 INVX1_371 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_k_7_), .Y(_6033_) );
AOI21X1 AOI21X1_1100 ( .gnd(gnd), .vdd(vdd), .A(_6033_), .B(_6025_), .C(_4594__bF_buf7), .Y(_4495__7_) );
NAND2X1 NAND2X1_804 ( .gnd(gnd), .vdd(vdd), .A(_8690_), .B(_4630_), .Y(_6034_) );
NOR2X1 NOR2X1_1012 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe21_bF_buf0), .B(micro_hash_ucr_2_pipe23), .Y(_6035_) );
INVX1 INVX1_372 ( .gnd(gnd), .vdd(vdd), .A(_6035_), .Y(_6036_) );
NOR2X1 NOR2X1_1013 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe39), .B(micro_hash_ucr_2_pipe37), .Y(_6037_) );
INVX1 INVX1_373 ( .gnd(gnd), .vdd(vdd), .A(_6037_), .Y(_6038_) );
NOR2X1 NOR2X1_1014 ( .gnd(gnd), .vdd(vdd), .A(_6036_), .B(_6038_), .Y(_6039_) );
NOR2X1 NOR2X1_1015 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe27), .B(micro_hash_ucr_2_pipe29_bF_buf3), .Y(_6040_) );
AND2X2 AND2X2_432 ( .gnd(gnd), .vdd(vdd), .A(_6040_), .B(_5108__bF_buf1), .Y(_6041_) );
AND2X2 AND2X2_433 ( .gnd(gnd), .vdd(vdd), .A(_6039_), .B(_6041_), .Y(_6042_) );
NAND3X1 NAND3X1_280 ( .gnd(gnd), .vdd(vdd), .A(_5107_), .B(_5112__bF_buf1), .C(_5174_), .Y(_6043_) );
NOR2X1 NOR2X1_1016 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe25), .B(micro_hash_ucr_2_pipe19), .Y(_6044_) );
NAND2X1 NAND2X1_805 ( .gnd(gnd), .vdd(vdd), .A(_5168_), .B(_5494_), .Y(_6045_) );
INVX1 INVX1_374 ( .gnd(gnd), .vdd(vdd), .A(_6045_), .Y(_6046_) );
NAND2X1 NAND2X1_806 ( .gnd(gnd), .vdd(vdd), .A(_6044_), .B(_6046_), .Y(_6047_) );
NOR2X1 NOR2X1_1017 ( .gnd(gnd), .vdd(vdd), .A(_6043_), .B(_6047_), .Y(_6048_) );
NAND2X1 NAND2X1_807 ( .gnd(gnd), .vdd(vdd), .A(_6042_), .B(_6048_), .Y(_6049_) );
INVX4 INVX4_106 ( .gnd(gnd), .vdd(vdd), .A(_6049_), .Y(_6050_) );
AOI21X1 AOI21X1_1101 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_0_bF_buf0_), .B(micro_hash_ucr_2_a_0_), .C(_6050_), .Y(_6051_) );
NOR2X1 NOR2X1_1018 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe45_bF_buf1), .B(micro_hash_ucr_2_pipe47), .Y(_6052_) );
NAND3X1 NAND3X1_281 ( .gnd(gnd), .vdd(vdd), .A(_5100__bF_buf1), .B(_5102_), .C(_6052_), .Y(_6053_) );
NOR2X1 NOR2X1_1019 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe55), .B(micro_hash_ucr_2_pipe51), .Y(_6054_) );
NAND3X1 NAND3X1_282 ( .gnd(gnd), .vdd(vdd), .A(_5090_), .B(_5094_), .C(_6054_), .Y(_6055_) );
NOR2X1 NOR2X1_1020 ( .gnd(gnd), .vdd(vdd), .A(_6053_), .B(_6055_), .Y(_6056_) );
NOR2X1 NOR2X1_1021 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe67), .B(micro_hash_ucr_2_pipe65_bF_buf3), .Y(_6057_) );
INVX2 INVX2_218 ( .gnd(gnd), .vdd(vdd), .A(_6057_), .Y(_6058_) );
NOR2X1 NOR2X1_1022 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe63), .B(micro_hash_ucr_2_pipe61_bF_buf1), .Y(_6059_) );
NAND3X1 NAND3X1_283 ( .gnd(gnd), .vdd(vdd), .A(_5083_), .B(_5084__bF_buf0), .C(_6059_), .Y(_6060_) );
NOR2X1 NOR2X1_1023 ( .gnd(gnd), .vdd(vdd), .A(_6058_), .B(_6060_), .Y(_6061_) );
NAND2X1 NAND2X1_808 ( .gnd(gnd), .vdd(vdd), .A(_6061_), .B(_6056_), .Y(_6062_) );
OAI21X1 OAI21X1_1694 ( .gnd(gnd), .vdd(vdd), .A(_6051_), .B(_6062_), .C(_6034_), .Y(_6063_) );
INVX2 INVX2_219 ( .gnd(gnd), .vdd(vdd), .A(_6056_), .Y(_6064_) );
NOR2X1 NOR2X1_1024 ( .gnd(gnd), .vdd(vdd), .A(_6060_), .B(_6064_), .Y(_6065_) );
NOR2X1 NOR2X1_1025 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe19), .B(_6036_), .Y(_6066_) );
NAND3X1 NAND3X1_284 ( .gnd(gnd), .vdd(vdd), .A(_5107_), .B(micro_hash_ucr_2_x_0_), .C(_5168_), .Y(_6067_) );
NOR2X1 NOR2X1_1026 ( .gnd(gnd), .vdd(vdd), .A(_6058_), .B(_6067_), .Y(_6068_) );
NAND2X1 NAND2X1_809 ( .gnd(gnd), .vdd(vdd), .A(_6066_), .B(_6068_), .Y(_6069_) );
NOR2X1 NOR2X1_1027 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe31), .B(micro_hash_ucr_2_pipe29_bF_buf2), .Y(_6070_) );
NAND3X1 NAND3X1_285 ( .gnd(gnd), .vdd(vdd), .A(_5174_), .B(_5494_), .C(_6070_), .Y(_6071_) );
NOR2X1 NOR2X1_1028 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe27), .B(micro_hash_ucr_2_pipe25), .Y(_6072_) );
NAND3X1 NAND3X1_286 ( .gnd(gnd), .vdd(vdd), .A(_5108__bF_buf0), .B(_6037_), .C(_6072_), .Y(_6073_) );
OR2X2 OR2X2_48 ( .gnd(gnd), .vdd(vdd), .A(_6071_), .B(_6073_), .Y(_6074_) );
NOR2X1 NOR2X1_1029 ( .gnd(gnd), .vdd(vdd), .A(_6074_), .B(_6069_), .Y(_6075_) );
AOI21X1 AOI21X1_1102 ( .gnd(gnd), .vdd(vdd), .A(_6065_), .B(_6075_), .C(micro_hash_ucr_2_pipe69), .Y(_6076_) );
OAI21X1 OAI21X1_1695 ( .gnd(gnd), .vdd(vdd), .A(_5073__bF_buf3), .B(_6034_), .C(_4496__bF_buf10), .Y(_6077_) );
AOI21X1 AOI21X1_1103 ( .gnd(gnd), .vdd(vdd), .A(_6076_), .B(_6063_), .C(_6077_), .Y(_4569__0_) );
NAND2X1 NAND2X1_810 ( .gnd(gnd), .vdd(vdd), .A(_8696_), .B(_4636_), .Y(_6078_) );
AOI21X1 AOI21X1_1104 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_1_bF_buf0_), .B(micro_hash_ucr_2_a_1_bF_buf2_), .C(_6050_), .Y(_6079_) );
OAI21X1 OAI21X1_1696 ( .gnd(gnd), .vdd(vdd), .A(_6079_), .B(_6062_), .C(_6078_), .Y(_6080_) );
INVX1 INVX1_375 ( .gnd(gnd), .vdd(vdd), .A(_6065_), .Y(_6081_) );
NAND2X1 NAND2X1_811 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_x_1_), .B(_6057_), .Y(_6082_) );
NOR2X1 NOR2X1_1030 ( .gnd(gnd), .vdd(vdd), .A(_6082_), .B(_6081_), .Y(_6083_) );
AOI21X1 AOI21X1_1105 ( .gnd(gnd), .vdd(vdd), .A(_6050_), .B(_6083_), .C(micro_hash_ucr_2_pipe69), .Y(_6084_) );
OAI21X1 OAI21X1_1697 ( .gnd(gnd), .vdd(vdd), .A(_5073__bF_buf2), .B(_6078_), .C(_4496__bF_buf9), .Y(_6085_) );
AOI21X1 AOI21X1_1106 ( .gnd(gnd), .vdd(vdd), .A(_6084_), .B(_6080_), .C(_6085_), .Y(_4569__1_) );
AOI21X1 AOI21X1_1107 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_2_bF_buf0_), .B(micro_hash_ucr_2_a_2_), .C(_6050_), .Y(_6086_) );
NOR2X1 NOR2X1_1031 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe69), .B(_6058_), .Y(_6087_) );
NAND2X1 NAND2X1_812 ( .gnd(gnd), .vdd(vdd), .A(_6087_), .B(_6065_), .Y(_6088_) );
OAI22X1 OAI22X1_90 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_2_bF_buf3_), .B(micro_hash_ucr_2_a_2_), .C(_6086_), .D(_6088_), .Y(_6089_) );
NAND3X1 NAND3X1_287 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_x_2_), .B(_6035_), .C(_6040_), .Y(_6090_) );
NOR2X1 NOR2X1_1032 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe35), .B(_6038_), .Y(_6091_) );
NAND2X1 NAND2X1_813 ( .gnd(gnd), .vdd(vdd), .A(_6091_), .B(_6087_), .Y(_6092_) );
NOR2X1 NOR2X1_1033 ( .gnd(gnd), .vdd(vdd), .A(_6090_), .B(_6092_), .Y(_6093_) );
NAND3X1 NAND3X1_288 ( .gnd(gnd), .vdd(vdd), .A(_6048_), .B(_6093_), .C(_6065_), .Y(_6094_) );
AOI21X1 AOI21X1_1108 ( .gnd(gnd), .vdd(vdd), .A(_6094_), .B(_6089_), .C(_4594__bF_buf6), .Y(_4569__2_) );
AOI21X1 AOI21X1_1109 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_3_bF_buf0_), .B(micro_hash_ucr_2_a_3_), .C(_6050_), .Y(_6095_) );
OAI22X1 OAI22X1_91 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_3_bF_buf3_), .B(micro_hash_ucr_2_a_3_), .C(_6095_), .D(_6088_), .Y(_6096_) );
NOR2X1 NOR2X1_1034 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe33_bF_buf1), .B(_6073_), .Y(_6097_) );
NAND2X1 NAND2X1_814 ( .gnd(gnd), .vdd(vdd), .A(_5125__bF_buf1), .B(_5494_), .Y(_6098_) );
NAND3X1 NAND3X1_289 ( .gnd(gnd), .vdd(vdd), .A(_5073__bF_buf1), .B(micro_hash_ucr_2_x_3_), .C(_6070_), .Y(_6099_) );
NOR2X1 NOR2X1_1035 ( .gnd(gnd), .vdd(vdd), .A(_6098_), .B(_6099_), .Y(_6100_) );
AND2X2 AND2X2_434 ( .gnd(gnd), .vdd(vdd), .A(_6056_), .B(_6100_), .Y(_6101_) );
NOR2X1 NOR2X1_1036 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe19), .B(micro_hash_ucr_2_pipe17_bF_buf3), .Y(_6102_) );
NAND3X1 NAND3X1_290 ( .gnd(gnd), .vdd(vdd), .A(_5168_), .B(_6035_), .C(_6102_), .Y(_6103_) );
INVX2 INVX2_220 ( .gnd(gnd), .vdd(vdd), .A(_6061_), .Y(_6104_) );
NOR2X1 NOR2X1_1037 ( .gnd(gnd), .vdd(vdd), .A(_6103_), .B(_6104_), .Y(_6105_) );
NAND3X1 NAND3X1_291 ( .gnd(gnd), .vdd(vdd), .A(_6097_), .B(_6105_), .C(_6101_), .Y(_6106_) );
AOI21X1 AOI21X1_1110 ( .gnd(gnd), .vdd(vdd), .A(_6106_), .B(_6096_), .C(_4594__bF_buf5), .Y(_4569__3_) );
NOR2X1 NOR2X1_1038 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_4_bF_buf3_), .B(micro_hash_ucr_2_a_4_), .Y(_6107_) );
OAI21X1 OAI21X1_1698 ( .gnd(gnd), .vdd(vdd), .A(_6058_), .B(_6107_), .C(_6104_), .Y(_6108_) );
NAND2X1 NAND2X1_815 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_x_4_), .B(_6050_), .Y(_6109_) );
NOR2X1 NOR2X1_1039 ( .gnd(gnd), .vdd(vdd), .A(_5593_), .B(_4668__bF_buf1), .Y(_6110_) );
NOR2X1 NOR2X1_1040 ( .gnd(gnd), .vdd(vdd), .A(_6107_), .B(_6110_), .Y(_6111_) );
AOI21X1 AOI21X1_1111 ( .gnd(gnd), .vdd(vdd), .A(_6111_), .B(_6049_), .C(_6064_), .Y(_6112_) );
AOI22X1 AOI22X1_50 ( .gnd(gnd), .vdd(vdd), .A(_6064_), .B(_6107_), .C(_6109_), .D(_6112_), .Y(_6113_) );
OAI21X1 OAI21X1_1699 ( .gnd(gnd), .vdd(vdd), .A(_6113_), .B(_6060_), .C(_6108_), .Y(_6114_) );
INVX1 INVX1_376 ( .gnd(gnd), .vdd(vdd), .A(_6107_), .Y(_6115_) );
AOI21X1 AOI21X1_1112 ( .gnd(gnd), .vdd(vdd), .A(_6058_), .B(_6115_), .C(micro_hash_ucr_2_pipe69), .Y(_6116_) );
OAI21X1 OAI21X1_1700 ( .gnd(gnd), .vdd(vdd), .A(_5073__bF_buf0), .B(_6115_), .C(_4496__bF_buf8), .Y(_6117_) );
AOI21X1 AOI21X1_1113 ( .gnd(gnd), .vdd(vdd), .A(_6116_), .B(_6114_), .C(_6117_), .Y(_4569__4_) );
AOI21X1 AOI21X1_1114 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_5_bF_buf3_), .B(micro_hash_ucr_2_a_5_bF_buf0_), .C(_6050_), .Y(_6118_) );
OAI22X1 OAI22X1_92 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_5_bF_buf2_), .B(micro_hash_ucr_2_a_5_bF_buf3_), .C(_6118_), .D(_6088_), .Y(_6119_) );
NAND3X1 NAND3X1_292 ( .gnd(gnd), .vdd(vdd), .A(_5107_), .B(_5108__bF_buf3), .C(_5112__bF_buf0), .Y(_6120_) );
NAND2X1 NAND2X1_816 ( .gnd(gnd), .vdd(vdd), .A(_6046_), .B(_6087_), .Y(_6121_) );
NOR2X1 NOR2X1_1041 ( .gnd(gnd), .vdd(vdd), .A(_6120_), .B(_6121_), .Y(_6122_) );
NAND2X1 NAND2X1_817 ( .gnd(gnd), .vdd(vdd), .A(_6044_), .B(_6039_), .Y(_6123_) );
NAND3X1 NAND3X1_293 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_x_5_), .B(_5174_), .C(_6040_), .Y(_6124_) );
NOR2X1 NOR2X1_1042 ( .gnd(gnd), .vdd(vdd), .A(_6124_), .B(_6123_), .Y(_6125_) );
NAND3X1 NAND3X1_294 ( .gnd(gnd), .vdd(vdd), .A(_6122_), .B(_6125_), .C(_6065_), .Y(_6126_) );
AOI21X1 AOI21X1_1115 ( .gnd(gnd), .vdd(vdd), .A(_6126_), .B(_6119_), .C(_4594__bF_buf4), .Y(_4569__5_) );
AOI21X1 AOI21X1_1116 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_6_), .B(micro_hash_ucr_2_a_6_bF_buf2_), .C(_6050_), .Y(_6127_) );
OAI22X1 OAI22X1_93 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_6_), .B(micro_hash_ucr_2_a_6_bF_buf1_), .C(_6127_), .D(_6088_), .Y(_6128_) );
NAND3X1 NAND3X1_295 ( .gnd(gnd), .vdd(vdd), .A(_5073__bF_buf3), .B(micro_hash_ucr_2_x_6_), .C(_6040_), .Y(_6129_) );
NOR2X1 NOR2X1_1043 ( .gnd(gnd), .vdd(vdd), .A(_6120_), .B(_6129_), .Y(_6130_) );
NAND2X1 NAND2X1_818 ( .gnd(gnd), .vdd(vdd), .A(_5174_), .B(_6046_), .Y(_6131_) );
OR2X2 OR2X2_49 ( .gnd(gnd), .vdd(vdd), .A(_6104_), .B(_6123_), .Y(_6132_) );
NOR2X1 NOR2X1_1044 ( .gnd(gnd), .vdd(vdd), .A(_6131_), .B(_6132_), .Y(_6133_) );
NAND3X1 NAND3X1_296 ( .gnd(gnd), .vdd(vdd), .A(_6056_), .B(_6130_), .C(_6133_), .Y(_6134_) );
AOI21X1 AOI21X1_1117 ( .gnd(gnd), .vdd(vdd), .A(_6134_), .B(_6128_), .C(_4594__bF_buf3), .Y(_4569__6_) );
INVX8 INVX8_183 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_7_bF_buf0_), .Y(_6135_) );
NAND2X1 NAND2X1_819 ( .gnd(gnd), .vdd(vdd), .A(_6135__bF_buf3), .B(_5915__bF_buf3), .Y(_6136_) );
AOI21X1 AOI21X1_1118 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_7_bF_buf3_), .B(micro_hash_ucr_2_a_7_), .C(_6050_), .Y(_6137_) );
OAI21X1 OAI21X1_1701 ( .gnd(gnd), .vdd(vdd), .A(_6137_), .B(_6062_), .C(_6136_), .Y(_6138_) );
AND2X2 AND2X2_435 ( .gnd(gnd), .vdd(vdd), .A(_6070_), .B(_5107_), .Y(_6139_) );
NAND3X1 NAND3X1_297 ( .gnd(gnd), .vdd(vdd), .A(_6072_), .B(_6139_), .C(_6091_), .Y(_6140_) );
NOR2X1 NOR2X1_1045 ( .gnd(gnd), .vdd(vdd), .A(_6131_), .B(_6140_), .Y(_6141_) );
NAND3X1 NAND3X1_298 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_x_7_), .B(_6057_), .C(_6066_), .Y(_6142_) );
NOR2X1 NOR2X1_1046 ( .gnd(gnd), .vdd(vdd), .A(_6142_), .B(_6081_), .Y(_6143_) );
AOI21X1 AOI21X1_1119 ( .gnd(gnd), .vdd(vdd), .A(_6141_), .B(_6143_), .C(micro_hash_ucr_2_pipe69), .Y(_6144_) );
OAI21X1 OAI21X1_1702 ( .gnd(gnd), .vdd(vdd), .A(_5073__bF_buf2), .B(_6136_), .C(_4496__bF_buf7), .Y(_6145_) );
AOI21X1 AOI21X1_1120 ( .gnd(gnd), .vdd(vdd), .A(_6144_), .B(_6138_), .C(_6145_), .Y(_4569__7_) );
NOR2X1 NOR2X1_1047 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe69), .B(_4594__bF_buf2), .Y(_6146_) );
INVX4 INVX4_107 ( .gnd(gnd), .vdd(vdd), .A(_6146_), .Y(_6147_) );
INVX1 INVX1_377 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_232_), .Y(_6148_) );
NOR2X1 NOR2X1_1048 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_k_0_), .B(micro_hash_ucr_2_x_0_), .Y(_6149_) );
NAND2X1 NAND2X1_820 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_k_0_), .B(micro_hash_ucr_2_x_0_), .Y(_6150_) );
INVX8 INVX8_184 ( .gnd(gnd), .vdd(vdd), .A(_6150_), .Y(_6151_) );
OAI21X1 OAI21X1_1703 ( .gnd(gnd), .vdd(vdd), .A(_6151_), .B(_6149_), .C(_6148_), .Y(_6152_) );
NOR2X1 NOR2X1_1049 ( .gnd(gnd), .vdd(vdd), .A(_6149_), .B(_6151_), .Y(_6153_) );
INVX8 INVX8_185 ( .gnd(gnd), .vdd(vdd), .A(_6153__bF_buf5), .Y(_6154_) );
NOR2X1 NOR2X1_1050 ( .gnd(gnd), .vdd(vdd), .A(_6148_), .B(_6154__bF_buf3), .Y(_6155_) );
INVX2 INVX2_221 ( .gnd(gnd), .vdd(vdd), .A(_6155_), .Y(_6156_) );
NAND2X1 NAND2X1_821 ( .gnd(gnd), .vdd(vdd), .A(_6152_), .B(_6156_), .Y(_6157_) );
OAI21X1 OAI21X1_1704 ( .gnd(gnd), .vdd(vdd), .A(_6151_), .B(_6149_), .C(_5026_), .Y(_6158_) );
NOR2X1 NOR2X1_1051 ( .gnd(gnd), .vdd(vdd), .A(_5026_), .B(_6154__bF_buf2), .Y(_6159_) );
INVX2 INVX2_222 ( .gnd(gnd), .vdd(vdd), .A(_6159_), .Y(_6160_) );
NAND2X1 NAND2X1_822 ( .gnd(gnd), .vdd(vdd), .A(_6158_), .B(_6160_), .Y(_6161_) );
INVX1 INVX1_378 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_32_), .Y(_6162_) );
OAI21X1 OAI21X1_1705 ( .gnd(gnd), .vdd(vdd), .A(_6151_), .B(_6149_), .C(_6162_), .Y(_6163_) );
NAND2X1 NAND2X1_823 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_32_), .B(_6153__bF_buf4), .Y(_6164_) );
AOI21X1 AOI21X1_1121 ( .gnd(gnd), .vdd(vdd), .A(_6163_), .B(_6164_), .C(_5127__bF_buf1), .Y(_6165_) );
NOR2X1 NOR2X1_1052 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_8_), .B(_6153__bF_buf3), .Y(_6166_) );
AND2X2 AND2X2_436 ( .gnd(gnd), .vdd(vdd), .A(_6153__bF_buf2), .B(micro_hash_ucr_2_Wx_8_), .Y(_6167_) );
OAI21X1 OAI21X1_1706 ( .gnd(gnd), .vdd(vdd), .A(_6167_), .B(_6166_), .C(micro_hash_ucr_2_pipe10), .Y(_6168_) );
INVX1 INVX1_379 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_0_), .Y(_6169_) );
NOR2X1 NOR2X1_1053 ( .gnd(gnd), .vdd(vdd), .A(_6169_), .B(_6154__bF_buf1), .Y(_6170_) );
OAI21X1 OAI21X1_1707 ( .gnd(gnd), .vdd(vdd), .A(_6153__bF_buf1), .B(micro_hash_ucr_2_Wx_0_), .C(micro_hash_ucr_2_pipe8), .Y(_6171_) );
NOR2X1 NOR2X1_1054 ( .gnd(gnd), .vdd(vdd), .A(_6171_), .B(_6170_), .Y(_6172_) );
NOR2X1 NOR2X1_1055 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_0_bF_buf0_), .B(micro_hash_ucr_2_pipe6), .Y(_6173_) );
OAI21X1 OAI21X1_1708 ( .gnd(gnd), .vdd(vdd), .A(_5134_), .B(H_2_16_), .C(_5135_), .Y(_6174_) );
OAI21X1 OAI21X1_1709 ( .gnd(gnd), .vdd(vdd), .A(_6174_), .B(_6173_), .C(_5133_), .Y(_6175_) );
OAI21X1 OAI21X1_1710 ( .gnd(gnd), .vdd(vdd), .A(_6172_), .B(_6175_), .C(_6168_), .Y(_6176_) );
XOR2X1 XOR2X1_88 ( .gnd(gnd), .vdd(vdd), .A(_6153__bF_buf0), .B(micro_hash_ucr_2_Wx_16_), .Y(_6177_) );
AOI21X1 AOI21X1_1122 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe12_bF_buf0), .B(_6177_), .C(micro_hash_ucr_2_pipe14_bF_buf1), .Y(_6178_) );
OAI21X1 OAI21X1_1711 ( .gnd(gnd), .vdd(vdd), .A(_6176_), .B(micro_hash_ucr_2_pipe12_bF_buf3), .C(_6178_), .Y(_6179_) );
NOR2X1 NOR2X1_1056 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_24_), .B(_6153__bF_buf5), .Y(_6180_) );
INVX1 INVX1_380 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_24_), .Y(_6181_) );
NOR2X1 NOR2X1_1057 ( .gnd(gnd), .vdd(vdd), .A(_6181_), .B(_6154__bF_buf0), .Y(_6182_) );
OAI21X1 OAI21X1_1712 ( .gnd(gnd), .vdd(vdd), .A(_6182_), .B(_6180_), .C(micro_hash_ucr_2_pipe14_bF_buf0), .Y(_6183_) );
AOI21X1 AOI21X1_1123 ( .gnd(gnd), .vdd(vdd), .A(_6183_), .B(_6179_), .C(micro_hash_ucr_2_pipe16_bF_buf0), .Y(_6184_) );
OAI21X1 OAI21X1_1713 ( .gnd(gnd), .vdd(vdd), .A(_6184_), .B(_6165_), .C(_5122__bF_buf0), .Y(_6185_) );
NOR2X1 NOR2X1_1058 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_40_), .B(_6153__bF_buf4), .Y(_6186_) );
NAND2X1 NAND2X1_824 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_40_), .B(_6153__bF_buf3), .Y(_6187_) );
INVX1 INVX1_381 ( .gnd(gnd), .vdd(vdd), .A(_6187_), .Y(_6188_) );
OAI21X1 OAI21X1_1714 ( .gnd(gnd), .vdd(vdd), .A(_6188_), .B(_6186_), .C(micro_hash_ucr_2_pipe18_bF_buf4), .Y(_6189_) );
NAND2X1 NAND2X1_825 ( .gnd(gnd), .vdd(vdd), .A(_6189_), .B(_6185_), .Y(_6190_) );
NOR2X1 NOR2X1_1059 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe20_bF_buf0), .B(_6190_), .Y(_6191_) );
AND2X2 AND2X2_437 ( .gnd(gnd), .vdd(vdd), .A(_6153__bF_buf2), .B(micro_hash_ucr_2_Wx_48_), .Y(_6192_) );
OAI21X1 OAI21X1_1715 ( .gnd(gnd), .vdd(vdd), .A(_6153__bF_buf1), .B(micro_hash_ucr_2_Wx_48_), .C(micro_hash_ucr_2_pipe20_bF_buf3), .Y(_6193_) );
OAI21X1 OAI21X1_1716 ( .gnd(gnd), .vdd(vdd), .A(_6192_), .B(_6193_), .C(_5121__bF_buf1), .Y(_6194_) );
NOR2X1 NOR2X1_1060 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_56_), .B(_6153__bF_buf0), .Y(_6195_) );
NOR2X1 NOR2X1_1061 ( .gnd(gnd), .vdd(vdd), .A(_5004_), .B(_6154__bF_buf3), .Y(_6196_) );
OAI21X1 OAI21X1_1717 ( .gnd(gnd), .vdd(vdd), .A(_6196_), .B(_6195_), .C(micro_hash_ucr_2_pipe22_bF_buf3), .Y(_6197_) );
OAI21X1 OAI21X1_1718 ( .gnd(gnd), .vdd(vdd), .A(_6191_), .B(_6194_), .C(_6197_), .Y(_6198_) );
NAND2X1 NAND2X1_826 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_64_), .B(_6153__bF_buf5), .Y(_6199_) );
OAI21X1 OAI21X1_1719 ( .gnd(gnd), .vdd(vdd), .A(_6151_), .B(_6149_), .C(_5050_), .Y(_6200_) );
AOI21X1 AOI21X1_1124 ( .gnd(gnd), .vdd(vdd), .A(_6200_), .B(_6199_), .C(_5116__bF_buf3), .Y(_6201_) );
AOI21X1 AOI21X1_1125 ( .gnd(gnd), .vdd(vdd), .A(_5116__bF_buf2), .B(_6198_), .C(_6201_), .Y(_6202_) );
NAND2X1 NAND2X1_827 ( .gnd(gnd), .vdd(vdd), .A(_5117__bF_buf2), .B(_6202_), .Y(_6203_) );
OAI21X1 OAI21X1_1720 ( .gnd(gnd), .vdd(vdd), .A(_5117__bF_buf1), .B(_6161_), .C(_6203_), .Y(_6204_) );
NOR2X1 NOR2X1_1062 ( .gnd(gnd), .vdd(vdd), .A(_4935_), .B(_6154__bF_buf2), .Y(_6205_) );
NOR2X1 NOR2X1_1063 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_80_), .B(_6153__bF_buf4), .Y(_6206_) );
OAI21X1 OAI21X1_1721 ( .gnd(gnd), .vdd(vdd), .A(_6205_), .B(_6206_), .C(micro_hash_ucr_2_pipe28_bF_buf0), .Y(_6207_) );
OAI21X1 OAI21X1_1722 ( .gnd(gnd), .vdd(vdd), .A(_6204_), .B(micro_hash_ucr_2_pipe28_bF_buf3), .C(_6207_), .Y(_6208_) );
OAI21X1 OAI21X1_1723 ( .gnd(gnd), .vdd(vdd), .A(_6151_), .B(_6149_), .C(_4975_), .Y(_6209_) );
NOR2X1 NOR2X1_1064 ( .gnd(gnd), .vdd(vdd), .A(_4975_), .B(_6154__bF_buf1), .Y(_6210_) );
NOR2X1 NOR2X1_1065 ( .gnd(gnd), .vdd(vdd), .A(_5110__bF_buf3), .B(_6210_), .Y(_6211_) );
AOI21X1 AOI21X1_1126 ( .gnd(gnd), .vdd(vdd), .A(_6209_), .B(_6211_), .C(micro_hash_ucr_2_pipe32_bF_buf0), .Y(_6212_) );
OAI21X1 OAI21X1_1724 ( .gnd(gnd), .vdd(vdd), .A(_6208_), .B(micro_hash_ucr_2_pipe30_bF_buf4), .C(_6212_), .Y(_6213_) );
NOR2X1 NOR2X1_1066 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_96_), .B(_6153__bF_buf3), .Y(_6214_) );
NOR2X1 NOR2X1_1067 ( .gnd(gnd), .vdd(vdd), .A(_4840_), .B(_6154__bF_buf0), .Y(_6215_) );
OAI21X1 OAI21X1_1725 ( .gnd(gnd), .vdd(vdd), .A(_6215_), .B(_6214_), .C(micro_hash_ucr_2_pipe32_bF_buf3), .Y(_6216_) );
NAND3X1 NAND3X1_299 ( .gnd(gnd), .vdd(vdd), .A(_5109__bF_buf4), .B(_6216_), .C(_6213_), .Y(_6217_) );
NOR2X1 NOR2X1_1068 ( .gnd(gnd), .vdd(vdd), .A(_4869_), .B(_6154__bF_buf3), .Y(_6218_) );
OAI21X1 OAI21X1_1726 ( .gnd(gnd), .vdd(vdd), .A(_6153__bF_buf2), .B(micro_hash_ucr_2_Wx_104_), .C(micro_hash_ucr_2_pipe34_bF_buf3), .Y(_6219_) );
OAI21X1 OAI21X1_1727 ( .gnd(gnd), .vdd(vdd), .A(_6218_), .B(_6219_), .C(_6217_), .Y(_6220_) );
XNOR2X1 XNOR2X1_212 ( .gnd(gnd), .vdd(vdd), .A(_6153__bF_buf1), .B(micro_hash_ucr_2_Wx_112_), .Y(_6221_) );
AOI21X1 AOI21X1_1127 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe36_bF_buf3), .B(_6221_), .C(micro_hash_ucr_2_pipe38_bF_buf2), .Y(_6222_) );
OAI21X1 OAI21X1_1728 ( .gnd(gnd), .vdd(vdd), .A(_6220_), .B(micro_hash_ucr_2_pipe36_bF_buf2), .C(_6222_), .Y(_6223_) );
NOR2X1 NOR2X1_1069 ( .gnd(gnd), .vdd(vdd), .A(_4754_), .B(_6154__bF_buf2), .Y(_6224_) );
OAI21X1 OAI21X1_1729 ( .gnd(gnd), .vdd(vdd), .A(_6153__bF_buf0), .B(micro_hash_ucr_2_Wx_120_), .C(micro_hash_ucr_2_pipe38_bF_buf1), .Y(_6225_) );
OAI21X1 OAI21X1_1730 ( .gnd(gnd), .vdd(vdd), .A(_6224_), .B(_6225_), .C(_6223_), .Y(_6226_) );
NOR2X1 NOR2X1_1070 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_128_), .B(_6153__bF_buf5), .Y(_6227_) );
NOR2X1 NOR2X1_1071 ( .gnd(gnd), .vdd(vdd), .A(_4781_), .B(_6154__bF_buf1), .Y(_6228_) );
OAI21X1 OAI21X1_1731 ( .gnd(gnd), .vdd(vdd), .A(_6228_), .B(_6227_), .C(micro_hash_ucr_2_pipe40_bF_buf3), .Y(_6229_) );
OAI21X1 OAI21X1_1732 ( .gnd(gnd), .vdd(vdd), .A(_6226_), .B(micro_hash_ucr_2_pipe40_bF_buf2), .C(_6229_), .Y(_6230_) );
NOR2X1 NOR2X1_1072 ( .gnd(gnd), .vdd(vdd), .A(_4976_), .B(_6154__bF_buf0), .Y(_6231_) );
OAI21X1 OAI21X1_1733 ( .gnd(gnd), .vdd(vdd), .A(_6153__bF_buf4), .B(micro_hash_ucr_2_Wx_136_), .C(micro_hash_ucr_2_pipe42_bF_buf1), .Y(_6232_) );
OAI22X1 OAI22X1_94 ( .gnd(gnd), .vdd(vdd), .A(_6231_), .B(_6232_), .C(_6230_), .D(micro_hash_ucr_2_pipe42_bF_buf0), .Y(_6233_) );
NOR2X1 NOR2X1_1073 ( .gnd(gnd), .vdd(vdd), .A(_4811_), .B(_6154__bF_buf3), .Y(_6234_) );
OAI21X1 OAI21X1_1734 ( .gnd(gnd), .vdd(vdd), .A(_6153__bF_buf3), .B(micro_hash_ucr_2_Wx_144_), .C(micro_hash_ucr_2_pipe44_bF_buf0), .Y(_6235_) );
OAI21X1 OAI21X1_1735 ( .gnd(gnd), .vdd(vdd), .A(_6234_), .B(_6235_), .C(_5097__bF_buf1), .Y(_6236_) );
AOI21X1 AOI21X1_1128 ( .gnd(gnd), .vdd(vdd), .A(_5099__bF_buf3), .B(_6233_), .C(_6236_), .Y(_6237_) );
NOR2X1 NOR2X1_1074 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_152_), .B(_6153__bF_buf2), .Y(_6238_) );
NOR2X1 NOR2X1_1075 ( .gnd(gnd), .vdd(vdd), .A(_4697_), .B(_6154__bF_buf2), .Y(_6239_) );
OAI21X1 OAI21X1_1736 ( .gnd(gnd), .vdd(vdd), .A(_6239_), .B(_6238_), .C(micro_hash_ucr_2_pipe46_bF_buf2), .Y(_6240_) );
NAND2X1 NAND2X1_828 ( .gnd(gnd), .vdd(vdd), .A(_5092__bF_buf1), .B(_6240_), .Y(_6241_) );
OAI21X1 OAI21X1_1737 ( .gnd(gnd), .vdd(vdd), .A(_6153__bF_buf1), .B(micro_hash_ucr_2_Wx_160_), .C(micro_hash_ucr_2_pipe48_bF_buf4), .Y(_6242_) );
AOI21X1 AOI21X1_1129 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_160_), .B(_6153__bF_buf0), .C(_6242_), .Y(_6243_) );
NOR2X1 NOR2X1_1076 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe50_bF_buf1), .B(_6243_), .Y(_6244_) );
OAI21X1 OAI21X1_1738 ( .gnd(gnd), .vdd(vdd), .A(_6237_), .B(_6241_), .C(_6244_), .Y(_6245_) );
XOR2X1 XOR2X1_89 ( .gnd(gnd), .vdd(vdd), .A(_6153__bF_buf5), .B(micro_hash_ucr_2_Wx_168_), .Y(_6246_) );
OAI21X1 OAI21X1_1739 ( .gnd(gnd), .vdd(vdd), .A(_5093__bF_buf1), .B(_6246_), .C(_6245_), .Y(_6247_) );
OAI21X1 OAI21X1_1740 ( .gnd(gnd), .vdd(vdd), .A(_6151_), .B(_6149_), .C(_4782_), .Y(_6248_) );
NOR2X1 NOR2X1_1077 ( .gnd(gnd), .vdd(vdd), .A(_4782_), .B(_6154__bF_buf1), .Y(_6249_) );
NOR2X1 NOR2X1_1078 ( .gnd(gnd), .vdd(vdd), .A(_5091__bF_buf4), .B(_6249_), .Y(_6250_) );
AOI21X1 AOI21X1_1130 ( .gnd(gnd), .vdd(vdd), .A(_6248_), .B(_6250_), .C(micro_hash_ucr_2_pipe54_bF_buf3), .Y(_6251_) );
OAI21X1 OAI21X1_1741 ( .gnd(gnd), .vdd(vdd), .A(_6247_), .B(micro_hash_ucr_2_pipe52_bF_buf3), .C(_6251_), .Y(_6252_) );
NOR2X1 NOR2X1_1079 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_184_), .B(_6153__bF_buf4), .Y(_6253_) );
AND2X2 AND2X2_438 ( .gnd(gnd), .vdd(vdd), .A(_6153__bF_buf3), .B(micro_hash_ucr_2_Wx_184_), .Y(_6254_) );
OAI21X1 OAI21X1_1742 ( .gnd(gnd), .vdd(vdd), .A(_6254_), .B(_6253_), .C(micro_hash_ucr_2_pipe54_bF_buf2), .Y(_6255_) );
NAND3X1 NAND3X1_300 ( .gnd(gnd), .vdd(vdd), .A(_5087__bF_buf1), .B(_6255_), .C(_6252_), .Y(_6256_) );
NOR2X1 NOR2X1_1080 ( .gnd(gnd), .vdd(vdd), .A(_4812_), .B(_6154__bF_buf0), .Y(_6257_) );
OAI21X1 OAI21X1_1743 ( .gnd(gnd), .vdd(vdd), .A(_6153__bF_buf2), .B(micro_hash_ucr_2_Wx_192_), .C(micro_hash_ucr_2_pipe56_bF_buf1), .Y(_6258_) );
OAI21X1 OAI21X1_1744 ( .gnd(gnd), .vdd(vdd), .A(_6257_), .B(_6258_), .C(_6256_), .Y(_6259_) );
OAI21X1 OAI21X1_1745 ( .gnd(gnd), .vdd(vdd), .A(_6151_), .B(_6149_), .C(_4698_), .Y(_6260_) );
NOR2X1 NOR2X1_1081 ( .gnd(gnd), .vdd(vdd), .A(_4698_), .B(_6154__bF_buf3), .Y(_6261_) );
INVX1 INVX1_382 ( .gnd(gnd), .vdd(vdd), .A(_6261_), .Y(_6262_) );
NAND2X1 NAND2X1_829 ( .gnd(gnd), .vdd(vdd), .A(_6260_), .B(_6262_), .Y(_6263_) );
AOI21X1 AOI21X1_1131 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe58_bF_buf3), .B(_6263_), .C(micro_hash_ucr_2_pipe60_bF_buf4), .Y(_6264_) );
OAI21X1 OAI21X1_1746 ( .gnd(gnd), .vdd(vdd), .A(_6259_), .B(micro_hash_ucr_2_pipe58_bF_buf2), .C(_6264_), .Y(_6265_) );
AND2X2 AND2X2_439 ( .gnd(gnd), .vdd(vdd), .A(_6153__bF_buf1), .B(micro_hash_ucr_2_Wx_208_), .Y(_6266_) );
OAI21X1 OAI21X1_1747 ( .gnd(gnd), .vdd(vdd), .A(_6153__bF_buf0), .B(micro_hash_ucr_2_Wx_208_), .C(micro_hash_ucr_2_pipe60_bF_buf3), .Y(_6267_) );
OAI21X1 OAI21X1_1748 ( .gnd(gnd), .vdd(vdd), .A(_6266_), .B(_6267_), .C(_6265_), .Y(_6268_) );
NOR2X1 NOR2X1_1082 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_216_), .B(_6153__bF_buf5), .Y(_6269_) );
NOR2X1 NOR2X1_1083 ( .gnd(gnd), .vdd(vdd), .A(_4726_), .B(_6154__bF_buf2), .Y(_6270_) );
OAI21X1 OAI21X1_1749 ( .gnd(gnd), .vdd(vdd), .A(_6270_), .B(_6269_), .C(micro_hash_ucr_2_pipe62_bF_buf4), .Y(_6271_) );
OAI21X1 OAI21X1_1750 ( .gnd(gnd), .vdd(vdd), .A(_6268_), .B(micro_hash_ucr_2_pipe62_bF_buf3), .C(_6271_), .Y(_6272_) );
AND2X2 AND2X2_440 ( .gnd(gnd), .vdd(vdd), .A(_6153__bF_buf4), .B(micro_hash_ucr_2_Wx_224_), .Y(_6273_) );
OAI21X1 OAI21X1_1751 ( .gnd(gnd), .vdd(vdd), .A(_6153__bF_buf3), .B(micro_hash_ucr_2_Wx_224_), .C(micro_hash_ucr_2_pipe64_bF_buf1), .Y(_6274_) );
OAI22X1 OAI22X1_95 ( .gnd(gnd), .vdd(vdd), .A(_6273_), .B(_6274_), .C(_6272_), .D(micro_hash_ucr_2_pipe64_bF_buf0), .Y(_6275_) );
NAND2X1 NAND2X1_830 ( .gnd(gnd), .vdd(vdd), .A(_5074__bF_buf0), .B(_6275_), .Y(_6276_) );
OAI21X1 OAI21X1_1752 ( .gnd(gnd), .vdd(vdd), .A(_5074__bF_buf3), .B(_6157_), .C(_6276_), .Y(_6277_) );
NOR2X1 NOR2X1_1084 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_240_), .B(_6153__bF_buf2), .Y(_6278_) );
AND2X2 AND2X2_441 ( .gnd(gnd), .vdd(vdd), .A(_6153__bF_buf1), .B(micro_hash_ucr_2_Wx_240_), .Y(_6279_) );
OAI21X1 OAI21X1_1753 ( .gnd(gnd), .vdd(vdd), .A(_6279_), .B(_6278_), .C(micro_hash_ucr_2_pipe68), .Y(_6280_) );
OAI21X1 OAI21X1_1754 ( .gnd(gnd), .vdd(vdd), .A(_6277_), .B(micro_hash_ucr_2_pipe68), .C(_6280_), .Y(_6281_) );
INVX2 INVX2_223 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_248_), .Y(_6282_) );
AOI21X1 AOI21X1_1132 ( .gnd(gnd), .vdd(vdd), .A(_6282_), .B(_6154__bF_buf1), .C(_4594__bF_buf1), .Y(_6283_) );
OAI21X1 OAI21X1_1755 ( .gnd(gnd), .vdd(vdd), .A(_6282_), .B(_6154__bF_buf0), .C(_6283_), .Y(_6284_) );
AOI22X1 AOI22X1_51 ( .gnd(gnd), .vdd(vdd), .A(_6147_), .B(_6284_), .C(_6281_), .D(_5073__bF_buf1), .Y(_4493__0_) );
INVX1 INVX1_383 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_9_), .Y(_6285_) );
NOR2X1 NOR2X1_1085 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_k_1_), .B(micro_hash_ucr_2_x_1_), .Y(_6286_) );
AND2X2 AND2X2_442 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_k_1_), .B(micro_hash_ucr_2_x_1_), .Y(_6287_) );
NOR2X1 NOR2X1_1086 ( .gnd(gnd), .vdd(vdd), .A(_6286_), .B(_6287_), .Y(_6288_) );
AND2X2 AND2X2_443 ( .gnd(gnd), .vdd(vdd), .A(_6288_), .B(_6151_), .Y(_6289_) );
NOR2X1 NOR2X1_1087 ( .gnd(gnd), .vdd(vdd), .A(_6151_), .B(_6288_), .Y(_6290_) );
OAI21X1 OAI21X1_1756 ( .gnd(gnd), .vdd(vdd), .A(_6289_), .B(_6290_), .C(_6285_), .Y(_6291_) );
INVX1 INVX1_384 ( .gnd(gnd), .vdd(vdd), .A(_6291_), .Y(_6292_) );
NOR2X1 NOR2X1_1088 ( .gnd(gnd), .vdd(vdd), .A(_6290_), .B(_6289_), .Y(_6293_) );
INVX8 INVX8_186 ( .gnd(gnd), .vdd(vdd), .A(_6293__bF_buf4), .Y(_6294_) );
NOR2X1 NOR2X1_1089 ( .gnd(gnd), .vdd(vdd), .A(_6285_), .B(_6294__bF_buf4), .Y(_6295_) );
NOR2X1 NOR2X1_1090 ( .gnd(gnd), .vdd(vdd), .A(_6292_), .B(_6295_), .Y(_6296_) );
XNOR2X1 XNOR2X1_213 ( .gnd(gnd), .vdd(vdd), .A(_6296_), .B(_6167_), .Y(_6297_) );
NAND2X1 NAND2X1_831 ( .gnd(gnd), .vdd(vdd), .A(H_2_17_), .B(micro_hash_ucr_2_pipe6), .Y(_6298_) );
OAI21X1 OAI21X1_1757 ( .gnd(gnd), .vdd(vdd), .A(_5255_), .B(micro_hash_ucr_2_pipe6), .C(_6298_), .Y(_6299_) );
NOR2X1 NOR2X1_1091 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_1_), .B(_6293__bF_buf3), .Y(_6300_) );
INVX1 INVX1_385 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_1_), .Y(_6301_) );
NOR2X1 NOR2X1_1092 ( .gnd(gnd), .vdd(vdd), .A(_6301_), .B(_6294__bF_buf3), .Y(_6302_) );
NOR2X1 NOR2X1_1093 ( .gnd(gnd), .vdd(vdd), .A(_6300_), .B(_6302_), .Y(_6303_) );
AND2X2 AND2X2_444 ( .gnd(gnd), .vdd(vdd), .A(_6303_), .B(_6170_), .Y(_6304_) );
NOR2X1 NOR2X1_1094 ( .gnd(gnd), .vdd(vdd), .A(_6170_), .B(_6303_), .Y(_6305_) );
OAI21X1 OAI21X1_1758 ( .gnd(gnd), .vdd(vdd), .A(_6305_), .B(_6304_), .C(micro_hash_ucr_2_pipe8), .Y(_6306_) );
OAI21X1 OAI21X1_1759 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe8), .B(_6299_), .C(_6306_), .Y(_6307_) );
MUX2X1 MUX2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_6307_), .B(_6297_), .S(_5133_), .Y(_6308_) );
NAND2X1 NAND2X1_832 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_16_), .B(_6153__bF_buf0), .Y(_6309_) );
NOR2X1 NOR2X1_1095 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_17_), .B(_6293__bF_buf2), .Y(_6310_) );
INVX1 INVX1_386 ( .gnd(gnd), .vdd(vdd), .A(_6310_), .Y(_6311_) );
NAND2X1 NAND2X1_833 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_17_), .B(_6293__bF_buf1), .Y(_6312_) );
NAND2X1 NAND2X1_834 ( .gnd(gnd), .vdd(vdd), .A(_6312_), .B(_6311_), .Y(_6313_) );
AND2X2 AND2X2_445 ( .gnd(gnd), .vdd(vdd), .A(_6313_), .B(_6309_), .Y(_6314_) );
NOR2X1 NOR2X1_1096 ( .gnd(gnd), .vdd(vdd), .A(_6309_), .B(_6313_), .Y(_6315_) );
OAI21X1 OAI21X1_1760 ( .gnd(gnd), .vdd(vdd), .A(_6314_), .B(_6315_), .C(micro_hash_ucr_2_pipe12_bF_buf2), .Y(_6316_) );
OAI21X1 OAI21X1_1761 ( .gnd(gnd), .vdd(vdd), .A(_6308_), .B(micro_hash_ucr_2_pipe12_bF_buf1), .C(_6316_), .Y(_6317_) );
INVX1 INVX1_387 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_25_), .Y(_6318_) );
OAI21X1 OAI21X1_1762 ( .gnd(gnd), .vdd(vdd), .A(_6289_), .B(_6290_), .C(_6318_), .Y(_6319_) );
INVX1 INVX1_388 ( .gnd(gnd), .vdd(vdd), .A(_6319_), .Y(_6320_) );
NOR2X1 NOR2X1_1097 ( .gnd(gnd), .vdd(vdd), .A(_6318_), .B(_6294__bF_buf2), .Y(_6321_) );
NOR2X1 NOR2X1_1098 ( .gnd(gnd), .vdd(vdd), .A(_6320_), .B(_6321_), .Y(_6322_) );
XOR2X1 XOR2X1_90 ( .gnd(gnd), .vdd(vdd), .A(_6322_), .B(_6182_), .Y(_6323_) );
NAND2X1 NAND2X1_835 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe14_bF_buf4), .B(_6323_), .Y(_6324_) );
OAI21X1 OAI21X1_1763 ( .gnd(gnd), .vdd(vdd), .A(_6317_), .B(micro_hash_ucr_2_pipe14_bF_buf3), .C(_6324_), .Y(_6325_) );
NOR2X1 NOR2X1_1099 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_33_), .B(_6293__bF_buf0), .Y(_6326_) );
INVX1 INVX1_389 ( .gnd(gnd), .vdd(vdd), .A(_6326_), .Y(_6327_) );
NAND2X1 NAND2X1_836 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_33_), .B(_6293__bF_buf4), .Y(_6328_) );
NAND2X1 NAND2X1_837 ( .gnd(gnd), .vdd(vdd), .A(_6328_), .B(_6327_), .Y(_6329_) );
NOR2X1 NOR2X1_1100 ( .gnd(gnd), .vdd(vdd), .A(_6164_), .B(_6329_), .Y(_6330_) );
AND2X2 AND2X2_446 ( .gnd(gnd), .vdd(vdd), .A(_6329_), .B(_6164_), .Y(_6331_) );
OAI21X1 OAI21X1_1764 ( .gnd(gnd), .vdd(vdd), .A(_6331_), .B(_6330_), .C(micro_hash_ucr_2_pipe16_bF_buf4), .Y(_6332_) );
OAI21X1 OAI21X1_1765 ( .gnd(gnd), .vdd(vdd), .A(_6325_), .B(micro_hash_ucr_2_pipe16_bF_buf3), .C(_6332_), .Y(_6333_) );
NAND2X1 NAND2X1_838 ( .gnd(gnd), .vdd(vdd), .A(_5122__bF_buf4), .B(_6333_), .Y(_6334_) );
INVX1 INVX1_390 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_41_), .Y(_6335_) );
OAI21X1 OAI21X1_1766 ( .gnd(gnd), .vdd(vdd), .A(_6289_), .B(_6290_), .C(_6335_), .Y(_6336_) );
INVX1 INVX1_391 ( .gnd(gnd), .vdd(vdd), .A(_6336_), .Y(_6337_) );
NOR2X1 NOR2X1_1101 ( .gnd(gnd), .vdd(vdd), .A(_6335_), .B(_6294__bF_buf1), .Y(_6338_) );
NOR2X1 NOR2X1_1102 ( .gnd(gnd), .vdd(vdd), .A(_6337_), .B(_6338_), .Y(_6339_) );
XNOR2X1 XNOR2X1_214 ( .gnd(gnd), .vdd(vdd), .A(_6339_), .B(_6187_), .Y(_6340_) );
OAI21X1 OAI21X1_1767 ( .gnd(gnd), .vdd(vdd), .A(_5122__bF_buf3), .B(_6340_), .C(_6334_), .Y(_6341_) );
INVX2 INVX2_224 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_49_), .Y(_6342_) );
XNOR2X1 XNOR2X1_215 ( .gnd(gnd), .vdd(vdd), .A(_6293__bF_buf3), .B(_6342_), .Y(_6343_) );
NAND2X1 NAND2X1_839 ( .gnd(gnd), .vdd(vdd), .A(_6192_), .B(_6343_), .Y(_6344_) );
NOR2X1 NOR2X1_1103 ( .gnd(gnd), .vdd(vdd), .A(_6192_), .B(_6343_), .Y(_6345_) );
NOR2X1 NOR2X1_1104 ( .gnd(gnd), .vdd(vdd), .A(_5123__bF_buf2), .B(_6345_), .Y(_6346_) );
AOI21X1 AOI21X1_1133 ( .gnd(gnd), .vdd(vdd), .A(_6344_), .B(_6346_), .C(micro_hash_ucr_2_pipe22_bF_buf2), .Y(_6347_) );
OAI21X1 OAI21X1_1768 ( .gnd(gnd), .vdd(vdd), .A(_6341_), .B(micro_hash_ucr_2_pipe20_bF_buf2), .C(_6347_), .Y(_6348_) );
INVX1 INVX1_392 ( .gnd(gnd), .vdd(vdd), .A(_6196_), .Y(_6349_) );
OAI21X1 OAI21X1_1769 ( .gnd(gnd), .vdd(vdd), .A(_6289_), .B(_6290_), .C(_5007_), .Y(_6350_) );
NOR2X1 NOR2X1_1105 ( .gnd(gnd), .vdd(vdd), .A(_5007_), .B(_6294__bF_buf0), .Y(_6351_) );
INVX2 INVX2_225 ( .gnd(gnd), .vdd(vdd), .A(_6351_), .Y(_6352_) );
NAND2X1 NAND2X1_840 ( .gnd(gnd), .vdd(vdd), .A(_6350_), .B(_6352_), .Y(_6353_) );
NOR2X1 NOR2X1_1106 ( .gnd(gnd), .vdd(vdd), .A(_6349_), .B(_6353_), .Y(_6354_) );
AOI21X1 AOI21X1_1134 ( .gnd(gnd), .vdd(vdd), .A(_6350_), .B(_6352_), .C(_6196_), .Y(_6355_) );
OAI21X1 OAI21X1_1770 ( .gnd(gnd), .vdd(vdd), .A(_6354_), .B(_6355_), .C(micro_hash_ucr_2_pipe22_bF_buf1), .Y(_6356_) );
AOI21X1 AOI21X1_1135 ( .gnd(gnd), .vdd(vdd), .A(_6356_), .B(_6348_), .C(micro_hash_ucr_2_pipe24_bF_buf3), .Y(_6357_) );
XNOR2X1 XNOR2X1_216 ( .gnd(gnd), .vdd(vdd), .A(_6293__bF_buf2), .B(micro_hash_ucr_2_Wx_65_), .Y(_6358_) );
NOR2X1 NOR2X1_1107 ( .gnd(gnd), .vdd(vdd), .A(_6199_), .B(_6358_), .Y(_6359_) );
INVX1 INVX1_393 ( .gnd(gnd), .vdd(vdd), .A(_6359_), .Y(_6360_) );
OAI21X1 OAI21X1_1771 ( .gnd(gnd), .vdd(vdd), .A(_5050_), .B(_6154__bF_buf3), .C(_6358_), .Y(_6361_) );
AOI21X1 AOI21X1_1136 ( .gnd(gnd), .vdd(vdd), .A(_6361_), .B(_6360_), .C(_5116__bF_buf1), .Y(_6362_) );
OAI21X1 OAI21X1_1772 ( .gnd(gnd), .vdd(vdd), .A(_6357_), .B(_6362_), .C(_5117__bF_buf0), .Y(_6363_) );
OAI21X1 OAI21X1_1773 ( .gnd(gnd), .vdd(vdd), .A(_6289_), .B(_6290_), .C(_5029_), .Y(_6364_) );
INVX1 INVX1_394 ( .gnd(gnd), .vdd(vdd), .A(_6364_), .Y(_6365_) );
NOR2X1 NOR2X1_1108 ( .gnd(gnd), .vdd(vdd), .A(_5029_), .B(_6294__bF_buf4), .Y(_6366_) );
NOR2X1 NOR2X1_1109 ( .gnd(gnd), .vdd(vdd), .A(_6365_), .B(_6366_), .Y(_6367_) );
XNOR2X1 XNOR2X1_217 ( .gnd(gnd), .vdd(vdd), .A(_6367_), .B(_6160_), .Y(_6368_) );
OAI21X1 OAI21X1_1774 ( .gnd(gnd), .vdd(vdd), .A(_5117__bF_buf4), .B(_6368_), .C(_6363_), .Y(_6369_) );
XNOR2X1 XNOR2X1_218 ( .gnd(gnd), .vdd(vdd), .A(_6293__bF_buf1), .B(_4938_), .Y(_6370_) );
XOR2X1 XOR2X1_91 ( .gnd(gnd), .vdd(vdd), .A(_6370_), .B(_6205_), .Y(_6371_) );
AOI21X1 AOI21X1_1137 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe28_bF_buf2), .B(_6371_), .C(micro_hash_ucr_2_pipe30_bF_buf3), .Y(_6372_) );
OAI21X1 OAI21X1_1775 ( .gnd(gnd), .vdd(vdd), .A(_6369_), .B(micro_hash_ucr_2_pipe28_bF_buf1), .C(_6372_), .Y(_6373_) );
INVX1 INVX1_395 ( .gnd(gnd), .vdd(vdd), .A(_6210_), .Y(_6374_) );
OAI21X1 OAI21X1_1776 ( .gnd(gnd), .vdd(vdd), .A(_6289_), .B(_6290_), .C(_4979_), .Y(_6375_) );
NOR2X1 NOR2X1_1110 ( .gnd(gnd), .vdd(vdd), .A(_4979_), .B(_6294__bF_buf3), .Y(_6376_) );
INVX2 INVX2_226 ( .gnd(gnd), .vdd(vdd), .A(_6376_), .Y(_6377_) );
NAND2X1 NAND2X1_841 ( .gnd(gnd), .vdd(vdd), .A(_6375_), .B(_6377_), .Y(_6378_) );
NOR2X1 NOR2X1_1111 ( .gnd(gnd), .vdd(vdd), .A(_6374_), .B(_6378_), .Y(_6379_) );
AOI21X1 AOI21X1_1138 ( .gnd(gnd), .vdd(vdd), .A(_6375_), .B(_6377_), .C(_6210_), .Y(_6380_) );
OAI21X1 OAI21X1_1777 ( .gnd(gnd), .vdd(vdd), .A(_6379_), .B(_6380_), .C(micro_hash_ucr_2_pipe30_bF_buf2), .Y(_6381_) );
AOI21X1 AOI21X1_1139 ( .gnd(gnd), .vdd(vdd), .A(_6381_), .B(_6373_), .C(micro_hash_ucr_2_pipe32_bF_buf2), .Y(_6382_) );
XNOR2X1 XNOR2X1_219 ( .gnd(gnd), .vdd(vdd), .A(_6293__bF_buf0), .B(_4843_), .Y(_6383_) );
NAND2X1 NAND2X1_842 ( .gnd(gnd), .vdd(vdd), .A(_6215_), .B(_6383_), .Y(_6384_) );
OR2X2 OR2X2_50 ( .gnd(gnd), .vdd(vdd), .A(_6383_), .B(_6215_), .Y(_6385_) );
AOI21X1 AOI21X1_1140 ( .gnd(gnd), .vdd(vdd), .A(_6384_), .B(_6385_), .C(_5111__bF_buf3), .Y(_6386_) );
OAI21X1 OAI21X1_1778 ( .gnd(gnd), .vdd(vdd), .A(_6382_), .B(_6386_), .C(_5109__bF_buf3), .Y(_6387_) );
OAI21X1 OAI21X1_1779 ( .gnd(gnd), .vdd(vdd), .A(_6289_), .B(_6290_), .C(_4872_), .Y(_6388_) );
INVX1 INVX1_396 ( .gnd(gnd), .vdd(vdd), .A(_6388_), .Y(_6389_) );
NOR2X1 NOR2X1_1112 ( .gnd(gnd), .vdd(vdd), .A(_4872_), .B(_6294__bF_buf2), .Y(_6390_) );
NOR2X1 NOR2X1_1113 ( .gnd(gnd), .vdd(vdd), .A(_6389_), .B(_6390_), .Y(_6391_) );
XOR2X1 XOR2X1_92 ( .gnd(gnd), .vdd(vdd), .A(_6391_), .B(_6218_), .Y(_6392_) );
OAI21X1 OAI21X1_1780 ( .gnd(gnd), .vdd(vdd), .A(_5109__bF_buf2), .B(_6392_), .C(_6387_), .Y(_6393_) );
NOR2X1 NOR2X1_1114 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe36_bF_buf1), .B(_6393_), .Y(_6394_) );
NOR2X1 NOR2X1_1115 ( .gnd(gnd), .vdd(vdd), .A(_4913_), .B(_6154__bF_buf2), .Y(_6395_) );
XNOR2X1 XNOR2X1_220 ( .gnd(gnd), .vdd(vdd), .A(_6293__bF_buf4), .B(_4916_), .Y(_6396_) );
NOR2X1 NOR2X1_1116 ( .gnd(gnd), .vdd(vdd), .A(_6395_), .B(_6396_), .Y(_6397_) );
NAND2X1 NAND2X1_843 ( .gnd(gnd), .vdd(vdd), .A(_6395_), .B(_6396_), .Y(_6398_) );
NAND2X1 NAND2X1_844 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe36_bF_buf0), .B(_6398_), .Y(_6399_) );
OAI21X1 OAI21X1_1781 ( .gnd(gnd), .vdd(vdd), .A(_6399_), .B(_6397_), .C(_5105__bF_buf0), .Y(_6400_) );
OAI21X1 OAI21X1_1782 ( .gnd(gnd), .vdd(vdd), .A(_6289_), .B(_6290_), .C(_4895_), .Y(_6401_) );
INVX1 INVX1_397 ( .gnd(gnd), .vdd(vdd), .A(_6401_), .Y(_6402_) );
NOR2X1 NOR2X1_1117 ( .gnd(gnd), .vdd(vdd), .A(_4895_), .B(_6294__bF_buf1), .Y(_6403_) );
NOR2X1 NOR2X1_1118 ( .gnd(gnd), .vdd(vdd), .A(_6402_), .B(_6403_), .Y(_6404_) );
XOR2X1 XOR2X1_93 ( .gnd(gnd), .vdd(vdd), .A(_6404_), .B(_6224_), .Y(_6405_) );
OAI22X1 OAI22X1_96 ( .gnd(gnd), .vdd(vdd), .A(_5105__bF_buf4), .B(_6405_), .C(_6394_), .D(_6400_), .Y(_6406_) );
XNOR2X1 XNOR2X1_221 ( .gnd(gnd), .vdd(vdd), .A(_6293__bF_buf3), .B(_4785_), .Y(_6407_) );
XOR2X1 XOR2X1_94 ( .gnd(gnd), .vdd(vdd), .A(_6407_), .B(_6228_), .Y(_6408_) );
AOI21X1 AOI21X1_1141 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe40_bF_buf1), .B(_6408_), .C(micro_hash_ucr_2_pipe42_bF_buf3), .Y(_6409_) );
OAI21X1 OAI21X1_1783 ( .gnd(gnd), .vdd(vdd), .A(_6406_), .B(micro_hash_ucr_2_pipe40_bF_buf0), .C(_6409_), .Y(_6410_) );
XNOR2X1 XNOR2X1_222 ( .gnd(gnd), .vdd(vdd), .A(_6293__bF_buf2), .B(_4980_), .Y(_6411_) );
AND2X2 AND2X2_447 ( .gnd(gnd), .vdd(vdd), .A(_6411_), .B(_6231_), .Y(_6412_) );
NOR2X1 NOR2X1_1119 ( .gnd(gnd), .vdd(vdd), .A(_6231_), .B(_6411_), .Y(_6413_) );
OAI21X1 OAI21X1_1784 ( .gnd(gnd), .vdd(vdd), .A(_6412_), .B(_6413_), .C(micro_hash_ucr_2_pipe42_bF_buf2), .Y(_6414_) );
NAND3X1 NAND3X1_301 ( .gnd(gnd), .vdd(vdd), .A(_5099__bF_buf2), .B(_6414_), .C(_6410_), .Y(_6415_) );
XNOR2X1 XNOR2X1_223 ( .gnd(gnd), .vdd(vdd), .A(_6293__bF_buf1), .B(_4815_), .Y(_6416_) );
NAND2X1 NAND2X1_845 ( .gnd(gnd), .vdd(vdd), .A(_6234_), .B(_6416_), .Y(_6417_) );
INVX1 INVX1_398 ( .gnd(gnd), .vdd(vdd), .A(_6417_), .Y(_6418_) );
OAI21X1 OAI21X1_1785 ( .gnd(gnd), .vdd(vdd), .A(_6416_), .B(_6234_), .C(micro_hash_ucr_2_pipe44_bF_buf3), .Y(_6419_) );
OAI21X1 OAI21X1_1786 ( .gnd(gnd), .vdd(vdd), .A(_6418_), .B(_6419_), .C(_6415_), .Y(_6420_) );
XNOR2X1 XNOR2X1_224 ( .gnd(gnd), .vdd(vdd), .A(_6293__bF_buf0), .B(_4701_), .Y(_6421_) );
AND2X2 AND2X2_448 ( .gnd(gnd), .vdd(vdd), .A(_6421_), .B(_6239_), .Y(_6422_) );
NOR2X1 NOR2X1_1120 ( .gnd(gnd), .vdd(vdd), .A(_6239_), .B(_6421_), .Y(_6423_) );
OAI21X1 OAI21X1_1787 ( .gnd(gnd), .vdd(vdd), .A(_6422_), .B(_6423_), .C(micro_hash_ucr_2_pipe46_bF_buf1), .Y(_6424_) );
OAI21X1 OAI21X1_1788 ( .gnd(gnd), .vdd(vdd), .A(_6420_), .B(micro_hash_ucr_2_pipe46_bF_buf0), .C(_6424_), .Y(_6425_) );
NAND2X1 NAND2X1_846 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_160_), .B(_6153__bF_buf5), .Y(_6426_) );
XNOR2X1 XNOR2X1_225 ( .gnd(gnd), .vdd(vdd), .A(_6293__bF_buf4), .B(micro_hash_ucr_2_Wx_161_), .Y(_6427_) );
NOR2X1 NOR2X1_1121 ( .gnd(gnd), .vdd(vdd), .A(_6426_), .B(_6427_), .Y(_6428_) );
INVX1 INVX1_399 ( .gnd(gnd), .vdd(vdd), .A(_6428_), .Y(_6429_) );
AOI21X1 AOI21X1_1142 ( .gnd(gnd), .vdd(vdd), .A(_6426_), .B(_6427_), .C(_5092__bF_buf0), .Y(_6430_) );
AOI21X1 AOI21X1_1143 ( .gnd(gnd), .vdd(vdd), .A(_6430_), .B(_6429_), .C(micro_hash_ucr_2_pipe50_bF_buf0), .Y(_6431_) );
OAI21X1 OAI21X1_1789 ( .gnd(gnd), .vdd(vdd), .A(_6425_), .B(micro_hash_ucr_2_pipe48_bF_buf3), .C(_6431_), .Y(_6432_) );
NAND2X1 NAND2X1_847 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_168_), .B(_6153__bF_buf4), .Y(_6433_) );
OAI21X1 OAI21X1_1790 ( .gnd(gnd), .vdd(vdd), .A(_6289_), .B(_6290_), .C(_4728_), .Y(_6434_) );
NAND2X1 NAND2X1_848 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_169_), .B(_6293__bF_buf3), .Y(_6435_) );
NAND2X1 NAND2X1_849 ( .gnd(gnd), .vdd(vdd), .A(_6434_), .B(_6435_), .Y(_6436_) );
XOR2X1 XOR2X1_95 ( .gnd(gnd), .vdd(vdd), .A(_6436_), .B(_6433_), .Y(_6437_) );
OAI21X1 OAI21X1_1791 ( .gnd(gnd), .vdd(vdd), .A(_5093__bF_buf0), .B(_6437_), .C(_6432_), .Y(_6438_) );
XNOR2X1 XNOR2X1_226 ( .gnd(gnd), .vdd(vdd), .A(_6293__bF_buf2), .B(_4786_), .Y(_6439_) );
XOR2X1 XOR2X1_96 ( .gnd(gnd), .vdd(vdd), .A(_6439_), .B(_6249_), .Y(_6440_) );
AOI21X1 AOI21X1_1144 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe52_bF_buf2), .B(_6440_), .C(micro_hash_ucr_2_pipe54_bF_buf1), .Y(_6441_) );
OAI21X1 OAI21X1_1792 ( .gnd(gnd), .vdd(vdd), .A(_6438_), .B(micro_hash_ucr_2_pipe52_bF_buf1), .C(_6441_), .Y(_6442_) );
XNOR2X1 XNOR2X1_227 ( .gnd(gnd), .vdd(vdd), .A(_6293__bF_buf1), .B(_4844_), .Y(_6443_) );
AND2X2 AND2X2_449 ( .gnd(gnd), .vdd(vdd), .A(_6443_), .B(_6254_), .Y(_6444_) );
NOR2X1 NOR2X1_1122 ( .gnd(gnd), .vdd(vdd), .A(_6254_), .B(_6443_), .Y(_6445_) );
OAI21X1 OAI21X1_1793 ( .gnd(gnd), .vdd(vdd), .A(_6444_), .B(_6445_), .C(micro_hash_ucr_2_pipe54_bF_buf0), .Y(_6446_) );
NAND3X1 NAND3X1_302 ( .gnd(gnd), .vdd(vdd), .A(_5087__bF_buf0), .B(_6446_), .C(_6442_), .Y(_6447_) );
XNOR2X1 XNOR2X1_228 ( .gnd(gnd), .vdd(vdd), .A(_6293__bF_buf0), .B(_4816_), .Y(_6448_) );
NAND2X1 NAND2X1_850 ( .gnd(gnd), .vdd(vdd), .A(_6257_), .B(_6448_), .Y(_6449_) );
INVX1 INVX1_400 ( .gnd(gnd), .vdd(vdd), .A(_6449_), .Y(_6450_) );
OAI21X1 OAI21X1_1794 ( .gnd(gnd), .vdd(vdd), .A(_6448_), .B(_6257_), .C(micro_hash_ucr_2_pipe56_bF_buf0), .Y(_6451_) );
OAI21X1 OAI21X1_1795 ( .gnd(gnd), .vdd(vdd), .A(_6450_), .B(_6451_), .C(_6447_), .Y(_6452_) );
XNOR2X1 XNOR2X1_229 ( .gnd(gnd), .vdd(vdd), .A(_6293__bF_buf4), .B(_4702_), .Y(_6453_) );
NOR2X1 NOR2X1_1123 ( .gnd(gnd), .vdd(vdd), .A(_6261_), .B(_6453_), .Y(_6454_) );
AND2X2 AND2X2_450 ( .gnd(gnd), .vdd(vdd), .A(_6453_), .B(_6261_), .Y(_6455_) );
OAI21X1 OAI21X1_1796 ( .gnd(gnd), .vdd(vdd), .A(_6455_), .B(_6454_), .C(micro_hash_ucr_2_pipe58_bF_buf1), .Y(_6456_) );
OAI21X1 OAI21X1_1797 ( .gnd(gnd), .vdd(vdd), .A(_6452_), .B(micro_hash_ucr_2_pipe58_bF_buf0), .C(_6456_), .Y(_6457_) );
NAND2X1 NAND2X1_851 ( .gnd(gnd), .vdd(vdd), .A(_5080__bF_buf3), .B(_6457_), .Y(_6458_) );
NAND2X1 NAND2X1_852 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_208_), .B(_6153__bF_buf3), .Y(_6459_) );
NOR2X1 NOR2X1_1124 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_209_), .B(_6293__bF_buf3), .Y(_6460_) );
INVX1 INVX1_401 ( .gnd(gnd), .vdd(vdd), .A(_6460_), .Y(_6461_) );
NAND2X1 NAND2X1_853 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_209_), .B(_6293__bF_buf2), .Y(_6462_) );
NAND2X1 NAND2X1_854 ( .gnd(gnd), .vdd(vdd), .A(_6462_), .B(_6461_), .Y(_6463_) );
NOR2X1 NOR2X1_1125 ( .gnd(gnd), .vdd(vdd), .A(_6459_), .B(_6463_), .Y(_6464_) );
AOI21X1 AOI21X1_1145 ( .gnd(gnd), .vdd(vdd), .A(_6462_), .B(_6461_), .C(_6266_), .Y(_6465_) );
OAI21X1 OAI21X1_1798 ( .gnd(gnd), .vdd(vdd), .A(_6464_), .B(_6465_), .C(micro_hash_ucr_2_pipe60_bF_buf2), .Y(_6466_) );
NAND3X1 NAND3X1_303 ( .gnd(gnd), .vdd(vdd), .A(_5081__bF_buf3), .B(_6466_), .C(_6458_), .Y(_6467_) );
OAI21X1 OAI21X1_1799 ( .gnd(gnd), .vdd(vdd), .A(_6289_), .B(_6290_), .C(_4729_), .Y(_6468_) );
INVX1 INVX1_402 ( .gnd(gnd), .vdd(vdd), .A(_6468_), .Y(_6469_) );
NOR2X1 NOR2X1_1126 ( .gnd(gnd), .vdd(vdd), .A(_4729_), .B(_6294__bF_buf0), .Y(_6470_) );
NOR2X1 NOR2X1_1127 ( .gnd(gnd), .vdd(vdd), .A(_6469_), .B(_6470_), .Y(_6471_) );
AND2X2 AND2X2_451 ( .gnd(gnd), .vdd(vdd), .A(_6471_), .B(_6270_), .Y(_6472_) );
OAI21X1 OAI21X1_1800 ( .gnd(gnd), .vdd(vdd), .A(_6471_), .B(_6270_), .C(micro_hash_ucr_2_pipe62_bF_buf2), .Y(_6473_) );
OAI21X1 OAI21X1_1801 ( .gnd(gnd), .vdd(vdd), .A(_6472_), .B(_6473_), .C(_6467_), .Y(_6474_) );
NOR2X1 NOR2X1_1128 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe64_bF_buf4), .B(_6474_), .Y(_6475_) );
INVX2 INVX2_227 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_225_), .Y(_6476_) );
XNOR2X1 XNOR2X1_230 ( .gnd(gnd), .vdd(vdd), .A(_6293__bF_buf1), .B(_6476_), .Y(_6477_) );
OR2X2 OR2X2_51 ( .gnd(gnd), .vdd(vdd), .A(_6477_), .B(_6273_), .Y(_6478_) );
NAND2X1 NAND2X1_855 ( .gnd(gnd), .vdd(vdd), .A(_6273_), .B(_6477_), .Y(_6479_) );
AOI21X1 AOI21X1_1146 ( .gnd(gnd), .vdd(vdd), .A(_6479_), .B(_6478_), .C(_5079__bF_buf4), .Y(_6480_) );
OAI21X1 OAI21X1_1802 ( .gnd(gnd), .vdd(vdd), .A(_6475_), .B(_6480_), .C(_5074__bF_buf2), .Y(_6481_) );
INVX1 INVX1_403 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_233_), .Y(_6482_) );
OAI21X1 OAI21X1_1803 ( .gnd(gnd), .vdd(vdd), .A(_6289_), .B(_6290_), .C(_6482_), .Y(_6483_) );
NOR2X1 NOR2X1_1129 ( .gnd(gnd), .vdd(vdd), .A(_6482_), .B(_6294__bF_buf4), .Y(_6484_) );
INVX2 INVX2_228 ( .gnd(gnd), .vdd(vdd), .A(_6484_), .Y(_6485_) );
NAND2X1 NAND2X1_856 ( .gnd(gnd), .vdd(vdd), .A(_6483_), .B(_6485_), .Y(_6486_) );
NOR2X1 NOR2X1_1130 ( .gnd(gnd), .vdd(vdd), .A(_6156_), .B(_6486_), .Y(_6487_) );
AOI21X1 AOI21X1_1147 ( .gnd(gnd), .vdd(vdd), .A(_6483_), .B(_6485_), .C(_6155_), .Y(_6488_) );
OAI21X1 OAI21X1_1804 ( .gnd(gnd), .vdd(vdd), .A(_6487_), .B(_6488_), .C(micro_hash_ucr_2_pipe66_bF_buf3), .Y(_6489_) );
NAND3X1 NAND3X1_304 ( .gnd(gnd), .vdd(vdd), .A(_5075__bF_buf0), .B(_6489_), .C(_6481_), .Y(_6490_) );
INVX2 INVX2_229 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_241_), .Y(_6491_) );
XNOR2X1 XNOR2X1_231 ( .gnd(gnd), .vdd(vdd), .A(_6293__bF_buf0), .B(_6491_), .Y(_6492_) );
XOR2X1 XOR2X1_97 ( .gnd(gnd), .vdd(vdd), .A(_6492_), .B(_6279_), .Y(_6493_) );
AOI21X1 AOI21X1_1148 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe68), .B(_6493_), .C(micro_hash_ucr_2_pipe69), .Y(_6494_) );
NOR2X1 NOR2X1_1131 ( .gnd(gnd), .vdd(vdd), .A(_6282_), .B(_6154__bF_buf1), .Y(_6495_) );
INVX2 INVX2_230 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_249_), .Y(_6496_) );
OAI21X1 OAI21X1_1805 ( .gnd(gnd), .vdd(vdd), .A(_6289_), .B(_6290_), .C(_6496_), .Y(_6497_) );
INVX1 INVX1_404 ( .gnd(gnd), .vdd(vdd), .A(_6497_), .Y(_6498_) );
NOR2X1 NOR2X1_1132 ( .gnd(gnd), .vdd(vdd), .A(_6496_), .B(_6294__bF_buf3), .Y(_6499_) );
NOR2X1 NOR2X1_1133 ( .gnd(gnd), .vdd(vdd), .A(_6498_), .B(_6499_), .Y(_6500_) );
AOI21X1 AOI21X1_1149 ( .gnd(gnd), .vdd(vdd), .A(_6495_), .B(_6500_), .C(_4594__bF_buf0), .Y(_6501_) );
OAI21X1 OAI21X1_1806 ( .gnd(gnd), .vdd(vdd), .A(_6495_), .B(_6500_), .C(_6501_), .Y(_6502_) );
AOI22X1 AOI22X1_52 ( .gnd(gnd), .vdd(vdd), .A(_6147_), .B(_6502_), .C(_6490_), .D(_6494_), .Y(_4493__1_) );
OAI21X1 OAI21X1_1807 ( .gnd(gnd), .vdd(vdd), .A(_6476_), .B(_6294__bF_buf2), .C(_6479_), .Y(_6503_) );
INVX2 INVX2_231 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_226_), .Y(_6504_) );
INVX2 INVX2_232 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_k_2_), .Y(_6505_) );
INVX2 INVX2_233 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_x_2_), .Y(_6506_) );
NAND2X1 NAND2X1_857 ( .gnd(gnd), .vdd(vdd), .A(_6505_), .B(_6506_), .Y(_6507_) );
NOR2X1 NOR2X1_1134 ( .gnd(gnd), .vdd(vdd), .A(_6505_), .B(_6506_), .Y(_6508_) );
INVX1 INVX1_405 ( .gnd(gnd), .vdd(vdd), .A(_6508_), .Y(_6509_) );
AND2X2 AND2X2_452 ( .gnd(gnd), .vdd(vdd), .A(_6509_), .B(_6507_), .Y(_6510_) );
OAI21X1 OAI21X1_1808 ( .gnd(gnd), .vdd(vdd), .A(_6289_), .B(_6287_), .C(_6510_), .Y(_6511_) );
INVX8 INVX8_187 ( .gnd(gnd), .vdd(vdd), .A(_6511_), .Y(_6512_) );
OR2X2 OR2X2_52 ( .gnd(gnd), .vdd(vdd), .A(_6289_), .B(_6287_), .Y(_6513_) );
NOR2X1 NOR2X1_1135 ( .gnd(gnd), .vdd(vdd), .A(_6510_), .B(_6513_), .Y(_6514_) );
OAI21X1 OAI21X1_1809 ( .gnd(gnd), .vdd(vdd), .A(_6514__bF_buf3), .B(_6512__bF_buf3), .C(_6504_), .Y(_6515_) );
NOR2X1 NOR2X1_1136 ( .gnd(gnd), .vdd(vdd), .A(_6512__bF_buf2), .B(_6514__bF_buf2), .Y(_6516_) );
INVX8 INVX8_188 ( .gnd(gnd), .vdd(vdd), .A(_6516_), .Y(_6517_) );
NOR2X1 NOR2X1_1137 ( .gnd(gnd), .vdd(vdd), .A(_6504_), .B(_6517__bF_buf5), .Y(_6518_) );
INVX1 INVX1_406 ( .gnd(gnd), .vdd(vdd), .A(_6518_), .Y(_6519_) );
NAND2X1 NAND2X1_858 ( .gnd(gnd), .vdd(vdd), .A(_6515_), .B(_6519_), .Y(_6520_) );
XOR2X1 XOR2X1_98 ( .gnd(gnd), .vdd(vdd), .A(_6520_), .B(_6503_), .Y(_6521_) );
OR2X2 OR2X2_53 ( .gnd(gnd), .vdd(vdd), .A(_6304_), .B(_6302_), .Y(_6522_) );
NOR2X1 NOR2X1_1138 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_2_), .B(_6516_), .Y(_6523_) );
AND2X2 AND2X2_453 ( .gnd(gnd), .vdd(vdd), .A(_6516_), .B(micro_hash_ucr_2_Wx_2_), .Y(_6524_) );
NOR2X1 NOR2X1_1139 ( .gnd(gnd), .vdd(vdd), .A(_6523_), .B(_6524_), .Y(_6525_) );
AND2X2 AND2X2_454 ( .gnd(gnd), .vdd(vdd), .A(_6522_), .B(_6525_), .Y(_6526_) );
NOR2X1 NOR2X1_1140 ( .gnd(gnd), .vdd(vdd), .A(_6525_), .B(_6522_), .Y(_6527_) );
OAI21X1 OAI21X1_1810 ( .gnd(gnd), .vdd(vdd), .A(_6526_), .B(_6527_), .C(micro_hash_ucr_2_pipe8), .Y(_6528_) );
AOI21X1 AOI21X1_1150 ( .gnd(gnd), .vdd(vdd), .A(_6167_), .B(_6291_), .C(_6295_), .Y(_6529_) );
XNOR2X1 XNOR2X1_232 ( .gnd(gnd), .vdd(vdd), .A(_6516_), .B(micro_hash_ucr_2_Wx_10_), .Y(_6530_) );
XOR2X1 XOR2X1_99 ( .gnd(gnd), .vdd(vdd), .A(_6530_), .B(_6529_), .Y(_6531_) );
NAND2X1 NAND2X1_859 ( .gnd(gnd), .vdd(vdd), .A(_5372_), .B(_5134_), .Y(_6532_) );
OAI21X1 OAI21X1_1811 ( .gnd(gnd), .vdd(vdd), .A(H_2_18_), .B(_5134_), .C(_6532_), .Y(_6533_) );
AOI21X1 AOI21X1_1151 ( .gnd(gnd), .vdd(vdd), .A(_5135_), .B(_6533_), .C(micro_hash_ucr_2_pipe10), .Y(_6534_) );
AOI22X1 AOI22X1_53 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe10), .B(_6531_), .C(_6528_), .D(_6534_), .Y(_6535_) );
OAI21X1 OAI21X1_1812 ( .gnd(gnd), .vdd(vdd), .A(_6310_), .B(_6309_), .C(_6312_), .Y(_6536_) );
INVX1 INVX1_407 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_18_), .Y(_6537_) );
OAI21X1 OAI21X1_1813 ( .gnd(gnd), .vdd(vdd), .A(_6514__bF_buf1), .B(_6512__bF_buf1), .C(_6537_), .Y(_6538_) );
INVX1 INVX1_408 ( .gnd(gnd), .vdd(vdd), .A(_6538_), .Y(_6539_) );
NOR2X1 NOR2X1_1141 ( .gnd(gnd), .vdd(vdd), .A(_6537_), .B(_6517__bF_buf4), .Y(_6540_) );
NOR2X1 NOR2X1_1142 ( .gnd(gnd), .vdd(vdd), .A(_6539_), .B(_6540_), .Y(_6541_) );
XOR2X1 XOR2X1_100 ( .gnd(gnd), .vdd(vdd), .A(_6541_), .B(_6536_), .Y(_6542_) );
AOI21X1 AOI21X1_1152 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe12_bF_buf0), .B(_6542_), .C(micro_hash_ucr_2_pipe14_bF_buf2), .Y(_6543_) );
OAI21X1 OAI21X1_1814 ( .gnd(gnd), .vdd(vdd), .A(_6535_), .B(micro_hash_ucr_2_pipe12_bF_buf3), .C(_6543_), .Y(_6544_) );
AOI21X1 AOI21X1_1153 ( .gnd(gnd), .vdd(vdd), .A(_6182_), .B(_6319_), .C(_6321_), .Y(_6545_) );
INVX1 INVX1_409 ( .gnd(gnd), .vdd(vdd), .A(_6545_), .Y(_6546_) );
INVX2 INVX2_234 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_26_), .Y(_6547_) );
XNOR2X1 XNOR2X1_233 ( .gnd(gnd), .vdd(vdd), .A(_6516_), .B(_6547_), .Y(_6548_) );
NAND2X1 NAND2X1_860 ( .gnd(gnd), .vdd(vdd), .A(_6546_), .B(_6548_), .Y(_6549_) );
INVX1 INVX1_410 ( .gnd(gnd), .vdd(vdd), .A(_6549_), .Y(_6550_) );
NOR2X1 NOR2X1_1143 ( .gnd(gnd), .vdd(vdd), .A(_6546_), .B(_6548_), .Y(_6551_) );
OAI21X1 OAI21X1_1815 ( .gnd(gnd), .vdd(vdd), .A(_6550_), .B(_6551_), .C(micro_hash_ucr_2_pipe14_bF_buf1), .Y(_6552_) );
AOI21X1 AOI21X1_1154 ( .gnd(gnd), .vdd(vdd), .A(_6552_), .B(_6544_), .C(micro_hash_ucr_2_pipe16_bF_buf2), .Y(_6553_) );
OAI21X1 OAI21X1_1816 ( .gnd(gnd), .vdd(vdd), .A(_6326_), .B(_6164_), .C(_6328_), .Y(_6554_) );
INVX1 INVX1_411 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_34_), .Y(_6555_) );
OAI21X1 OAI21X1_1817 ( .gnd(gnd), .vdd(vdd), .A(_6514__bF_buf0), .B(_6512__bF_buf0), .C(_6555_), .Y(_6556_) );
NOR2X1 NOR2X1_1144 ( .gnd(gnd), .vdd(vdd), .A(_6555_), .B(_6517__bF_buf3), .Y(_6557_) );
INVX1 INVX1_412 ( .gnd(gnd), .vdd(vdd), .A(_6557_), .Y(_6558_) );
NAND2X1 NAND2X1_861 ( .gnd(gnd), .vdd(vdd), .A(_6556_), .B(_6558_), .Y(_6559_) );
XNOR2X1 XNOR2X1_234 ( .gnd(gnd), .vdd(vdd), .A(_6559_), .B(_6554_), .Y(_6560_) );
OAI21X1 OAI21X1_1818 ( .gnd(gnd), .vdd(vdd), .A(_6560_), .B(_5127__bF_buf0), .C(_5122__bF_buf2), .Y(_6561_) );
NOR2X1 NOR2X1_1145 ( .gnd(gnd), .vdd(vdd), .A(_6561_), .B(_6553_), .Y(_6562_) );
AOI21X1 AOI21X1_1155 ( .gnd(gnd), .vdd(vdd), .A(_6188_), .B(_6336_), .C(_6338_), .Y(_6563_) );
INVX2 INVX2_235 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_42_), .Y(_6564_) );
OAI21X1 OAI21X1_1819 ( .gnd(gnd), .vdd(vdd), .A(_6514__bF_buf3), .B(_6512__bF_buf3), .C(_6564_), .Y(_6565_) );
INVX1 INVX1_413 ( .gnd(gnd), .vdd(vdd), .A(_6565_), .Y(_6566_) );
NOR2X1 NOR2X1_1146 ( .gnd(gnd), .vdd(vdd), .A(_6564_), .B(_6517__bF_buf2), .Y(_6567_) );
OAI21X1 OAI21X1_1820 ( .gnd(gnd), .vdd(vdd), .A(_6567_), .B(_6566_), .C(_6563_), .Y(_6568_) );
INVX1 INVX1_414 ( .gnd(gnd), .vdd(vdd), .A(_6563_), .Y(_6569_) );
NOR2X1 NOR2X1_1147 ( .gnd(gnd), .vdd(vdd), .A(_6566_), .B(_6567_), .Y(_6570_) );
NAND2X1 NAND2X1_862 ( .gnd(gnd), .vdd(vdd), .A(_6569_), .B(_6570_), .Y(_6571_) );
NAND2X1 NAND2X1_863 ( .gnd(gnd), .vdd(vdd), .A(_6568_), .B(_6571_), .Y(_6572_) );
OAI21X1 OAI21X1_1821 ( .gnd(gnd), .vdd(vdd), .A(_6572_), .B(_5122__bF_buf1), .C(_5123__bF_buf1), .Y(_6573_) );
OAI21X1 OAI21X1_1822 ( .gnd(gnd), .vdd(vdd), .A(_6342_), .B(_6294__bF_buf1), .C(_6344_), .Y(_6574_) );
INVX2 INVX2_236 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_50_), .Y(_6575_) );
OAI21X1 OAI21X1_1823 ( .gnd(gnd), .vdd(vdd), .A(_6514__bF_buf2), .B(_6512__bF_buf2), .C(_6575_), .Y(_6576_) );
NOR2X1 NOR2X1_1148 ( .gnd(gnd), .vdd(vdd), .A(_6575_), .B(_6517__bF_buf1), .Y(_6577_) );
INVX1 INVX1_415 ( .gnd(gnd), .vdd(vdd), .A(_6577_), .Y(_6578_) );
NAND2X1 NAND2X1_864 ( .gnd(gnd), .vdd(vdd), .A(_6576_), .B(_6578_), .Y(_6579_) );
XOR2X1 XOR2X1_101 ( .gnd(gnd), .vdd(vdd), .A(_6579_), .B(_6574_), .Y(_6580_) );
AOI21X1 AOI21X1_1156 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe20_bF_buf1), .B(_6580_), .C(micro_hash_ucr_2_pipe22_bF_buf0), .Y(_6581_) );
OAI21X1 OAI21X1_1824 ( .gnd(gnd), .vdd(vdd), .A(_6562_), .B(_6573_), .C(_6581_), .Y(_6582_) );
XNOR2X1 XNOR2X1_235 ( .gnd(gnd), .vdd(vdd), .A(_6516_), .B(_5010_), .Y(_6583_) );
OAI21X1 OAI21X1_1825 ( .gnd(gnd), .vdd(vdd), .A(_6354_), .B(_6351_), .C(_6583_), .Y(_6584_) );
INVX1 INVX1_416 ( .gnd(gnd), .vdd(vdd), .A(_6584_), .Y(_6585_) );
OAI21X1 OAI21X1_1826 ( .gnd(gnd), .vdd(vdd), .A(_6353_), .B(_6349_), .C(_6352_), .Y(_6586_) );
OAI21X1 OAI21X1_1827 ( .gnd(gnd), .vdd(vdd), .A(_6586_), .B(_6583_), .C(micro_hash_ucr_2_pipe22_bF_buf4), .Y(_6587_) );
OAI21X1 OAI21X1_1828 ( .gnd(gnd), .vdd(vdd), .A(_6585_), .B(_6587_), .C(_6582_), .Y(_6588_) );
OAI21X1 OAI21X1_1829 ( .gnd(gnd), .vdd(vdd), .A(_5053_), .B(_6294__bF_buf0), .C(_6360_), .Y(_6589_) );
XNOR2X1 XNOR2X1_236 ( .gnd(gnd), .vdd(vdd), .A(_6516_), .B(_5056_), .Y(_6590_) );
NAND2X1 NAND2X1_865 ( .gnd(gnd), .vdd(vdd), .A(_6590_), .B(_6589_), .Y(_6591_) );
INVX1 INVX1_417 ( .gnd(gnd), .vdd(vdd), .A(_6591_), .Y(_6592_) );
NOR2X1 NOR2X1_1149 ( .gnd(gnd), .vdd(vdd), .A(_6590_), .B(_6589_), .Y(_6593_) );
OAI21X1 OAI21X1_1830 ( .gnd(gnd), .vdd(vdd), .A(_6592_), .B(_6593_), .C(micro_hash_ucr_2_pipe24_bF_buf2), .Y(_6594_) );
OAI21X1 OAI21X1_1831 ( .gnd(gnd), .vdd(vdd), .A(_6588_), .B(micro_hash_ucr_2_pipe24_bF_buf1), .C(_6594_), .Y(_6595_) );
AOI21X1 AOI21X1_1157 ( .gnd(gnd), .vdd(vdd), .A(_6159_), .B(_6364_), .C(_6366_), .Y(_6596_) );
OAI21X1 OAI21X1_1832 ( .gnd(gnd), .vdd(vdd), .A(_6514__bF_buf1), .B(_6512__bF_buf1), .C(_5032_), .Y(_6597_) );
INVX1 INVX1_418 ( .gnd(gnd), .vdd(vdd), .A(_6597_), .Y(_6598_) );
NOR2X1 NOR2X1_1150 ( .gnd(gnd), .vdd(vdd), .A(_5032_), .B(_6517__bF_buf0), .Y(_6599_) );
OAI21X1 OAI21X1_1833 ( .gnd(gnd), .vdd(vdd), .A(_6599_), .B(_6598_), .C(_6596_), .Y(_6600_) );
INVX1 INVX1_419 ( .gnd(gnd), .vdd(vdd), .A(_6596_), .Y(_6601_) );
NOR2X1 NOR2X1_1151 ( .gnd(gnd), .vdd(vdd), .A(_6598_), .B(_6599_), .Y(_6602_) );
NAND2X1 NAND2X1_866 ( .gnd(gnd), .vdd(vdd), .A(_6601_), .B(_6602_), .Y(_6603_) );
AOI21X1 AOI21X1_1158 ( .gnd(gnd), .vdd(vdd), .A(_6600_), .B(_6603_), .C(_5117__bF_buf3), .Y(_6604_) );
AOI21X1 AOI21X1_1159 ( .gnd(gnd), .vdd(vdd), .A(_5117__bF_buf2), .B(_6595_), .C(_6604_), .Y(_6605_) );
NAND2X1 NAND2X1_867 ( .gnd(gnd), .vdd(vdd), .A(_6205_), .B(_6370_), .Y(_6606_) );
OAI21X1 OAI21X1_1834 ( .gnd(gnd), .vdd(vdd), .A(_4938_), .B(_6294__bF_buf4), .C(_6606_), .Y(_6607_) );
OAI21X1 OAI21X1_1835 ( .gnd(gnd), .vdd(vdd), .A(_6514__bF_buf0), .B(_6512__bF_buf0), .C(_4941_), .Y(_6608_) );
NOR2X1 NOR2X1_1152 ( .gnd(gnd), .vdd(vdd), .A(_4941_), .B(_6517__bF_buf5), .Y(_6609_) );
INVX1 INVX1_420 ( .gnd(gnd), .vdd(vdd), .A(_6609_), .Y(_6610_) );
NAND2X1 NAND2X1_868 ( .gnd(gnd), .vdd(vdd), .A(_6608_), .B(_6610_), .Y(_6611_) );
XOR2X1 XOR2X1_102 ( .gnd(gnd), .vdd(vdd), .A(_6611_), .B(_6607_), .Y(_6612_) );
AOI21X1 AOI21X1_1160 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe28_bF_buf0), .B(_6612_), .C(micro_hash_ucr_2_pipe30_bF_buf1), .Y(_6613_) );
OAI21X1 OAI21X1_1836 ( .gnd(gnd), .vdd(vdd), .A(_6605_), .B(micro_hash_ucr_2_pipe28_bF_buf3), .C(_6613_), .Y(_6614_) );
XNOR2X1 XNOR2X1_237 ( .gnd(gnd), .vdd(vdd), .A(_6516_), .B(_4983_), .Y(_6615_) );
OAI21X1 OAI21X1_1837 ( .gnd(gnd), .vdd(vdd), .A(_6379_), .B(_6376_), .C(_6615_), .Y(_6616_) );
INVX1 INVX1_421 ( .gnd(gnd), .vdd(vdd), .A(_6616_), .Y(_6617_) );
OAI21X1 OAI21X1_1838 ( .gnd(gnd), .vdd(vdd), .A(_6378_), .B(_6374_), .C(_6377_), .Y(_6618_) );
OAI21X1 OAI21X1_1839 ( .gnd(gnd), .vdd(vdd), .A(_6618_), .B(_6615_), .C(micro_hash_ucr_2_pipe30_bF_buf0), .Y(_6619_) );
OAI21X1 OAI21X1_1840 ( .gnd(gnd), .vdd(vdd), .A(_6617_), .B(_6619_), .C(_6614_), .Y(_6620_) );
OAI21X1 OAI21X1_1841 ( .gnd(gnd), .vdd(vdd), .A(_4843_), .B(_6294__bF_buf3), .C(_6384_), .Y(_6621_) );
OAI21X1 OAI21X1_1842 ( .gnd(gnd), .vdd(vdd), .A(_6514__bF_buf3), .B(_6512__bF_buf3), .C(_4847_), .Y(_6622_) );
NOR2X1 NOR2X1_1153 ( .gnd(gnd), .vdd(vdd), .A(_4847_), .B(_6517__bF_buf4), .Y(_6623_) );
INVX1 INVX1_422 ( .gnd(gnd), .vdd(vdd), .A(_6623_), .Y(_6624_) );
NAND2X1 NAND2X1_869 ( .gnd(gnd), .vdd(vdd), .A(_6622_), .B(_6624_), .Y(_6625_) );
XNOR2X1 XNOR2X1_238 ( .gnd(gnd), .vdd(vdd), .A(_6625_), .B(_6621_), .Y(_6626_) );
MUX2X1 MUX2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_6620_), .B(_6626_), .S(_5111__bF_buf2), .Y(_6627_) );
AOI21X1 AOI21X1_1161 ( .gnd(gnd), .vdd(vdd), .A(_6218_), .B(_6388_), .C(_6390_), .Y(_6628_) );
OAI21X1 OAI21X1_1843 ( .gnd(gnd), .vdd(vdd), .A(_6514__bF_buf2), .B(_6512__bF_buf2), .C(_4875_), .Y(_6629_) );
INVX1 INVX1_423 ( .gnd(gnd), .vdd(vdd), .A(_6629_), .Y(_6630_) );
NOR2X1 NOR2X1_1154 ( .gnd(gnd), .vdd(vdd), .A(_4875_), .B(_6517__bF_buf3), .Y(_6631_) );
OAI21X1 OAI21X1_1844 ( .gnd(gnd), .vdd(vdd), .A(_6631_), .B(_6630_), .C(_6628_), .Y(_6632_) );
INVX1 INVX1_424 ( .gnd(gnd), .vdd(vdd), .A(_6628_), .Y(_6633_) );
NOR2X1 NOR2X1_1155 ( .gnd(gnd), .vdd(vdd), .A(_6630_), .B(_6631_), .Y(_6634_) );
NAND2X1 NAND2X1_870 ( .gnd(gnd), .vdd(vdd), .A(_6633_), .B(_6634_), .Y(_6635_) );
AOI21X1 AOI21X1_1162 ( .gnd(gnd), .vdd(vdd), .A(_6632_), .B(_6635_), .C(_5109__bF_buf1), .Y(_6636_) );
AOI21X1 AOI21X1_1163 ( .gnd(gnd), .vdd(vdd), .A(_5109__bF_buf0), .B(_6627_), .C(_6636_), .Y(_6637_) );
OAI21X1 OAI21X1_1845 ( .gnd(gnd), .vdd(vdd), .A(_4916_), .B(_6294__bF_buf2), .C(_6398_), .Y(_6638_) );
OAI21X1 OAI21X1_1846 ( .gnd(gnd), .vdd(vdd), .A(_6514__bF_buf1), .B(_6512__bF_buf1), .C(_4919_), .Y(_6639_) );
NOR2X1 NOR2X1_1156 ( .gnd(gnd), .vdd(vdd), .A(_4919_), .B(_6517__bF_buf2), .Y(_6640_) );
INVX1 INVX1_425 ( .gnd(gnd), .vdd(vdd), .A(_6640_), .Y(_6641_) );
NAND2X1 NAND2X1_871 ( .gnd(gnd), .vdd(vdd), .A(_6639_), .B(_6641_), .Y(_6642_) );
XOR2X1 XOR2X1_103 ( .gnd(gnd), .vdd(vdd), .A(_6642_), .B(_6638_), .Y(_6643_) );
AOI21X1 AOI21X1_1164 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe36_bF_buf3), .B(_6643_), .C(micro_hash_ucr_2_pipe38_bF_buf0), .Y(_6644_) );
OAI21X1 OAI21X1_1847 ( .gnd(gnd), .vdd(vdd), .A(_6637_), .B(micro_hash_ucr_2_pipe36_bF_buf2), .C(_6644_), .Y(_6645_) );
AOI21X1 AOI21X1_1165 ( .gnd(gnd), .vdd(vdd), .A(_6224_), .B(_6401_), .C(_6403_), .Y(_6646_) );
OAI21X1 OAI21X1_1848 ( .gnd(gnd), .vdd(vdd), .A(_6514__bF_buf0), .B(_6512__bF_buf0), .C(_4898_), .Y(_6647_) );
INVX1 INVX1_426 ( .gnd(gnd), .vdd(vdd), .A(_6647_), .Y(_6648_) );
NOR2X1 NOR2X1_1157 ( .gnd(gnd), .vdd(vdd), .A(_4898_), .B(_6517__bF_buf1), .Y(_6649_) );
NOR2X1 NOR2X1_1158 ( .gnd(gnd), .vdd(vdd), .A(_6648_), .B(_6649_), .Y(_6650_) );
INVX1 INVX1_427 ( .gnd(gnd), .vdd(vdd), .A(_6650_), .Y(_6651_) );
NOR2X1 NOR2X1_1159 ( .gnd(gnd), .vdd(vdd), .A(_6646_), .B(_6651_), .Y(_6652_) );
INVX1 INVX1_428 ( .gnd(gnd), .vdd(vdd), .A(_6652_), .Y(_6653_) );
OAI21X1 OAI21X1_1849 ( .gnd(gnd), .vdd(vdd), .A(_6649_), .B(_6648_), .C(_6646_), .Y(_6654_) );
NAND2X1 NAND2X1_872 ( .gnd(gnd), .vdd(vdd), .A(_6654_), .B(_6653_), .Y(_6655_) );
OAI21X1 OAI21X1_1850 ( .gnd(gnd), .vdd(vdd), .A(_5105__bF_buf3), .B(_6655_), .C(_6645_), .Y(_6656_) );
NOR2X1 NOR2X1_1160 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe40_bF_buf4), .B(_6656_), .Y(_6657_) );
NAND2X1 NAND2X1_873 ( .gnd(gnd), .vdd(vdd), .A(_6228_), .B(_6407_), .Y(_6658_) );
OAI21X1 OAI21X1_1851 ( .gnd(gnd), .vdd(vdd), .A(_4785_), .B(_6294__bF_buf1), .C(_6658_), .Y(_6659_) );
OAI21X1 OAI21X1_1852 ( .gnd(gnd), .vdd(vdd), .A(_6514__bF_buf3), .B(_6512__bF_buf3), .C(_4789_), .Y(_6660_) );
NOR2X1 NOR2X1_1161 ( .gnd(gnd), .vdd(vdd), .A(_4789_), .B(_6517__bF_buf0), .Y(_6661_) );
INVX1 INVX1_429 ( .gnd(gnd), .vdd(vdd), .A(_6661_), .Y(_6662_) );
NAND2X1 NAND2X1_874 ( .gnd(gnd), .vdd(vdd), .A(_6660_), .B(_6662_), .Y(_6663_) );
XNOR2X1 XNOR2X1_239 ( .gnd(gnd), .vdd(vdd), .A(_6663_), .B(_6659_), .Y(_6664_) );
OAI21X1 OAI21X1_1853 ( .gnd(gnd), .vdd(vdd), .A(_6664_), .B(_5103__bF_buf0), .C(_5098__bF_buf1), .Y(_6665_) );
NOR2X1 NOR2X1_1162 ( .gnd(gnd), .vdd(vdd), .A(_4980_), .B(_6294__bF_buf0), .Y(_6666_) );
OAI21X1 OAI21X1_1854 ( .gnd(gnd), .vdd(vdd), .A(_6514__bF_buf2), .B(_6512__bF_buf2), .C(_4984_), .Y(_6667_) );
INVX1 INVX1_430 ( .gnd(gnd), .vdd(vdd), .A(_6667_), .Y(_6668_) );
NOR2X1 NOR2X1_1163 ( .gnd(gnd), .vdd(vdd), .A(_4984_), .B(_6517__bF_buf5), .Y(_6669_) );
NOR2X1 NOR2X1_1164 ( .gnd(gnd), .vdd(vdd), .A(_6668_), .B(_6669_), .Y(_6670_) );
OAI21X1 OAI21X1_1855 ( .gnd(gnd), .vdd(vdd), .A(_6666_), .B(_6412_), .C(_6670_), .Y(_6671_) );
NOR2X1 NOR2X1_1165 ( .gnd(gnd), .vdd(vdd), .A(_6666_), .B(_6412_), .Y(_6672_) );
OAI21X1 OAI21X1_1856 ( .gnd(gnd), .vdd(vdd), .A(_6669_), .B(_6668_), .C(_6672_), .Y(_6673_) );
NAND2X1 NAND2X1_875 ( .gnd(gnd), .vdd(vdd), .A(_6673_), .B(_6671_), .Y(_6674_) );
OAI22X1 OAI22X1_97 ( .gnd(gnd), .vdd(vdd), .A(_5098__bF_buf0), .B(_6674_), .C(_6657_), .D(_6665_), .Y(_6675_) );
OAI21X1 OAI21X1_1857 ( .gnd(gnd), .vdd(vdd), .A(_4815_), .B(_6294__bF_buf4), .C(_6417_), .Y(_6676_) );
XNOR2X1 XNOR2X1_240 ( .gnd(gnd), .vdd(vdd), .A(_6516_), .B(_4819_), .Y(_6677_) );
NOR2X1 NOR2X1_1166 ( .gnd(gnd), .vdd(vdd), .A(_6676_), .B(_6677_), .Y(_6678_) );
NOR2X1 NOR2X1_1167 ( .gnd(gnd), .vdd(vdd), .A(_4815_), .B(_6294__bF_buf3), .Y(_6679_) );
OAI21X1 OAI21X1_1858 ( .gnd(gnd), .vdd(vdd), .A(_6418_), .B(_6679_), .C(_6677_), .Y(_6680_) );
INVX1 INVX1_431 ( .gnd(gnd), .vdd(vdd), .A(_6680_), .Y(_6681_) );
OAI21X1 OAI21X1_1859 ( .gnd(gnd), .vdd(vdd), .A(_6681_), .B(_6678_), .C(micro_hash_ucr_2_pipe44_bF_buf2), .Y(_6682_) );
OAI21X1 OAI21X1_1860 ( .gnd(gnd), .vdd(vdd), .A(_6675_), .B(micro_hash_ucr_2_pipe44_bF_buf1), .C(_6682_), .Y(_6683_) );
NAND2X1 NAND2X1_876 ( .gnd(gnd), .vdd(vdd), .A(_6239_), .B(_6421_), .Y(_6684_) );
OAI21X1 OAI21X1_1861 ( .gnd(gnd), .vdd(vdd), .A(_4701_), .B(_6294__bF_buf2), .C(_6684_), .Y(_6685_) );
OAI21X1 OAI21X1_1862 ( .gnd(gnd), .vdd(vdd), .A(_6514__bF_buf1), .B(_6512__bF_buf1), .C(_4705_), .Y(_6686_) );
NOR2X1 NOR2X1_1168 ( .gnd(gnd), .vdd(vdd), .A(_4705_), .B(_6517__bF_buf4), .Y(_6687_) );
INVX1 INVX1_432 ( .gnd(gnd), .vdd(vdd), .A(_6687_), .Y(_6688_) );
NAND2X1 NAND2X1_877 ( .gnd(gnd), .vdd(vdd), .A(_6686_), .B(_6688_), .Y(_6689_) );
XNOR2X1 XNOR2X1_241 ( .gnd(gnd), .vdd(vdd), .A(_6689_), .B(_6685_), .Y(_6690_) );
OAI21X1 OAI21X1_1863 ( .gnd(gnd), .vdd(vdd), .A(_6690_), .B(_5097__bF_buf0), .C(_5092__bF_buf4), .Y(_6691_) );
AOI21X1 AOI21X1_1166 ( .gnd(gnd), .vdd(vdd), .A(_5097__bF_buf3), .B(_6683_), .C(_6691_), .Y(_6692_) );
OAI21X1 OAI21X1_1864 ( .gnd(gnd), .vdd(vdd), .A(_4757_), .B(_6294__bF_buf1), .C(_6429_), .Y(_6693_) );
XNOR2X1 XNOR2X1_242 ( .gnd(gnd), .vdd(vdd), .A(_6516_), .B(_4760_), .Y(_6694_) );
NAND2X1 NAND2X1_878 ( .gnd(gnd), .vdd(vdd), .A(_6694_), .B(_6693_), .Y(_6695_) );
INVX1 INVX1_433 ( .gnd(gnd), .vdd(vdd), .A(_6695_), .Y(_6696_) );
OAI21X1 OAI21X1_1865 ( .gnd(gnd), .vdd(vdd), .A(_6693_), .B(_6694_), .C(micro_hash_ucr_2_pipe48_bF_buf2), .Y(_6697_) );
OAI21X1 OAI21X1_1866 ( .gnd(gnd), .vdd(vdd), .A(_6696_), .B(_6697_), .C(_5093__bF_buf4), .Y(_6698_) );
OAI21X1 OAI21X1_1867 ( .gnd(gnd), .vdd(vdd), .A(_6436_), .B(_6433_), .C(_6435_), .Y(_6699_) );
OAI21X1 OAI21X1_1868 ( .gnd(gnd), .vdd(vdd), .A(_6514__bF_buf0), .B(_6512__bF_buf0), .C(_4732_), .Y(_6700_) );
NOR2X1 NOR2X1_1169 ( .gnd(gnd), .vdd(vdd), .A(_4732_), .B(_6517__bF_buf3), .Y(_6701_) );
INVX1 INVX1_434 ( .gnd(gnd), .vdd(vdd), .A(_6701_), .Y(_6702_) );
NAND2X1 NAND2X1_879 ( .gnd(gnd), .vdd(vdd), .A(_6700_), .B(_6702_), .Y(_6703_) );
XOR2X1 XOR2X1_104 ( .gnd(gnd), .vdd(vdd), .A(_6703_), .B(_6699_), .Y(_6704_) );
AOI21X1 AOI21X1_1167 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe50_bF_buf3), .B(_6704_), .C(micro_hash_ucr_2_pipe52_bF_buf0), .Y(_6705_) );
OAI21X1 OAI21X1_1869 ( .gnd(gnd), .vdd(vdd), .A(_6692_), .B(_6698_), .C(_6705_), .Y(_6706_) );
NAND2X1 NAND2X1_880 ( .gnd(gnd), .vdd(vdd), .A(_6249_), .B(_6439_), .Y(_6707_) );
OAI21X1 OAI21X1_1870 ( .gnd(gnd), .vdd(vdd), .A(_4786_), .B(_6294__bF_buf0), .C(_6707_), .Y(_6708_) );
XNOR2X1 XNOR2X1_243 ( .gnd(gnd), .vdd(vdd), .A(_6516_), .B(_4790_), .Y(_6709_) );
NAND2X1 NAND2X1_881 ( .gnd(gnd), .vdd(vdd), .A(_6708_), .B(_6709_), .Y(_6710_) );
INVX1 INVX1_435 ( .gnd(gnd), .vdd(vdd), .A(_6710_), .Y(_6711_) );
OAI21X1 OAI21X1_1871 ( .gnd(gnd), .vdd(vdd), .A(_6709_), .B(_6708_), .C(micro_hash_ucr_2_pipe52_bF_buf3), .Y(_6712_) );
OAI21X1 OAI21X1_1872 ( .gnd(gnd), .vdd(vdd), .A(_6711_), .B(_6712_), .C(_6706_), .Y(_6713_) );
NOR2X1 NOR2X1_1170 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe54_bF_buf4), .B(_6713_), .Y(_6714_) );
NAND2X1 NAND2X1_882 ( .gnd(gnd), .vdd(vdd), .A(_6254_), .B(_6443_), .Y(_6715_) );
OAI21X1 OAI21X1_1873 ( .gnd(gnd), .vdd(vdd), .A(_4844_), .B(_6294__bF_buf4), .C(_6715_), .Y(_6716_) );
OAI21X1 OAI21X1_1874 ( .gnd(gnd), .vdd(vdd), .A(_6514__bF_buf3), .B(_6512__bF_buf3), .C(_4848_), .Y(_6717_) );
NOR2X1 NOR2X1_1171 ( .gnd(gnd), .vdd(vdd), .A(_4848_), .B(_6517__bF_buf2), .Y(_6718_) );
INVX1 INVX1_436 ( .gnd(gnd), .vdd(vdd), .A(_6718_), .Y(_6719_) );
NAND2X1 NAND2X1_883 ( .gnd(gnd), .vdd(vdd), .A(_6717_), .B(_6719_), .Y(_6720_) );
XNOR2X1 XNOR2X1_244 ( .gnd(gnd), .vdd(vdd), .A(_6720_), .B(_6716_), .Y(_6721_) );
OAI21X1 OAI21X1_1875 ( .gnd(gnd), .vdd(vdd), .A(_6721_), .B(_5086__bF_buf0), .C(_5087__bF_buf4), .Y(_6722_) );
NOR2X1 NOR2X1_1172 ( .gnd(gnd), .vdd(vdd), .A(_4816_), .B(_6294__bF_buf3), .Y(_6723_) );
XNOR2X1 XNOR2X1_245 ( .gnd(gnd), .vdd(vdd), .A(_6516_), .B(_4820_), .Y(_6724_) );
OAI21X1 OAI21X1_1876 ( .gnd(gnd), .vdd(vdd), .A(_6723_), .B(_6450_), .C(_6724_), .Y(_6725_) );
INVX1 INVX1_437 ( .gnd(gnd), .vdd(vdd), .A(_6725_), .Y(_6726_) );
OAI21X1 OAI21X1_1877 ( .gnd(gnd), .vdd(vdd), .A(_4816_), .B(_6294__bF_buf2), .C(_6449_), .Y(_6727_) );
OAI21X1 OAI21X1_1878 ( .gnd(gnd), .vdd(vdd), .A(_6724_), .B(_6727_), .C(micro_hash_ucr_2_pipe56_bF_buf3), .Y(_6728_) );
OAI22X1 OAI22X1_98 ( .gnd(gnd), .vdd(vdd), .A(_6726_), .B(_6728_), .C(_6714_), .D(_6722_), .Y(_6729_) );
AOI21X1 AOI21X1_1168 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_201_), .B(_6293__bF_buf4), .C(_6455_), .Y(_6730_) );
XNOR2X1 XNOR2X1_246 ( .gnd(gnd), .vdd(vdd), .A(_6516_), .B(_4706_), .Y(_6731_) );
INVX1 INVX1_438 ( .gnd(gnd), .vdd(vdd), .A(_6731_), .Y(_6732_) );
NAND2X1 NAND2X1_884 ( .gnd(gnd), .vdd(vdd), .A(_6730_), .B(_6732_), .Y(_6733_) );
NOR2X1 NOR2X1_1173 ( .gnd(gnd), .vdd(vdd), .A(_6730_), .B(_6732_), .Y(_6734_) );
INVX1 INVX1_439 ( .gnd(gnd), .vdd(vdd), .A(_6734_), .Y(_6735_) );
NAND2X1 NAND2X1_885 ( .gnd(gnd), .vdd(vdd), .A(_6733_), .B(_6735_), .Y(_6736_) );
OAI21X1 OAI21X1_1879 ( .gnd(gnd), .vdd(vdd), .A(_6736_), .B(_5085__bF_buf0), .C(_5080__bF_buf2), .Y(_6737_) );
AOI21X1 AOI21X1_1169 ( .gnd(gnd), .vdd(vdd), .A(_5085__bF_buf3), .B(_6729_), .C(_6737_), .Y(_6738_) );
OAI21X1 OAI21X1_1880 ( .gnd(gnd), .vdd(vdd), .A(_6460_), .B(_6459_), .C(_6462_), .Y(_6739_) );
OAI21X1 OAI21X1_1881 ( .gnd(gnd), .vdd(vdd), .A(_6514__bF_buf2), .B(_6512__bF_buf2), .C(_4761_), .Y(_6740_) );
NOR2X1 NOR2X1_1174 ( .gnd(gnd), .vdd(vdd), .A(_4761_), .B(_6517__bF_buf1), .Y(_6741_) );
INVX1 INVX1_440 ( .gnd(gnd), .vdd(vdd), .A(_6741_), .Y(_6742_) );
NAND2X1 NAND2X1_886 ( .gnd(gnd), .vdd(vdd), .A(_6740_), .B(_6742_), .Y(_6743_) );
XNOR2X1 XNOR2X1_247 ( .gnd(gnd), .vdd(vdd), .A(_6743_), .B(_6739_), .Y(_6744_) );
OAI21X1 OAI21X1_1882 ( .gnd(gnd), .vdd(vdd), .A(_6744_), .B(_5080__bF_buf1), .C(_5081__bF_buf2), .Y(_6745_) );
NOR2X1 NOR2X1_1175 ( .gnd(gnd), .vdd(vdd), .A(_6745_), .B(_6738_), .Y(_6746_) );
NOR2X1 NOR2X1_1176 ( .gnd(gnd), .vdd(vdd), .A(_6470_), .B(_6472_), .Y(_6747_) );
INVX1 INVX1_441 ( .gnd(gnd), .vdd(vdd), .A(_6747_), .Y(_6748_) );
XNOR2X1 XNOR2X1_248 ( .gnd(gnd), .vdd(vdd), .A(_6516_), .B(_4733_), .Y(_6749_) );
OAI21X1 OAI21X1_1883 ( .gnd(gnd), .vdd(vdd), .A(_6748_), .B(_6749_), .C(micro_hash_ucr_2_pipe62_bF_buf1), .Y(_6750_) );
AOI21X1 AOI21X1_1170 ( .gnd(gnd), .vdd(vdd), .A(_6748_), .B(_6749_), .C(_6750_), .Y(_6751_) );
OAI21X1 OAI21X1_1884 ( .gnd(gnd), .vdd(vdd), .A(_6746_), .B(_6751_), .C(_5079__bF_buf3), .Y(_6752_) );
OAI21X1 OAI21X1_1885 ( .gnd(gnd), .vdd(vdd), .A(_5079__bF_buf2), .B(_6521_), .C(_6752_), .Y(_6753_) );
OAI21X1 OAI21X1_1886 ( .gnd(gnd), .vdd(vdd), .A(_6486_), .B(_6156_), .C(_6485_), .Y(_6754_) );
INVX2 INVX2_237 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_234_), .Y(_6755_) );
XNOR2X1 XNOR2X1_249 ( .gnd(gnd), .vdd(vdd), .A(_6516_), .B(_6755_), .Y(_6756_) );
NOR2X1 NOR2X1_1177 ( .gnd(gnd), .vdd(vdd), .A(_6756_), .B(_6754_), .Y(_6757_) );
OAI21X1 OAI21X1_1887 ( .gnd(gnd), .vdd(vdd), .A(_6487_), .B(_6484_), .C(_6756_), .Y(_6758_) );
NAND2X1 NAND2X1_887 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe66_bF_buf2), .B(_6758_), .Y(_6759_) );
OAI21X1 OAI21X1_1888 ( .gnd(gnd), .vdd(vdd), .A(_6759_), .B(_6757_), .C(_5075__bF_buf4), .Y(_6760_) );
AOI21X1 AOI21X1_1171 ( .gnd(gnd), .vdd(vdd), .A(_5074__bF_buf1), .B(_6753_), .C(_6760_), .Y(_6761_) );
NAND2X1 NAND2X1_888 ( .gnd(gnd), .vdd(vdd), .A(_6279_), .B(_6492_), .Y(_6762_) );
OAI21X1 OAI21X1_1889 ( .gnd(gnd), .vdd(vdd), .A(_6491_), .B(_6294__bF_buf1), .C(_6762_), .Y(_6763_) );
INVX2 INVX2_238 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_242_), .Y(_6764_) );
OAI21X1 OAI21X1_1890 ( .gnd(gnd), .vdd(vdd), .A(_6514__bF_buf1), .B(_6512__bF_buf1), .C(_6764_), .Y(_6765_) );
NOR2X1 NOR2X1_1178 ( .gnd(gnd), .vdd(vdd), .A(_6764_), .B(_6517__bF_buf0), .Y(_6766_) );
INVX1 INVX1_442 ( .gnd(gnd), .vdd(vdd), .A(_6766_), .Y(_6767_) );
NAND2X1 NAND2X1_889 ( .gnd(gnd), .vdd(vdd), .A(_6765_), .B(_6767_), .Y(_6768_) );
XNOR2X1 XNOR2X1_250 ( .gnd(gnd), .vdd(vdd), .A(_6768_), .B(_6763_), .Y(_6769_) );
OAI21X1 OAI21X1_1891 ( .gnd(gnd), .vdd(vdd), .A(_6769_), .B(_5075__bF_buf3), .C(_6146_), .Y(_6770_) );
NAND2X1 NAND2X1_890 ( .gnd(gnd), .vdd(vdd), .A(_6495_), .B(_6500_), .Y(_6771_) );
OAI21X1 OAI21X1_1892 ( .gnd(gnd), .vdd(vdd), .A(_6496_), .B(_6294__bF_buf0), .C(_6771_), .Y(_6772_) );
INVX1 INVX1_443 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_250_), .Y(_6773_) );
OAI21X1 OAI21X1_1893 ( .gnd(gnd), .vdd(vdd), .A(_6514__bF_buf0), .B(_6512__bF_buf0), .C(_6773_), .Y(_6774_) );
INVX1 INVX1_444 ( .gnd(gnd), .vdd(vdd), .A(_6774_), .Y(_6775_) );
NOR2X1 NOR2X1_1179 ( .gnd(gnd), .vdd(vdd), .A(_6773_), .B(_6517__bF_buf5), .Y(_6776_) );
NOR2X1 NOR2X1_1180 ( .gnd(gnd), .vdd(vdd), .A(_6775_), .B(_6776_), .Y(_6777_) );
AND2X2 AND2X2_455 ( .gnd(gnd), .vdd(vdd), .A(_6777_), .B(_6772_), .Y(_6778_) );
OAI21X1 OAI21X1_1894 ( .gnd(gnd), .vdd(vdd), .A(_6777_), .B(_6772_), .C(_4563_), .Y(_6779_) );
OAI22X1 OAI22X1_99 ( .gnd(gnd), .vdd(vdd), .A(_6778_), .B(_6779_), .C(_6761_), .D(_6770_), .Y(_4493__2_) );
NOR2X1 NOR2X1_1181 ( .gnd(gnd), .vdd(vdd), .A(_6524_), .B(_6526_), .Y(_6780_) );
INVX1 INVX1_445 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_3_), .Y(_6781_) );
OAI21X1 OAI21X1_1895 ( .gnd(gnd), .vdd(vdd), .A(_6505_), .B(_6506_), .C(_6511_), .Y(_6782_) );
XOR2X1 XOR2X1_105 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_k_3_), .B(micro_hash_ucr_2_x_3_), .Y(_6783_) );
AND2X2 AND2X2_456 ( .gnd(gnd), .vdd(vdd), .A(_6782_), .B(_6783_), .Y(_6784_) );
NOR2X1 NOR2X1_1182 ( .gnd(gnd), .vdd(vdd), .A(_6783_), .B(_6782_), .Y(_6785_) );
OAI21X1 OAI21X1_1896 ( .gnd(gnd), .vdd(vdd), .A(_6784__bF_buf4), .B(_6785__bF_buf4), .C(_6781_), .Y(_6786_) );
NOR2X1 NOR2X1_1183 ( .gnd(gnd), .vdd(vdd), .A(_6785__bF_buf3), .B(_6784__bF_buf3), .Y(_6787_) );
NAND2X1 NAND2X1_891 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_3_), .B(_6787_), .Y(_6788_) );
AND2X2 AND2X2_457 ( .gnd(gnd), .vdd(vdd), .A(_6788_), .B(_6786_), .Y(_6789_) );
OAI21X1 OAI21X1_1897 ( .gnd(gnd), .vdd(vdd), .A(_6780_), .B(_6789_), .C(micro_hash_ucr_2_pipe8), .Y(_6790_) );
AOI21X1 AOI21X1_1172 ( .gnd(gnd), .vdd(vdd), .A(_6780_), .B(_6789_), .C(_6790_), .Y(_6791_) );
NOR2X1 NOR2X1_1184 ( .gnd(gnd), .vdd(vdd), .A(_8653_), .B(_5134_), .Y(_6792_) );
OAI21X1 OAI21X1_1898 ( .gnd(gnd), .vdd(vdd), .A(_8654_), .B(micro_hash_ucr_2_pipe6), .C(_5135_), .Y(_6793_) );
OAI21X1 OAI21X1_1899 ( .gnd(gnd), .vdd(vdd), .A(_6793_), .B(_6792_), .C(_5133_), .Y(_6794_) );
NOR2X1 NOR2X1_1185 ( .gnd(gnd), .vdd(vdd), .A(_6529_), .B(_6530_), .Y(_6795_) );
AOI21X1 AOI21X1_1173 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_10_), .B(_6516_), .C(_6795_), .Y(_6796_) );
INVX1 INVX1_446 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_11_), .Y(_6797_) );
OAI21X1 OAI21X1_1900 ( .gnd(gnd), .vdd(vdd), .A(_6784__bF_buf2), .B(_6785__bF_buf2), .C(_6797_), .Y(_6798_) );
NAND2X1 NAND2X1_892 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_11_), .B(_6787_), .Y(_6799_) );
NAND2X1 NAND2X1_893 ( .gnd(gnd), .vdd(vdd), .A(_6798_), .B(_6799_), .Y(_6800_) );
XOR2X1 XOR2X1_106 ( .gnd(gnd), .vdd(vdd), .A(_6796_), .B(_6800_), .Y(_6801_) );
AOI21X1 AOI21X1_1174 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe10), .B(_6801_), .C(micro_hash_ucr_2_pipe12_bF_buf2), .Y(_6802_) );
OAI21X1 OAI21X1_1901 ( .gnd(gnd), .vdd(vdd), .A(_6791_), .B(_6794_), .C(_6802_), .Y(_6803_) );
AOI21X1 AOI21X1_1175 ( .gnd(gnd), .vdd(vdd), .A(_6536_), .B(_6538_), .C(_6540_), .Y(_6804_) );
INVX2 INVX2_239 ( .gnd(gnd), .vdd(vdd), .A(_6804_), .Y(_6805_) );
INVX1 INVX1_447 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_19_), .Y(_6806_) );
OAI21X1 OAI21X1_1902 ( .gnd(gnd), .vdd(vdd), .A(_6784__bF_buf1), .B(_6785__bF_buf1), .C(_6806_), .Y(_6807_) );
INVX8 INVX8_189 ( .gnd(gnd), .vdd(vdd), .A(_6787_), .Y(_6808_) );
NOR2X1 NOR2X1_1186 ( .gnd(gnd), .vdd(vdd), .A(_6806_), .B(_6808__bF_buf4), .Y(_6809_) );
INVX1 INVX1_448 ( .gnd(gnd), .vdd(vdd), .A(_6809_), .Y(_6810_) );
NAND2X1 NAND2X1_894 ( .gnd(gnd), .vdd(vdd), .A(_6807_), .B(_6810_), .Y(_6811_) );
AOI21X1 AOI21X1_1176 ( .gnd(gnd), .vdd(vdd), .A(_6805_), .B(_6811_), .C(_5128_), .Y(_6812_) );
OAI21X1 OAI21X1_1903 ( .gnd(gnd), .vdd(vdd), .A(_6805_), .B(_6811_), .C(_6812_), .Y(_6813_) );
AOI21X1 AOI21X1_1177 ( .gnd(gnd), .vdd(vdd), .A(_6813_), .B(_6803_), .C(micro_hash_ucr_2_pipe14_bF_buf0), .Y(_6814_) );
OAI21X1 OAI21X1_1904 ( .gnd(gnd), .vdd(vdd), .A(_6547_), .B(_6517__bF_buf4), .C(_6549_), .Y(_6815_) );
INVX1 INVX1_449 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_27_), .Y(_6816_) );
OAI21X1 OAI21X1_1905 ( .gnd(gnd), .vdd(vdd), .A(_6784__bF_buf0), .B(_6785__bF_buf0), .C(_6816_), .Y(_6817_) );
INVX1 INVX1_450 ( .gnd(gnd), .vdd(vdd), .A(_6817_), .Y(_6818_) );
NOR2X1 NOR2X1_1187 ( .gnd(gnd), .vdd(vdd), .A(_6816_), .B(_6808__bF_buf3), .Y(_6819_) );
NOR2X1 NOR2X1_1188 ( .gnd(gnd), .vdd(vdd), .A(_6818_), .B(_6819_), .Y(_6820_) );
XOR2X1 XOR2X1_107 ( .gnd(gnd), .vdd(vdd), .A(_6820_), .B(_6815_), .Y(_6821_) );
NOR2X1 NOR2X1_1189 ( .gnd(gnd), .vdd(vdd), .A(_5129_), .B(_6821_), .Y(_6822_) );
OAI21X1 OAI21X1_1906 ( .gnd(gnd), .vdd(vdd), .A(_6814_), .B(_6822_), .C(_5127__bF_buf3), .Y(_6823_) );
AOI21X1 AOI21X1_1178 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_33_), .B(_6293__bF_buf3), .C(_6330_), .Y(_6824_) );
OAI21X1 OAI21X1_1907 ( .gnd(gnd), .vdd(vdd), .A(_6559_), .B(_6824_), .C(_6558_), .Y(_6825_) );
INVX1 INVX1_451 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_35_), .Y(_6826_) );
OAI21X1 OAI21X1_1908 ( .gnd(gnd), .vdd(vdd), .A(_6784__bF_buf4), .B(_6785__bF_buf4), .C(_6826_), .Y(_6827_) );
NOR2X1 NOR2X1_1190 ( .gnd(gnd), .vdd(vdd), .A(_6826_), .B(_6808__bF_buf2), .Y(_6828_) );
INVX1 INVX1_452 ( .gnd(gnd), .vdd(vdd), .A(_6828_), .Y(_6829_) );
NAND2X1 NAND2X1_895 ( .gnd(gnd), .vdd(vdd), .A(_6827_), .B(_6829_), .Y(_6830_) );
AOI21X1 AOI21X1_1179 ( .gnd(gnd), .vdd(vdd), .A(_6830_), .B(_6825_), .C(_5127__bF_buf2), .Y(_6831_) );
OAI21X1 OAI21X1_1909 ( .gnd(gnd), .vdd(vdd), .A(_6825_), .B(_6830_), .C(_6831_), .Y(_6832_) );
AND2X2 AND2X2_458 ( .gnd(gnd), .vdd(vdd), .A(_6832_), .B(_5122__bF_buf0), .Y(_6833_) );
OAI21X1 OAI21X1_1910 ( .gnd(gnd), .vdd(vdd), .A(_6564_), .B(_6517__bF_buf3), .C(_6571_), .Y(_6834_) );
INVX1 INVX1_453 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_43_), .Y(_6835_) );
OAI21X1 OAI21X1_1911 ( .gnd(gnd), .vdd(vdd), .A(_6784__bF_buf3), .B(_6785__bF_buf3), .C(_6835_), .Y(_6836_) );
NOR2X1 NOR2X1_1191 ( .gnd(gnd), .vdd(vdd), .A(_6835_), .B(_6808__bF_buf1), .Y(_6837_) );
INVX1 INVX1_454 ( .gnd(gnd), .vdd(vdd), .A(_6837_), .Y(_6838_) );
NAND2X1 NAND2X1_896 ( .gnd(gnd), .vdd(vdd), .A(_6836_), .B(_6838_), .Y(_6839_) );
XOR2X1 XOR2X1_108 ( .gnd(gnd), .vdd(vdd), .A(_6834_), .B(_6839_), .Y(_6840_) );
OAI21X1 OAI21X1_1912 ( .gnd(gnd), .vdd(vdd), .A(_6840_), .B(_5122__bF_buf4), .C(_5123__bF_buf0), .Y(_6841_) );
AOI21X1 AOI21X1_1180 ( .gnd(gnd), .vdd(vdd), .A(_6833_), .B(_6823_), .C(_6841_), .Y(_6842_) );
NAND3X1 NAND3X1_305 ( .gnd(gnd), .vdd(vdd), .A(_6574_), .B(_6576_), .C(_6578_), .Y(_6843_) );
OAI21X1 OAI21X1_1913 ( .gnd(gnd), .vdd(vdd), .A(_6575_), .B(_6517__bF_buf2), .C(_6843_), .Y(_6844_) );
INVX1 INVX1_455 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_51_), .Y(_6845_) );
OAI21X1 OAI21X1_1914 ( .gnd(gnd), .vdd(vdd), .A(_6784__bF_buf2), .B(_6785__bF_buf2), .C(_6845_), .Y(_6846_) );
NOR2X1 NOR2X1_1192 ( .gnd(gnd), .vdd(vdd), .A(_6845_), .B(_6808__bF_buf0), .Y(_6847_) );
INVX1 INVX1_456 ( .gnd(gnd), .vdd(vdd), .A(_6847_), .Y(_6848_) );
NAND2X1 NAND2X1_897 ( .gnd(gnd), .vdd(vdd), .A(_6846_), .B(_6848_), .Y(_6849_) );
XNOR2X1 XNOR2X1_251 ( .gnd(gnd), .vdd(vdd), .A(_6844_), .B(_6849_), .Y(_6850_) );
OAI21X1 OAI21X1_1915 ( .gnd(gnd), .vdd(vdd), .A(_6850_), .B(_5123__bF_buf4), .C(_5121__bF_buf0), .Y(_6851_) );
OAI21X1 OAI21X1_1916 ( .gnd(gnd), .vdd(vdd), .A(_5010_), .B(_6517__bF_buf1), .C(_6584_), .Y(_6852_) );
OAI21X1 OAI21X1_1917 ( .gnd(gnd), .vdd(vdd), .A(_6784__bF_buf1), .B(_6785__bF_buf1), .C(_5013_), .Y(_6853_) );
INVX1 INVX1_457 ( .gnd(gnd), .vdd(vdd), .A(_6853_), .Y(_6854_) );
NOR2X1 NOR2X1_1193 ( .gnd(gnd), .vdd(vdd), .A(_5013_), .B(_6808__bF_buf4), .Y(_6855_) );
NOR2X1 NOR2X1_1194 ( .gnd(gnd), .vdd(vdd), .A(_6854_), .B(_6855_), .Y(_6856_) );
XOR2X1 XOR2X1_109 ( .gnd(gnd), .vdd(vdd), .A(_6852_), .B(_6856_), .Y(_6857_) );
AOI21X1 AOI21X1_1181 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe22_bF_buf3), .B(_6857_), .C(micro_hash_ucr_2_pipe24_bF_buf0), .Y(_6858_) );
OAI21X1 OAI21X1_1918 ( .gnd(gnd), .vdd(vdd), .A(_6842_), .B(_6851_), .C(_6858_), .Y(_6859_) );
OAI21X1 OAI21X1_1919 ( .gnd(gnd), .vdd(vdd), .A(_5056_), .B(_6517__bF_buf0), .C(_6591_), .Y(_6860_) );
OAI21X1 OAI21X1_1920 ( .gnd(gnd), .vdd(vdd), .A(_6784__bF_buf0), .B(_6785__bF_buf0), .C(_5059_), .Y(_6861_) );
NOR2X1 NOR2X1_1195 ( .gnd(gnd), .vdd(vdd), .A(_5059_), .B(_6808__bF_buf3), .Y(_6862_) );
INVX1 INVX1_458 ( .gnd(gnd), .vdd(vdd), .A(_6862_), .Y(_6863_) );
NAND2X1 NAND2X1_898 ( .gnd(gnd), .vdd(vdd), .A(_6861_), .B(_6863_), .Y(_6864_) );
AOI21X1 AOI21X1_1182 ( .gnd(gnd), .vdd(vdd), .A(_6860_), .B(_6864_), .C(_5116__bF_buf0), .Y(_6865_) );
OAI21X1 OAI21X1_1921 ( .gnd(gnd), .vdd(vdd), .A(_6860_), .B(_6864_), .C(_6865_), .Y(_6866_) );
AND2X2 AND2X2_459 ( .gnd(gnd), .vdd(vdd), .A(_6866_), .B(_5117__bF_buf1), .Y(_6867_) );
OAI21X1 OAI21X1_1922 ( .gnd(gnd), .vdd(vdd), .A(_5032_), .B(_6517__bF_buf5), .C(_6603_), .Y(_6868_) );
OAI21X1 OAI21X1_1923 ( .gnd(gnd), .vdd(vdd), .A(_6784__bF_buf4), .B(_6785__bF_buf4), .C(_5035_), .Y(_6869_) );
NOR2X1 NOR2X1_1196 ( .gnd(gnd), .vdd(vdd), .A(_5035_), .B(_6808__bF_buf2), .Y(_6870_) );
INVX1 INVX1_459 ( .gnd(gnd), .vdd(vdd), .A(_6870_), .Y(_6871_) );
NAND2X1 NAND2X1_899 ( .gnd(gnd), .vdd(vdd), .A(_6869_), .B(_6871_), .Y(_6872_) );
XOR2X1 XOR2X1_110 ( .gnd(gnd), .vdd(vdd), .A(_6868_), .B(_6872_), .Y(_6873_) );
OAI21X1 OAI21X1_1924 ( .gnd(gnd), .vdd(vdd), .A(_6873_), .B(_5117__bF_buf0), .C(_5115__bF_buf3), .Y(_6874_) );
AOI21X1 AOI21X1_1183 ( .gnd(gnd), .vdd(vdd), .A(_6867_), .B(_6859_), .C(_6874_), .Y(_6875_) );
NAND3X1 NAND3X1_306 ( .gnd(gnd), .vdd(vdd), .A(_6607_), .B(_6608_), .C(_6610_), .Y(_6876_) );
OAI21X1 OAI21X1_1925 ( .gnd(gnd), .vdd(vdd), .A(_4941_), .B(_6517__bF_buf4), .C(_6876_), .Y(_6877_) );
OAI21X1 OAI21X1_1926 ( .gnd(gnd), .vdd(vdd), .A(_6784__bF_buf3), .B(_6785__bF_buf3), .C(_4944_), .Y(_6878_) );
NOR2X1 NOR2X1_1197 ( .gnd(gnd), .vdd(vdd), .A(_4944_), .B(_6808__bF_buf1), .Y(_6879_) );
INVX1 INVX1_460 ( .gnd(gnd), .vdd(vdd), .A(_6879_), .Y(_6880_) );
NAND2X1 NAND2X1_900 ( .gnd(gnd), .vdd(vdd), .A(_6878_), .B(_6880_), .Y(_6881_) );
XNOR2X1 XNOR2X1_252 ( .gnd(gnd), .vdd(vdd), .A(_6877_), .B(_6881_), .Y(_6882_) );
OAI21X1 OAI21X1_1927 ( .gnd(gnd), .vdd(vdd), .A(_6882_), .B(_5115__bF_buf2), .C(_5110__bF_buf2), .Y(_6883_) );
OAI21X1 OAI21X1_1928 ( .gnd(gnd), .vdd(vdd), .A(_4983_), .B(_6517__bF_buf3), .C(_6616_), .Y(_6884_) );
OAI21X1 OAI21X1_1929 ( .gnd(gnd), .vdd(vdd), .A(_6784__bF_buf2), .B(_6785__bF_buf2), .C(_4987_), .Y(_6885_) );
INVX1 INVX1_461 ( .gnd(gnd), .vdd(vdd), .A(_6885_), .Y(_6886_) );
NOR2X1 NOR2X1_1198 ( .gnd(gnd), .vdd(vdd), .A(_4987_), .B(_6808__bF_buf0), .Y(_6887_) );
NOR2X1 NOR2X1_1199 ( .gnd(gnd), .vdd(vdd), .A(_6886_), .B(_6887_), .Y(_6888_) );
XOR2X1 XOR2X1_111 ( .gnd(gnd), .vdd(vdd), .A(_6884_), .B(_6888_), .Y(_6889_) );
AOI21X1 AOI21X1_1184 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe30_bF_buf4), .B(_6889_), .C(micro_hash_ucr_2_pipe32_bF_buf1), .Y(_6890_) );
OAI21X1 OAI21X1_1930 ( .gnd(gnd), .vdd(vdd), .A(_6875_), .B(_6883_), .C(_6890_), .Y(_6891_) );
NAND3X1 NAND3X1_307 ( .gnd(gnd), .vdd(vdd), .A(_6621_), .B(_6622_), .C(_6624_), .Y(_6892_) );
OAI21X1 OAI21X1_1931 ( .gnd(gnd), .vdd(vdd), .A(_4847_), .B(_6517__bF_buf2), .C(_6892_), .Y(_6893_) );
OAI21X1 OAI21X1_1932 ( .gnd(gnd), .vdd(vdd), .A(_6784__bF_buf1), .B(_6785__bF_buf1), .C(_4851_), .Y(_6894_) );
NOR2X1 NOR2X1_1200 ( .gnd(gnd), .vdd(vdd), .A(_4851_), .B(_6808__bF_buf4), .Y(_6895_) );
INVX1 INVX1_462 ( .gnd(gnd), .vdd(vdd), .A(_6895_), .Y(_6896_) );
NAND2X1 NAND2X1_901 ( .gnd(gnd), .vdd(vdd), .A(_6894_), .B(_6896_), .Y(_6897_) );
AOI21X1 AOI21X1_1185 ( .gnd(gnd), .vdd(vdd), .A(_6897_), .B(_6893_), .C(_5111__bF_buf1), .Y(_6898_) );
OAI21X1 OAI21X1_1933 ( .gnd(gnd), .vdd(vdd), .A(_6893_), .B(_6897_), .C(_6898_), .Y(_6899_) );
AND2X2 AND2X2_460 ( .gnd(gnd), .vdd(vdd), .A(_6899_), .B(_5109__bF_buf4), .Y(_6900_) );
OAI21X1 OAI21X1_1934 ( .gnd(gnd), .vdd(vdd), .A(_4875_), .B(_6517__bF_buf1), .C(_6635_), .Y(_6901_) );
OAI21X1 OAI21X1_1935 ( .gnd(gnd), .vdd(vdd), .A(_6784__bF_buf0), .B(_6785__bF_buf0), .C(_4878_), .Y(_6902_) );
NOR2X1 NOR2X1_1201 ( .gnd(gnd), .vdd(vdd), .A(_4878_), .B(_6808__bF_buf3), .Y(_6903_) );
INVX1 INVX1_463 ( .gnd(gnd), .vdd(vdd), .A(_6903_), .Y(_6904_) );
NAND2X1 NAND2X1_902 ( .gnd(gnd), .vdd(vdd), .A(_6902_), .B(_6904_), .Y(_6905_) );
XOR2X1 XOR2X1_112 ( .gnd(gnd), .vdd(vdd), .A(_6901_), .B(_6905_), .Y(_6906_) );
OAI21X1 OAI21X1_1936 ( .gnd(gnd), .vdd(vdd), .A(_6906_), .B(_5109__bF_buf3), .C(_5104__bF_buf4), .Y(_6907_) );
AOI21X1 AOI21X1_1186 ( .gnd(gnd), .vdd(vdd), .A(_6900_), .B(_6891_), .C(_6907_), .Y(_6908_) );
NAND3X1 NAND3X1_308 ( .gnd(gnd), .vdd(vdd), .A(_6638_), .B(_6639_), .C(_6641_), .Y(_6909_) );
OAI21X1 OAI21X1_1937 ( .gnd(gnd), .vdd(vdd), .A(_4919_), .B(_6517__bF_buf0), .C(_6909_), .Y(_6910_) );
XNOR2X1 XNOR2X1_253 ( .gnd(gnd), .vdd(vdd), .A(_6787_), .B(micro_hash_ucr_2_Wx_115_), .Y(_6911_) );
XNOR2X1 XNOR2X1_254 ( .gnd(gnd), .vdd(vdd), .A(_6910_), .B(_6911_), .Y(_6912_) );
OAI21X1 OAI21X1_1938 ( .gnd(gnd), .vdd(vdd), .A(_6912_), .B(_5104__bF_buf3), .C(_5105__bF_buf2), .Y(_6913_) );
OAI21X1 OAI21X1_1939 ( .gnd(gnd), .vdd(vdd), .A(_4898_), .B(_6517__bF_buf5), .C(_6653_), .Y(_6914_) );
OAI21X1 OAI21X1_1940 ( .gnd(gnd), .vdd(vdd), .A(_6784__bF_buf4), .B(_6785__bF_buf4), .C(_4901_), .Y(_6915_) );
NOR2X1 NOR2X1_1202 ( .gnd(gnd), .vdd(vdd), .A(_4901_), .B(_6808__bF_buf2), .Y(_6916_) );
INVX1 INVX1_464 ( .gnd(gnd), .vdd(vdd), .A(_6916_), .Y(_6917_) );
NAND2X1 NAND2X1_903 ( .gnd(gnd), .vdd(vdd), .A(_6915_), .B(_6917_), .Y(_6918_) );
XNOR2X1 XNOR2X1_255 ( .gnd(gnd), .vdd(vdd), .A(_6914_), .B(_6918_), .Y(_6919_) );
AOI21X1 AOI21X1_1187 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe38_bF_buf3), .B(_6919_), .C(micro_hash_ucr_2_pipe40_bF_buf3), .Y(_6920_) );
OAI21X1 OAI21X1_1941 ( .gnd(gnd), .vdd(vdd), .A(_6908_), .B(_6913_), .C(_6920_), .Y(_6921_) );
NAND3X1 NAND3X1_309 ( .gnd(gnd), .vdd(vdd), .A(_6659_), .B(_6660_), .C(_6662_), .Y(_6922_) );
OAI21X1 OAI21X1_1942 ( .gnd(gnd), .vdd(vdd), .A(_4789_), .B(_6517__bF_buf4), .C(_6922_), .Y(_6923_) );
OAI21X1 OAI21X1_1943 ( .gnd(gnd), .vdd(vdd), .A(_6784__bF_buf3), .B(_6785__bF_buf3), .C(_4793_), .Y(_6924_) );
NOR2X1 NOR2X1_1203 ( .gnd(gnd), .vdd(vdd), .A(_4793_), .B(_6808__bF_buf1), .Y(_6925_) );
INVX1 INVX1_465 ( .gnd(gnd), .vdd(vdd), .A(_6925_), .Y(_6926_) );
NAND2X1 NAND2X1_904 ( .gnd(gnd), .vdd(vdd), .A(_6924_), .B(_6926_), .Y(_6927_) );
AOI21X1 AOI21X1_1188 ( .gnd(gnd), .vdd(vdd), .A(_6927_), .B(_6923_), .C(_5103__bF_buf3), .Y(_6928_) );
OAI21X1 OAI21X1_1944 ( .gnd(gnd), .vdd(vdd), .A(_6923_), .B(_6927_), .C(_6928_), .Y(_6929_) );
AND2X2 AND2X2_461 ( .gnd(gnd), .vdd(vdd), .A(_6929_), .B(_5098__bF_buf4), .Y(_6930_) );
OAI21X1 OAI21X1_1945 ( .gnd(gnd), .vdd(vdd), .A(_4984_), .B(_6517__bF_buf3), .C(_6671_), .Y(_6931_) );
OAI21X1 OAI21X1_1946 ( .gnd(gnd), .vdd(vdd), .A(_6784__bF_buf2), .B(_6785__bF_buf2), .C(_4988_), .Y(_6932_) );
NOR2X1 NOR2X1_1204 ( .gnd(gnd), .vdd(vdd), .A(_4988_), .B(_6808__bF_buf0), .Y(_6933_) );
INVX1 INVX1_466 ( .gnd(gnd), .vdd(vdd), .A(_6933_), .Y(_6934_) );
NAND2X1 NAND2X1_905 ( .gnd(gnd), .vdd(vdd), .A(_6932_), .B(_6934_), .Y(_6935_) );
XOR2X1 XOR2X1_113 ( .gnd(gnd), .vdd(vdd), .A(_6931_), .B(_6935_), .Y(_6936_) );
OAI21X1 OAI21X1_1947 ( .gnd(gnd), .vdd(vdd), .A(_6936_), .B(_5098__bF_buf3), .C(_5099__bF_buf1), .Y(_6937_) );
AOI21X1 AOI21X1_1189 ( .gnd(gnd), .vdd(vdd), .A(_6930_), .B(_6921_), .C(_6937_), .Y(_6938_) );
OAI21X1 OAI21X1_1948 ( .gnd(gnd), .vdd(vdd), .A(_4819_), .B(_6517__bF_buf2), .C(_6680_), .Y(_6939_) );
OAI21X1 OAI21X1_1949 ( .gnd(gnd), .vdd(vdd), .A(_6784__bF_buf1), .B(_6785__bF_buf1), .C(_4823_), .Y(_6940_) );
NOR2X1 NOR2X1_1205 ( .gnd(gnd), .vdd(vdd), .A(_4823_), .B(_6808__bF_buf4), .Y(_6941_) );
INVX1 INVX1_467 ( .gnd(gnd), .vdd(vdd), .A(_6941_), .Y(_6942_) );
NAND2X1 NAND2X1_906 ( .gnd(gnd), .vdd(vdd), .A(_6940_), .B(_6942_), .Y(_6943_) );
XNOR2X1 XNOR2X1_256 ( .gnd(gnd), .vdd(vdd), .A(_6943_), .B(_6939_), .Y(_6944_) );
OAI21X1 OAI21X1_1950 ( .gnd(gnd), .vdd(vdd), .A(_6944_), .B(_5099__bF_buf0), .C(_5097__bF_buf2), .Y(_6945_) );
AOI21X1 AOI21X1_1190 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_153_), .B(_6293__bF_buf2), .C(_6422_), .Y(_6946_) );
OAI21X1 OAI21X1_1951 ( .gnd(gnd), .vdd(vdd), .A(_6689_), .B(_6946_), .C(_6688_), .Y(_6947_) );
OAI21X1 OAI21X1_1952 ( .gnd(gnd), .vdd(vdd), .A(_6784__bF_buf0), .B(_6785__bF_buf0), .C(_4709_), .Y(_6948_) );
INVX1 INVX1_468 ( .gnd(gnd), .vdd(vdd), .A(_6948_), .Y(_6949_) );
NOR2X1 NOR2X1_1206 ( .gnd(gnd), .vdd(vdd), .A(_4709_), .B(_6808__bF_buf3), .Y(_6950_) );
NOR2X1 NOR2X1_1207 ( .gnd(gnd), .vdd(vdd), .A(_6949_), .B(_6950_), .Y(_6951_) );
XOR2X1 XOR2X1_114 ( .gnd(gnd), .vdd(vdd), .A(_6947_), .B(_6951_), .Y(_6952_) );
AOI21X1 AOI21X1_1191 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe46_bF_buf4), .B(_6952_), .C(micro_hash_ucr_2_pipe48_bF_buf1), .Y(_6953_) );
OAI21X1 OAI21X1_1953 ( .gnd(gnd), .vdd(vdd), .A(_6938_), .B(_6945_), .C(_6953_), .Y(_6954_) );
OAI21X1 OAI21X1_1954 ( .gnd(gnd), .vdd(vdd), .A(_4760_), .B(_6517__bF_buf1), .C(_6695_), .Y(_6955_) );
OAI21X1 OAI21X1_1955 ( .gnd(gnd), .vdd(vdd), .A(_6784__bF_buf4), .B(_6785__bF_buf4), .C(_4764_), .Y(_6956_) );
NOR2X1 NOR2X1_1208 ( .gnd(gnd), .vdd(vdd), .A(_4764_), .B(_6808__bF_buf2), .Y(_6957_) );
INVX1 INVX1_469 ( .gnd(gnd), .vdd(vdd), .A(_6957_), .Y(_6958_) );
NAND2X1 NAND2X1_907 ( .gnd(gnd), .vdd(vdd), .A(_6956_), .B(_6958_), .Y(_6959_) );
AOI21X1 AOI21X1_1192 ( .gnd(gnd), .vdd(vdd), .A(_6955_), .B(_6959_), .C(_5092__bF_buf3), .Y(_6960_) );
OAI21X1 OAI21X1_1956 ( .gnd(gnd), .vdd(vdd), .A(_6955_), .B(_6959_), .C(_6960_), .Y(_6961_) );
AND2X2 AND2X2_462 ( .gnd(gnd), .vdd(vdd), .A(_6961_), .B(_5093__bF_buf3), .Y(_6962_) );
NAND3X1 NAND3X1_310 ( .gnd(gnd), .vdd(vdd), .A(_6699_), .B(_6700_), .C(_6702_), .Y(_6963_) );
OAI21X1 OAI21X1_1957 ( .gnd(gnd), .vdd(vdd), .A(_4732_), .B(_6517__bF_buf0), .C(_6963_), .Y(_6964_) );
OAI21X1 OAI21X1_1958 ( .gnd(gnd), .vdd(vdd), .A(_6784__bF_buf3), .B(_6785__bF_buf3), .C(_4736_), .Y(_6965_) );
NOR2X1 NOR2X1_1209 ( .gnd(gnd), .vdd(vdd), .A(_4736_), .B(_6808__bF_buf1), .Y(_6966_) );
INVX1 INVX1_470 ( .gnd(gnd), .vdd(vdd), .A(_6966_), .Y(_6967_) );
NAND2X1 NAND2X1_908 ( .gnd(gnd), .vdd(vdd), .A(_6965_), .B(_6967_), .Y(_6968_) );
XOR2X1 XOR2X1_115 ( .gnd(gnd), .vdd(vdd), .A(_6964_), .B(_6968_), .Y(_6969_) );
OAI21X1 OAI21X1_1959 ( .gnd(gnd), .vdd(vdd), .A(_6969_), .B(_5093__bF_buf2), .C(_5091__bF_buf3), .Y(_6970_) );
AOI21X1 AOI21X1_1193 ( .gnd(gnd), .vdd(vdd), .A(_6962_), .B(_6954_), .C(_6970_), .Y(_6971_) );
OAI21X1 OAI21X1_1960 ( .gnd(gnd), .vdd(vdd), .A(_4790_), .B(_6517__bF_buf5), .C(_6710_), .Y(_6972_) );
OAI21X1 OAI21X1_1961 ( .gnd(gnd), .vdd(vdd), .A(_6784__bF_buf2), .B(_6785__bF_buf2), .C(_4794_), .Y(_6973_) );
NOR2X1 NOR2X1_1210 ( .gnd(gnd), .vdd(vdd), .A(_4794_), .B(_6808__bF_buf0), .Y(_6974_) );
INVX1 INVX1_471 ( .gnd(gnd), .vdd(vdd), .A(_6974_), .Y(_6975_) );
NAND2X1 NAND2X1_909 ( .gnd(gnd), .vdd(vdd), .A(_6973_), .B(_6975_), .Y(_6976_) );
XNOR2X1 XNOR2X1_257 ( .gnd(gnd), .vdd(vdd), .A(_6976_), .B(_6972_), .Y(_6977_) );
OAI21X1 OAI21X1_1962 ( .gnd(gnd), .vdd(vdd), .A(_6977_), .B(_5091__bF_buf2), .C(_5086__bF_buf3), .Y(_6978_) );
AOI21X1 AOI21X1_1194 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_185_), .B(_6293__bF_buf1), .C(_6444_), .Y(_6979_) );
OAI21X1 OAI21X1_1963 ( .gnd(gnd), .vdd(vdd), .A(_6720_), .B(_6979_), .C(_6719_), .Y(_6980_) );
OAI21X1 OAI21X1_1964 ( .gnd(gnd), .vdd(vdd), .A(_6784__bF_buf1), .B(_6785__bF_buf1), .C(_4852_), .Y(_6981_) );
INVX1 INVX1_472 ( .gnd(gnd), .vdd(vdd), .A(_6981_), .Y(_6982_) );
NOR2X1 NOR2X1_1211 ( .gnd(gnd), .vdd(vdd), .A(_4852_), .B(_6808__bF_buf4), .Y(_6983_) );
NOR2X1 NOR2X1_1212 ( .gnd(gnd), .vdd(vdd), .A(_6982_), .B(_6983_), .Y(_6984_) );
XOR2X1 XOR2X1_116 ( .gnd(gnd), .vdd(vdd), .A(_6980_), .B(_6984_), .Y(_6985_) );
AOI21X1 AOI21X1_1195 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe54_bF_buf3), .B(_6985_), .C(micro_hash_ucr_2_pipe56_bF_buf2), .Y(_6986_) );
OAI21X1 OAI21X1_1965 ( .gnd(gnd), .vdd(vdd), .A(_6971_), .B(_6978_), .C(_6986_), .Y(_6987_) );
OAI21X1 OAI21X1_1966 ( .gnd(gnd), .vdd(vdd), .A(_4820_), .B(_6517__bF_buf4), .C(_6725_), .Y(_6988_) );
OAI21X1 OAI21X1_1967 ( .gnd(gnd), .vdd(vdd), .A(_6784__bF_buf0), .B(_6785__bF_buf0), .C(_4824_), .Y(_6989_) );
NOR2X1 NOR2X1_1213 ( .gnd(gnd), .vdd(vdd), .A(_4824_), .B(_6808__bF_buf3), .Y(_6990_) );
INVX1 INVX1_473 ( .gnd(gnd), .vdd(vdd), .A(_6990_), .Y(_6991_) );
NAND2X1 NAND2X1_910 ( .gnd(gnd), .vdd(vdd), .A(_6989_), .B(_6991_), .Y(_6992_) );
AOI21X1 AOI21X1_1196 ( .gnd(gnd), .vdd(vdd), .A(_6988_), .B(_6992_), .C(_5087__bF_buf3), .Y(_6993_) );
OAI21X1 OAI21X1_1968 ( .gnd(gnd), .vdd(vdd), .A(_6988_), .B(_6992_), .C(_6993_), .Y(_6994_) );
AND2X2 AND2X2_463 ( .gnd(gnd), .vdd(vdd), .A(_6994_), .B(_5085__bF_buf2), .Y(_6995_) );
OAI21X1 OAI21X1_1969 ( .gnd(gnd), .vdd(vdd), .A(_4706_), .B(_6517__bF_buf3), .C(_6735_), .Y(_6996_) );
OAI21X1 OAI21X1_1970 ( .gnd(gnd), .vdd(vdd), .A(_6784__bF_buf4), .B(_6785__bF_buf4), .C(_4710_), .Y(_6997_) );
NOR2X1 NOR2X1_1214 ( .gnd(gnd), .vdd(vdd), .A(_4710_), .B(_6808__bF_buf2), .Y(_6998_) );
INVX1 INVX1_474 ( .gnd(gnd), .vdd(vdd), .A(_6998_), .Y(_6999_) );
NAND2X1 NAND2X1_911 ( .gnd(gnd), .vdd(vdd), .A(_6997_), .B(_6999_), .Y(_7000_) );
XOR2X1 XOR2X1_117 ( .gnd(gnd), .vdd(vdd), .A(_6996_), .B(_7000_), .Y(_7001_) );
OAI21X1 OAI21X1_1971 ( .gnd(gnd), .vdd(vdd), .A(_7001_), .B(_5085__bF_buf1), .C(_5080__bF_buf0), .Y(_7002_) );
AOI21X1 AOI21X1_1197 ( .gnd(gnd), .vdd(vdd), .A(_6995_), .B(_6987_), .C(_7002_), .Y(_7003_) );
AOI21X1 AOI21X1_1198 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_209_), .B(_6293__bF_buf0), .C(_6464_), .Y(_7004_) );
OAI21X1 OAI21X1_1972 ( .gnd(gnd), .vdd(vdd), .A(_6743_), .B(_7004_), .C(_6742_), .Y(_7005_) );
OAI21X1 OAI21X1_1973 ( .gnd(gnd), .vdd(vdd), .A(_6784__bF_buf3), .B(_6785__bF_buf3), .C(_4765_), .Y(_7006_) );
NOR2X1 NOR2X1_1215 ( .gnd(gnd), .vdd(vdd), .A(_4765_), .B(_6808__bF_buf1), .Y(_7007_) );
INVX1 INVX1_475 ( .gnd(gnd), .vdd(vdd), .A(_7007_), .Y(_7008_) );
NAND2X1 NAND2X1_912 ( .gnd(gnd), .vdd(vdd), .A(_7006_), .B(_7008_), .Y(_7009_) );
XNOR2X1 XNOR2X1_258 ( .gnd(gnd), .vdd(vdd), .A(_7005_), .B(_7009_), .Y(_7010_) );
OAI21X1 OAI21X1_1974 ( .gnd(gnd), .vdd(vdd), .A(_7010_), .B(_5080__bF_buf3), .C(_5081__bF_buf1), .Y(_7011_) );
OAI21X1 OAI21X1_1975 ( .gnd(gnd), .vdd(vdd), .A(_6472_), .B(_6470_), .C(_6749_), .Y(_7012_) );
OAI21X1 OAI21X1_1976 ( .gnd(gnd), .vdd(vdd), .A(_4733_), .B(_6517__bF_buf2), .C(_7012_), .Y(_7013_) );
OAI21X1 OAI21X1_1977 ( .gnd(gnd), .vdd(vdd), .A(_6784__bF_buf2), .B(_6785__bF_buf2), .C(_4737_), .Y(_7014_) );
INVX1 INVX1_476 ( .gnd(gnd), .vdd(vdd), .A(_7014_), .Y(_7015_) );
NOR2X1 NOR2X1_1216 ( .gnd(gnd), .vdd(vdd), .A(_4737_), .B(_6808__bF_buf0), .Y(_7016_) );
NOR2X1 NOR2X1_1217 ( .gnd(gnd), .vdd(vdd), .A(_7015_), .B(_7016_), .Y(_7017_) );
XOR2X1 XOR2X1_118 ( .gnd(gnd), .vdd(vdd), .A(_7017_), .B(_7013_), .Y(_7018_) );
AOI21X1 AOI21X1_1199 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe62_bF_buf0), .B(_7018_), .C(micro_hash_ucr_2_pipe64_bF_buf3), .Y(_7019_) );
OAI21X1 OAI21X1_1978 ( .gnd(gnd), .vdd(vdd), .A(_7003_), .B(_7011_), .C(_7019_), .Y(_7020_) );
NAND3X1 NAND3X1_311 ( .gnd(gnd), .vdd(vdd), .A(_6503_), .B(_6515_), .C(_6519_), .Y(_7021_) );
OAI21X1 OAI21X1_1979 ( .gnd(gnd), .vdd(vdd), .A(_6504_), .B(_6517__bF_buf1), .C(_7021_), .Y(_7022_) );
INVX1 INVX1_477 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_227_), .Y(_7023_) );
OAI21X1 OAI21X1_1980 ( .gnd(gnd), .vdd(vdd), .A(_6784__bF_buf1), .B(_6785__bF_buf1), .C(_7023_), .Y(_7024_) );
NOR2X1 NOR2X1_1218 ( .gnd(gnd), .vdd(vdd), .A(_7023_), .B(_6808__bF_buf4), .Y(_7025_) );
INVX1 INVX1_478 ( .gnd(gnd), .vdd(vdd), .A(_7025_), .Y(_7026_) );
NAND2X1 NAND2X1_913 ( .gnd(gnd), .vdd(vdd), .A(_7024_), .B(_7026_), .Y(_7027_) );
AOI21X1 AOI21X1_1200 ( .gnd(gnd), .vdd(vdd), .A(_7027_), .B(_7022_), .C(_5079__bF_buf1), .Y(_7028_) );
OAI21X1 OAI21X1_1981 ( .gnd(gnd), .vdd(vdd), .A(_7022_), .B(_7027_), .C(_7028_), .Y(_7029_) );
AND2X2 AND2X2_464 ( .gnd(gnd), .vdd(vdd), .A(_7029_), .B(_5074__bF_buf0), .Y(_7030_) );
OAI21X1 OAI21X1_1982 ( .gnd(gnd), .vdd(vdd), .A(_6755_), .B(_6517__bF_buf0), .C(_6758_), .Y(_7031_) );
INVX1 INVX1_479 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_235_), .Y(_7032_) );
OAI21X1 OAI21X1_1983 ( .gnd(gnd), .vdd(vdd), .A(_6784__bF_buf0), .B(_6785__bF_buf0), .C(_7032_), .Y(_7033_) );
NOR2X1 NOR2X1_1219 ( .gnd(gnd), .vdd(vdd), .A(_7032_), .B(_6808__bF_buf3), .Y(_7034_) );
INVX1 INVX1_480 ( .gnd(gnd), .vdd(vdd), .A(_7034_), .Y(_7035_) );
NAND2X1 NAND2X1_914 ( .gnd(gnd), .vdd(vdd), .A(_7033_), .B(_7035_), .Y(_7036_) );
XOR2X1 XOR2X1_119 ( .gnd(gnd), .vdd(vdd), .A(_7036_), .B(_7031_), .Y(_7037_) );
OAI21X1 OAI21X1_1984 ( .gnd(gnd), .vdd(vdd), .A(_7037_), .B(_5074__bF_buf3), .C(_5075__bF_buf2), .Y(_7038_) );
AOI21X1 AOI21X1_1201 ( .gnd(gnd), .vdd(vdd), .A(_7030_), .B(_7020_), .C(_7038_), .Y(_7039_) );
NAND3X1 NAND3X1_312 ( .gnd(gnd), .vdd(vdd), .A(_6763_), .B(_6765_), .C(_6767_), .Y(_7040_) );
OAI21X1 OAI21X1_1985 ( .gnd(gnd), .vdd(vdd), .A(_6764_), .B(_6517__bF_buf5), .C(_7040_), .Y(_7041_) );
INVX1 INVX1_481 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_243_), .Y(_7042_) );
OAI21X1 OAI21X1_1986 ( .gnd(gnd), .vdd(vdd), .A(_6784__bF_buf4), .B(_6785__bF_buf4), .C(_7042_), .Y(_7043_) );
INVX1 INVX1_482 ( .gnd(gnd), .vdd(vdd), .A(_7043_), .Y(_7044_) );
NOR2X1 NOR2X1_1220 ( .gnd(gnd), .vdd(vdd), .A(_7042_), .B(_6808__bF_buf2), .Y(_7045_) );
NOR2X1 NOR2X1_1221 ( .gnd(gnd), .vdd(vdd), .A(_7044_), .B(_7045_), .Y(_7046_) );
XOR2X1 XOR2X1_120 ( .gnd(gnd), .vdd(vdd), .A(_7041_), .B(_7046_), .Y(_7047_) );
OAI21X1 OAI21X1_1987 ( .gnd(gnd), .vdd(vdd), .A(_7047_), .B(_5075__bF_buf1), .C(_6146_), .Y(_7048_) );
NOR2X1 NOR2X1_1222 ( .gnd(gnd), .vdd(vdd), .A(_6776_), .B(_6778_), .Y(_7049_) );
INVX2 INVX2_240 ( .gnd(gnd), .vdd(vdd), .A(_7049_), .Y(_7050_) );
INVX1 INVX1_483 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_251_), .Y(_7051_) );
OAI21X1 OAI21X1_1988 ( .gnd(gnd), .vdd(vdd), .A(_6784__bF_buf3), .B(_6785__bF_buf3), .C(_7051_), .Y(_7052_) );
INVX1 INVX1_484 ( .gnd(gnd), .vdd(vdd), .A(_7052_), .Y(_7053_) );
NOR2X1 NOR2X1_1223 ( .gnd(gnd), .vdd(vdd), .A(_7051_), .B(_6808__bF_buf1), .Y(_7054_) );
NOR2X1 NOR2X1_1224 ( .gnd(gnd), .vdd(vdd), .A(_7053_), .B(_7054_), .Y(_7055_) );
AND2X2 AND2X2_465 ( .gnd(gnd), .vdd(vdd), .A(_7050_), .B(_7055_), .Y(_7056_) );
OAI21X1 OAI21X1_1989 ( .gnd(gnd), .vdd(vdd), .A(_7050_), .B(_7055_), .C(_4563_), .Y(_7057_) );
OAI22X1 OAI22X1_100 ( .gnd(gnd), .vdd(vdd), .A(_7056_), .B(_7057_), .C(_7039_), .D(_7048_), .Y(_4493__3_) );
AOI21X1 AOI21X1_1202 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_k_3_), .B(micro_hash_ucr_2_x_3_), .C(_6784__bF_buf2), .Y(_7058_) );
NOR2X1 NOR2X1_1225 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_k_4_), .B(micro_hash_ucr_2_x_4_), .Y(_7059_) );
INVX1 INVX1_485 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_k_4_), .Y(_7060_) );
INVX1 INVX1_486 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_x_4_), .Y(_7061_) );
NOR2X1 NOR2X1_1226 ( .gnd(gnd), .vdd(vdd), .A(_7060_), .B(_7061_), .Y(_7062_) );
NOR2X1 NOR2X1_1227 ( .gnd(gnd), .vdd(vdd), .A(_7059_), .B(_7062_), .Y(_7063_) );
INVX1 INVX1_487 ( .gnd(gnd), .vdd(vdd), .A(_7063_), .Y(_7064_) );
OR2X2 OR2X2_54 ( .gnd(gnd), .vdd(vdd), .A(_7058_), .B(_7064_), .Y(_7065_) );
OAI21X1 OAI21X1_1990 ( .gnd(gnd), .vdd(vdd), .A(_7059_), .B(_7062_), .C(_7058_), .Y(_7066_) );
NAND2X1 NAND2X1_915 ( .gnd(gnd), .vdd(vdd), .A(_7066_), .B(_7065_), .Y(_7067_) );
XNOR2X1 XNOR2X1_259 ( .gnd(gnd), .vdd(vdd), .A(_7067__bF_buf5), .B(micro_hash_ucr_2_Wx_4_), .Y(_7068_) );
OAI21X1 OAI21X1_1991 ( .gnd(gnd), .vdd(vdd), .A(_6781_), .B(_6808__bF_buf0), .C(_6780_), .Y(_7069_) );
AND2X2 AND2X2_466 ( .gnd(gnd), .vdd(vdd), .A(_7069_), .B(_6786_), .Y(_7070_) );
NOR2X1 NOR2X1_1228 ( .gnd(gnd), .vdd(vdd), .A(_7068_), .B(_7070_), .Y(_7071_) );
AND2X2 AND2X2_467 ( .gnd(gnd), .vdd(vdd), .A(_7070_), .B(_7068_), .Y(_7072_) );
OAI21X1 OAI21X1_1992 ( .gnd(gnd), .vdd(vdd), .A(_7072_), .B(_7071_), .C(micro_hash_ucr_2_pipe8), .Y(_7073_) );
XOR2X1 XOR2X1_121 ( .gnd(gnd), .vdd(vdd), .A(_7067__bF_buf4), .B(micro_hash_ucr_2_Wx_12_), .Y(_7074_) );
INVX1 INVX1_488 ( .gnd(gnd), .vdd(vdd), .A(_6798_), .Y(_7075_) );
OAI21X1 OAI21X1_1993 ( .gnd(gnd), .vdd(vdd), .A(_6796_), .B(_7075_), .C(_6799_), .Y(_7076_) );
XNOR2X1 XNOR2X1_260 ( .gnd(gnd), .vdd(vdd), .A(_7076_), .B(_7074_), .Y(_7077_) );
NAND2X1 NAND2X1_916 ( .gnd(gnd), .vdd(vdd), .A(_5592_), .B(_5134_), .Y(_7078_) );
OAI21X1 OAI21X1_1994 ( .gnd(gnd), .vdd(vdd), .A(H_2_20_), .B(_5134_), .C(_7078_), .Y(_7079_) );
AOI21X1 AOI21X1_1203 ( .gnd(gnd), .vdd(vdd), .A(_5135_), .B(_7079_), .C(micro_hash_ucr_2_pipe10), .Y(_7080_) );
AOI22X1 AOI22X1_54 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe10), .B(_7077_), .C(_7073_), .D(_7080_), .Y(_7081_) );
INVX2 INVX2_241 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_20_), .Y(_7082_) );
XNOR2X1 XNOR2X1_261 ( .gnd(gnd), .vdd(vdd), .A(_7067__bF_buf3), .B(_7082_), .Y(_7083_) );
AOI21X1 AOI21X1_1204 ( .gnd(gnd), .vdd(vdd), .A(_6807_), .B(_6805_), .C(_6809_), .Y(_7084_) );
NAND2X1 NAND2X1_917 ( .gnd(gnd), .vdd(vdd), .A(_7084_), .B(_7083_), .Y(_7085_) );
NOR2X1 NOR2X1_1229 ( .gnd(gnd), .vdd(vdd), .A(_7084_), .B(_7083_), .Y(_7086_) );
INVX1 INVX1_489 ( .gnd(gnd), .vdd(vdd), .A(_7086_), .Y(_7087_) );
NAND3X1 NAND3X1_313 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe12_bF_buf1), .B(_7085_), .C(_7087_), .Y(_7088_) );
OAI21X1 OAI21X1_1995 ( .gnd(gnd), .vdd(vdd), .A(_7081_), .B(micro_hash_ucr_2_pipe12_bF_buf0), .C(_7088_), .Y(_7089_) );
XOR2X1 XOR2X1_122 ( .gnd(gnd), .vdd(vdd), .A(_7067__bF_buf2), .B(micro_hash_ucr_2_Wx_28_), .Y(_7090_) );
AOI21X1 AOI21X1_1205 ( .gnd(gnd), .vdd(vdd), .A(_6817_), .B(_6815_), .C(_6819_), .Y(_7091_) );
NOR2X1 NOR2X1_1230 ( .gnd(gnd), .vdd(vdd), .A(_7091_), .B(_7090_), .Y(_7092_) );
AND2X2 AND2X2_468 ( .gnd(gnd), .vdd(vdd), .A(_7090_), .B(_7091_), .Y(_7093_) );
OAI21X1 OAI21X1_1996 ( .gnd(gnd), .vdd(vdd), .A(_7093_), .B(_7092_), .C(micro_hash_ucr_2_pipe14_bF_buf4), .Y(_7094_) );
OAI21X1 OAI21X1_1997 ( .gnd(gnd), .vdd(vdd), .A(_7089_), .B(micro_hash_ucr_2_pipe14_bF_buf3), .C(_7094_), .Y(_7095_) );
XNOR2X1 XNOR2X1_262 ( .gnd(gnd), .vdd(vdd), .A(_7067__bF_buf1), .B(micro_hash_ucr_2_Wx_36_), .Y(_7096_) );
INVX1 INVX1_490 ( .gnd(gnd), .vdd(vdd), .A(_7096_), .Y(_7097_) );
AOI21X1 AOI21X1_1206 ( .gnd(gnd), .vdd(vdd), .A(_6827_), .B(_6825_), .C(_6828_), .Y(_7098_) );
AND2X2 AND2X2_469 ( .gnd(gnd), .vdd(vdd), .A(_7098_), .B(_7097_), .Y(_7099_) );
NOR2X1 NOR2X1_1231 ( .gnd(gnd), .vdd(vdd), .A(_7097_), .B(_7098_), .Y(_7100_) );
NOR2X1 NOR2X1_1232 ( .gnd(gnd), .vdd(vdd), .A(_7100_), .B(_7099_), .Y(_7101_) );
NAND2X1 NAND2X1_918 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe16_bF_buf1), .B(_7101_), .Y(_7102_) );
OAI21X1 OAI21X1_1998 ( .gnd(gnd), .vdd(vdd), .A(_7095_), .B(micro_hash_ucr_2_pipe16_bF_buf0), .C(_7102_), .Y(_7103_) );
XOR2X1 XOR2X1_123 ( .gnd(gnd), .vdd(vdd), .A(_7067__bF_buf0), .B(micro_hash_ucr_2_Wx_44_), .Y(_7104_) );
AOI21X1 AOI21X1_1207 ( .gnd(gnd), .vdd(vdd), .A(_6836_), .B(_6834_), .C(_6837_), .Y(_7105_) );
NOR2X1 NOR2X1_1233 ( .gnd(gnd), .vdd(vdd), .A(_7104_), .B(_7105_), .Y(_7106_) );
AND2X2 AND2X2_470 ( .gnd(gnd), .vdd(vdd), .A(_7105_), .B(_7104_), .Y(_7107_) );
OAI21X1 OAI21X1_1999 ( .gnd(gnd), .vdd(vdd), .A(_7107_), .B(_7106_), .C(micro_hash_ucr_2_pipe18_bF_buf3), .Y(_7108_) );
OAI21X1 OAI21X1_2000 ( .gnd(gnd), .vdd(vdd), .A(_7103_), .B(micro_hash_ucr_2_pipe18_bF_buf2), .C(_7108_), .Y(_7109_) );
XNOR2X1 XNOR2X1_263 ( .gnd(gnd), .vdd(vdd), .A(_7067__bF_buf5), .B(micro_hash_ucr_2_Wx_52_), .Y(_7110_) );
INVX1 INVX1_491 ( .gnd(gnd), .vdd(vdd), .A(_7110_), .Y(_7111_) );
AOI21X1 AOI21X1_1208 ( .gnd(gnd), .vdd(vdd), .A(_6846_), .B(_6844_), .C(_6847_), .Y(_7112_) );
NAND2X1 NAND2X1_919 ( .gnd(gnd), .vdd(vdd), .A(_7111_), .B(_7112_), .Y(_7113_) );
NOR2X1 NOR2X1_1234 ( .gnd(gnd), .vdd(vdd), .A(_7111_), .B(_7112_), .Y(_7114_) );
INVX1 INVX1_492 ( .gnd(gnd), .vdd(vdd), .A(_7114_), .Y(_7115_) );
NAND3X1 NAND3X1_314 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe20_bF_buf0), .B(_7113_), .C(_7115_), .Y(_7116_) );
OAI21X1 OAI21X1_2001 ( .gnd(gnd), .vdd(vdd), .A(_7109_), .B(micro_hash_ucr_2_pipe20_bF_buf3), .C(_7116_), .Y(_7117_) );
XNOR2X1 XNOR2X1_264 ( .gnd(gnd), .vdd(vdd), .A(_7067__bF_buf4), .B(micro_hash_ucr_2_Wx_60_), .Y(_7118_) );
INVX1 INVX1_493 ( .gnd(gnd), .vdd(vdd), .A(_7118_), .Y(_7119_) );
AOI21X1 AOI21X1_1209 ( .gnd(gnd), .vdd(vdd), .A(_6853_), .B(_6852_), .C(_6855_), .Y(_7120_) );
NAND2X1 NAND2X1_920 ( .gnd(gnd), .vdd(vdd), .A(_7120_), .B(_7119_), .Y(_7121_) );
NOR2X1 NOR2X1_1235 ( .gnd(gnd), .vdd(vdd), .A(_7120_), .B(_7119_), .Y(_7122_) );
INVX1 INVX1_494 ( .gnd(gnd), .vdd(vdd), .A(_7122_), .Y(_7123_) );
NAND2X1 NAND2X1_921 ( .gnd(gnd), .vdd(vdd), .A(_7121_), .B(_7123_), .Y(_7124_) );
OAI21X1 OAI21X1_2002 ( .gnd(gnd), .vdd(vdd), .A(_7124_), .B(_5121__bF_buf4), .C(_5116__bF_buf4), .Y(_7125_) );
AOI21X1 AOI21X1_1210 ( .gnd(gnd), .vdd(vdd), .A(_5121__bF_buf3), .B(_7117_), .C(_7125_), .Y(_7126_) );
XNOR2X1 XNOR2X1_265 ( .gnd(gnd), .vdd(vdd), .A(_7067__bF_buf3), .B(micro_hash_ucr_2_Wx_68_), .Y(_7127_) );
AOI21X1 AOI21X1_1211 ( .gnd(gnd), .vdd(vdd), .A(_6861_), .B(_6860_), .C(_6862_), .Y(_7128_) );
XOR2X1 XOR2X1_124 ( .gnd(gnd), .vdd(vdd), .A(_7128_), .B(_7127_), .Y(_7129_) );
AOI21X1 AOI21X1_1212 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe24_bF_buf3), .B(_7129_), .C(_7126_), .Y(_7130_) );
XNOR2X1 XNOR2X1_266 ( .gnd(gnd), .vdd(vdd), .A(_7067__bF_buf2), .B(_5038_), .Y(_7131_) );
AOI21X1 AOI21X1_1213 ( .gnd(gnd), .vdd(vdd), .A(_6869_), .B(_6868_), .C(_6870_), .Y(_7132_) );
NOR2X1 NOR2X1_1236 ( .gnd(gnd), .vdd(vdd), .A(_7131_), .B(_7132_), .Y(_7133_) );
AND2X2 AND2X2_471 ( .gnd(gnd), .vdd(vdd), .A(_7132_), .B(_7131_), .Y(_7134_) );
OAI21X1 OAI21X1_2003 ( .gnd(gnd), .vdd(vdd), .A(_7134_), .B(_7133_), .C(micro_hash_ucr_2_pipe26_bF_buf0), .Y(_7135_) );
OAI21X1 OAI21X1_2004 ( .gnd(gnd), .vdd(vdd), .A(_7130_), .B(micro_hash_ucr_2_pipe26_bF_buf3), .C(_7135_), .Y(_7136_) );
XNOR2X1 XNOR2X1_267 ( .gnd(gnd), .vdd(vdd), .A(_7067__bF_buf1), .B(micro_hash_ucr_2_Wx_84_), .Y(_7137_) );
INVX1 INVX1_495 ( .gnd(gnd), .vdd(vdd), .A(_7137_), .Y(_7138_) );
AOI21X1 AOI21X1_1214 ( .gnd(gnd), .vdd(vdd), .A(_6878_), .B(_6877_), .C(_6879_), .Y(_7139_) );
NAND2X1 NAND2X1_922 ( .gnd(gnd), .vdd(vdd), .A(_7138_), .B(_7139_), .Y(_7140_) );
NOR2X1 NOR2X1_1237 ( .gnd(gnd), .vdd(vdd), .A(_7138_), .B(_7139_), .Y(_7141_) );
INVX1 INVX1_496 ( .gnd(gnd), .vdd(vdd), .A(_7141_), .Y(_7142_) );
NAND3X1 NAND3X1_315 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe28_bF_buf2), .B(_7140_), .C(_7142_), .Y(_7143_) );
OAI21X1 OAI21X1_2005 ( .gnd(gnd), .vdd(vdd), .A(_7136_), .B(micro_hash_ucr_2_pipe28_bF_buf1), .C(_7143_), .Y(_7144_) );
XNOR2X1 XNOR2X1_268 ( .gnd(gnd), .vdd(vdd), .A(_7067__bF_buf0), .B(micro_hash_ucr_2_Wx_92_), .Y(_7145_) );
INVX1 INVX1_497 ( .gnd(gnd), .vdd(vdd), .A(_7145_), .Y(_7146_) );
AOI21X1 AOI21X1_1215 ( .gnd(gnd), .vdd(vdd), .A(_6885_), .B(_6884_), .C(_6887_), .Y(_7147_) );
NOR2X1 NOR2X1_1238 ( .gnd(gnd), .vdd(vdd), .A(_7147_), .B(_7146_), .Y(_7148_) );
INVX1 INVX1_498 ( .gnd(gnd), .vdd(vdd), .A(_7148_), .Y(_7149_) );
AOI21X1 AOI21X1_1216 ( .gnd(gnd), .vdd(vdd), .A(_7147_), .B(_7146_), .C(_5110__bF_buf1), .Y(_7150_) );
AOI22X1 AOI22X1_55 ( .gnd(gnd), .vdd(vdd), .A(_7149_), .B(_7150_), .C(_7144_), .D(_5110__bF_buf0), .Y(_7151_) );
NAND2X1 NAND2X1_923 ( .gnd(gnd), .vdd(vdd), .A(_5111__bF_buf0), .B(_7151_), .Y(_7152_) );
XNOR2X1 XNOR2X1_269 ( .gnd(gnd), .vdd(vdd), .A(_7067__bF_buf5), .B(micro_hash_ucr_2_Wx_100_), .Y(_7153_) );
INVX1 INVX1_499 ( .gnd(gnd), .vdd(vdd), .A(_7153_), .Y(_7154_) );
AOI21X1 AOI21X1_1217 ( .gnd(gnd), .vdd(vdd), .A(_6894_), .B(_6893_), .C(_6895_), .Y(_7155_) );
AND2X2 AND2X2_472 ( .gnd(gnd), .vdd(vdd), .A(_7155_), .B(_7154_), .Y(_7156_) );
NOR2X1 NOR2X1_1239 ( .gnd(gnd), .vdd(vdd), .A(_7154_), .B(_7155_), .Y(_7157_) );
OAI21X1 OAI21X1_2006 ( .gnd(gnd), .vdd(vdd), .A(_7156_), .B(_7157_), .C(micro_hash_ucr_2_pipe32_bF_buf0), .Y(_7158_) );
AOI21X1 AOI21X1_1218 ( .gnd(gnd), .vdd(vdd), .A(_7158_), .B(_7152_), .C(micro_hash_ucr_2_pipe34_bF_buf2), .Y(_7159_) );
XNOR2X1 XNOR2X1_270 ( .gnd(gnd), .vdd(vdd), .A(_7067__bF_buf4), .B(micro_hash_ucr_2_Wx_108_), .Y(_7160_) );
INVX1 INVX1_500 ( .gnd(gnd), .vdd(vdd), .A(_7160_), .Y(_7161_) );
AOI21X1 AOI21X1_1219 ( .gnd(gnd), .vdd(vdd), .A(_6902_), .B(_6901_), .C(_6903_), .Y(_7162_) );
NAND2X1 NAND2X1_924 ( .gnd(gnd), .vdd(vdd), .A(_7161_), .B(_7162_), .Y(_7163_) );
NOR2X1 NOR2X1_1240 ( .gnd(gnd), .vdd(vdd), .A(_7161_), .B(_7162_), .Y(_7164_) );
INVX1 INVX1_501 ( .gnd(gnd), .vdd(vdd), .A(_7164_), .Y(_7165_) );
AOI21X1 AOI21X1_1220 ( .gnd(gnd), .vdd(vdd), .A(_7163_), .B(_7165_), .C(_5109__bF_buf2), .Y(_7166_) );
OAI21X1 OAI21X1_2007 ( .gnd(gnd), .vdd(vdd), .A(_7159_), .B(_7166_), .C(_5104__bF_buf2), .Y(_7167_) );
XNOR2X1 XNOR2X1_271 ( .gnd(gnd), .vdd(vdd), .A(_7067__bF_buf3), .B(micro_hash_ucr_2_Wx_116_), .Y(_7168_) );
OAI21X1 OAI21X1_2008 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_115_), .B(_6787_), .C(_6910_), .Y(_7169_) );
OAI21X1 OAI21X1_2009 ( .gnd(gnd), .vdd(vdd), .A(_4922_), .B(_6808__bF_buf4), .C(_7169_), .Y(_7170_) );
NOR2X1 NOR2X1_1241 ( .gnd(gnd), .vdd(vdd), .A(_7168_), .B(_7170_), .Y(_7171_) );
NAND2X1 NAND2X1_925 ( .gnd(gnd), .vdd(vdd), .A(_7168_), .B(_7170_), .Y(_7172_) );
INVX1 INVX1_502 ( .gnd(gnd), .vdd(vdd), .A(_7172_), .Y(_7173_) );
OAI21X1 OAI21X1_2010 ( .gnd(gnd), .vdd(vdd), .A(_7173_), .B(_7171_), .C(micro_hash_ucr_2_pipe36_bF_buf1), .Y(_7174_) );
NAND3X1 NAND3X1_316 ( .gnd(gnd), .vdd(vdd), .A(_5105__bF_buf1), .B(_7174_), .C(_7167_), .Y(_7175_) );
XNOR2X1 XNOR2X1_272 ( .gnd(gnd), .vdd(vdd), .A(_7067__bF_buf2), .B(micro_hash_ucr_2_Wx_124_), .Y(_7176_) );
INVX1 INVX1_503 ( .gnd(gnd), .vdd(vdd), .A(_7176_), .Y(_7177_) );
AOI21X1 AOI21X1_1221 ( .gnd(gnd), .vdd(vdd), .A(_6915_), .B(_6914_), .C(_6916_), .Y(_7178_) );
NOR2X1 NOR2X1_1242 ( .gnd(gnd), .vdd(vdd), .A(_7177_), .B(_7178_), .Y(_7179_) );
INVX1 INVX1_504 ( .gnd(gnd), .vdd(vdd), .A(_7179_), .Y(_7180_) );
NAND2X1 NAND2X1_926 ( .gnd(gnd), .vdd(vdd), .A(_7177_), .B(_7178_), .Y(_7181_) );
NAND2X1 NAND2X1_927 ( .gnd(gnd), .vdd(vdd), .A(_7181_), .B(_7180_), .Y(_7182_) );
OAI21X1 OAI21X1_2011 ( .gnd(gnd), .vdd(vdd), .A(_5105__bF_buf0), .B(_7182_), .C(_7175_), .Y(_7183_) );
NOR2X1 NOR2X1_1243 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe40_bF_buf2), .B(_7183_), .Y(_7184_) );
XNOR2X1 XNOR2X1_273 ( .gnd(gnd), .vdd(vdd), .A(_7067__bF_buf1), .B(micro_hash_ucr_2_Wx_132_), .Y(_7185_) );
INVX1 INVX1_505 ( .gnd(gnd), .vdd(vdd), .A(_7185_), .Y(_7186_) );
AOI21X1 AOI21X1_1222 ( .gnd(gnd), .vdd(vdd), .A(_6924_), .B(_6923_), .C(_6925_), .Y(_7187_) );
NAND2X1 NAND2X1_928 ( .gnd(gnd), .vdd(vdd), .A(_7186_), .B(_7187_), .Y(_7188_) );
NOR2X1 NOR2X1_1244 ( .gnd(gnd), .vdd(vdd), .A(_7186_), .B(_7187_), .Y(_7189_) );
INVX1 INVX1_506 ( .gnd(gnd), .vdd(vdd), .A(_7189_), .Y(_7190_) );
AOI21X1 AOI21X1_1223 ( .gnd(gnd), .vdd(vdd), .A(_7188_), .B(_7190_), .C(_5103__bF_buf2), .Y(_7191_) );
OAI21X1 OAI21X1_2012 ( .gnd(gnd), .vdd(vdd), .A(_7184_), .B(_7191_), .C(_5098__bF_buf2), .Y(_7192_) );
XNOR2X1 XNOR2X1_274 ( .gnd(gnd), .vdd(vdd), .A(_7067__bF_buf0), .B(micro_hash_ucr_2_Wx_140_), .Y(_7193_) );
INVX1 INVX1_507 ( .gnd(gnd), .vdd(vdd), .A(_7193_), .Y(_7194_) );
AOI21X1 AOI21X1_1224 ( .gnd(gnd), .vdd(vdd), .A(_6932_), .B(_6931_), .C(_6933_), .Y(_7195_) );
AND2X2 AND2X2_473 ( .gnd(gnd), .vdd(vdd), .A(_7195_), .B(_7194_), .Y(_7196_) );
NOR2X1 NOR2X1_1245 ( .gnd(gnd), .vdd(vdd), .A(_7194_), .B(_7195_), .Y(_7197_) );
OAI21X1 OAI21X1_2013 ( .gnd(gnd), .vdd(vdd), .A(_7196_), .B(_7197_), .C(micro_hash_ucr_2_pipe42_bF_buf1), .Y(_7198_) );
NAND3X1 NAND3X1_317 ( .gnd(gnd), .vdd(vdd), .A(_5099__bF_buf4), .B(_7198_), .C(_7192_), .Y(_7199_) );
XNOR2X1 XNOR2X1_275 ( .gnd(gnd), .vdd(vdd), .A(_7067__bF_buf5), .B(micro_hash_ucr_2_Wx_148_), .Y(_7200_) );
INVX1 INVX1_508 ( .gnd(gnd), .vdd(vdd), .A(_7200_), .Y(_7201_) );
AOI21X1 AOI21X1_1225 ( .gnd(gnd), .vdd(vdd), .A(_6940_), .B(_6939_), .C(_6941_), .Y(_7202_) );
NOR2X1 NOR2X1_1246 ( .gnd(gnd), .vdd(vdd), .A(_7202_), .B(_7201_), .Y(_7203_) );
INVX1 INVX1_509 ( .gnd(gnd), .vdd(vdd), .A(_7203_), .Y(_7204_) );
NAND2X1 NAND2X1_929 ( .gnd(gnd), .vdd(vdd), .A(_7202_), .B(_7201_), .Y(_7205_) );
NAND2X1 NAND2X1_930 ( .gnd(gnd), .vdd(vdd), .A(_7205_), .B(_7204_), .Y(_7206_) );
OAI21X1 OAI21X1_2014 ( .gnd(gnd), .vdd(vdd), .A(_5099__bF_buf3), .B(_7206_), .C(_7199_), .Y(_7207_) );
NOR2X1 NOR2X1_1247 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe46_bF_buf3), .B(_7207_), .Y(_7208_) );
XNOR2X1 XNOR2X1_276 ( .gnd(gnd), .vdd(vdd), .A(_7067__bF_buf4), .B(micro_hash_ucr_2_Wx_156_), .Y(_7209_) );
INVX1 INVX1_510 ( .gnd(gnd), .vdd(vdd), .A(_7209_), .Y(_7210_) );
AOI21X1 AOI21X1_1226 ( .gnd(gnd), .vdd(vdd), .A(_6948_), .B(_6947_), .C(_6950_), .Y(_7211_) );
NAND2X1 NAND2X1_931 ( .gnd(gnd), .vdd(vdd), .A(_7210_), .B(_7211_), .Y(_7212_) );
NOR2X1 NOR2X1_1248 ( .gnd(gnd), .vdd(vdd), .A(_7210_), .B(_7211_), .Y(_7213_) );
INVX1 INVX1_511 ( .gnd(gnd), .vdd(vdd), .A(_7213_), .Y(_7214_) );
AOI21X1 AOI21X1_1227 ( .gnd(gnd), .vdd(vdd), .A(_7212_), .B(_7214_), .C(_5097__bF_buf1), .Y(_7215_) );
OAI21X1 OAI21X1_2015 ( .gnd(gnd), .vdd(vdd), .A(_7208_), .B(_7215_), .C(_5092__bF_buf2), .Y(_7216_) );
XNOR2X1 XNOR2X1_277 ( .gnd(gnd), .vdd(vdd), .A(_7067__bF_buf3), .B(micro_hash_ucr_2_Wx_164_), .Y(_7217_) );
INVX1 INVX1_512 ( .gnd(gnd), .vdd(vdd), .A(_7217_), .Y(_7218_) );
AOI21X1 AOI21X1_1228 ( .gnd(gnd), .vdd(vdd), .A(_6956_), .B(_6955_), .C(_6957_), .Y(_7219_) );
AND2X2 AND2X2_474 ( .gnd(gnd), .vdd(vdd), .A(_7218_), .B(_7219_), .Y(_7220_) );
NOR2X1 NOR2X1_1249 ( .gnd(gnd), .vdd(vdd), .A(_7219_), .B(_7218_), .Y(_7221_) );
OAI21X1 OAI21X1_2016 ( .gnd(gnd), .vdd(vdd), .A(_7220_), .B(_7221_), .C(micro_hash_ucr_2_pipe48_bF_buf0), .Y(_7222_) );
NAND3X1 NAND3X1_318 ( .gnd(gnd), .vdd(vdd), .A(_5093__bF_buf1), .B(_7222_), .C(_7216_), .Y(_7223_) );
XNOR2X1 XNOR2X1_278 ( .gnd(gnd), .vdd(vdd), .A(_7067__bF_buf2), .B(micro_hash_ucr_2_Wx_172_), .Y(_7224_) );
INVX1 INVX1_513 ( .gnd(gnd), .vdd(vdd), .A(_7224_), .Y(_7225_) );
AOI21X1 AOI21X1_1229 ( .gnd(gnd), .vdd(vdd), .A(_6965_), .B(_6964_), .C(_6966_), .Y(_7226_) );
OR2X2 OR2X2_55 ( .gnd(gnd), .vdd(vdd), .A(_7226_), .B(_7225_), .Y(_7227_) );
NAND2X1 NAND2X1_932 ( .gnd(gnd), .vdd(vdd), .A(_7225_), .B(_7226_), .Y(_7228_) );
NAND2X1 NAND2X1_933 ( .gnd(gnd), .vdd(vdd), .A(_7228_), .B(_7227_), .Y(_7229_) );
OAI21X1 OAI21X1_2017 ( .gnd(gnd), .vdd(vdd), .A(_5093__bF_buf0), .B(_7229_), .C(_7223_), .Y(_7230_) );
XNOR2X1 XNOR2X1_279 ( .gnd(gnd), .vdd(vdd), .A(_7067__bF_buf1), .B(_4798_), .Y(_7231_) );
AOI21X1 AOI21X1_1230 ( .gnd(gnd), .vdd(vdd), .A(_6973_), .B(_6972_), .C(_6974_), .Y(_7232_) );
AND2X2 AND2X2_475 ( .gnd(gnd), .vdd(vdd), .A(_7231_), .B(_7232_), .Y(_7233_) );
NOR2X1 NOR2X1_1250 ( .gnd(gnd), .vdd(vdd), .A(_7232_), .B(_7231_), .Y(_7234_) );
OAI21X1 OAI21X1_2018 ( .gnd(gnd), .vdd(vdd), .A(_7233_), .B(_7234_), .C(micro_hash_ucr_2_pipe52_bF_buf2), .Y(_7235_) );
OAI21X1 OAI21X1_2019 ( .gnd(gnd), .vdd(vdd), .A(_7230_), .B(micro_hash_ucr_2_pipe52_bF_buf1), .C(_7235_), .Y(_7236_) );
NAND2X1 NAND2X1_934 ( .gnd(gnd), .vdd(vdd), .A(_5086__bF_buf2), .B(_7236_), .Y(_7237_) );
XNOR2X1 XNOR2X1_280 ( .gnd(gnd), .vdd(vdd), .A(_7067__bF_buf0), .B(micro_hash_ucr_2_Wx_188_), .Y(_7238_) );
INVX1 INVX1_514 ( .gnd(gnd), .vdd(vdd), .A(_7238_), .Y(_7239_) );
AOI21X1 AOI21X1_1231 ( .gnd(gnd), .vdd(vdd), .A(_6981_), .B(_6980_), .C(_6983_), .Y(_7240_) );
AND2X2 AND2X2_476 ( .gnd(gnd), .vdd(vdd), .A(_7240_), .B(_7239_), .Y(_7241_) );
NOR2X1 NOR2X1_1251 ( .gnd(gnd), .vdd(vdd), .A(_7239_), .B(_7240_), .Y(_7242_) );
OAI21X1 OAI21X1_2020 ( .gnd(gnd), .vdd(vdd), .A(_7241_), .B(_7242_), .C(micro_hash_ucr_2_pipe54_bF_buf2), .Y(_7243_) );
AND2X2 AND2X2_477 ( .gnd(gnd), .vdd(vdd), .A(_7243_), .B(_5087__bF_buf2), .Y(_7244_) );
XNOR2X1 XNOR2X1_281 ( .gnd(gnd), .vdd(vdd), .A(_7067__bF_buf5), .B(micro_hash_ucr_2_Wx_196_), .Y(_7245_) );
INVX1 INVX1_515 ( .gnd(gnd), .vdd(vdd), .A(_7245_), .Y(_7246_) );
AOI21X1 AOI21X1_1232 ( .gnd(gnd), .vdd(vdd), .A(_6989_), .B(_6988_), .C(_6990_), .Y(_7247_) );
NOR2X1 NOR2X1_1252 ( .gnd(gnd), .vdd(vdd), .A(_7247_), .B(_7246_), .Y(_7248_) );
INVX1 INVX1_516 ( .gnd(gnd), .vdd(vdd), .A(_7248_), .Y(_7249_) );
AOI21X1 AOI21X1_1233 ( .gnd(gnd), .vdd(vdd), .A(_7247_), .B(_7246_), .C(_5087__bF_buf1), .Y(_7250_) );
AOI22X1 AOI22X1_56 ( .gnd(gnd), .vdd(vdd), .A(_7249_), .B(_7250_), .C(_7237_), .D(_7244_), .Y(_7251_) );
XNOR2X1 XNOR2X1_282 ( .gnd(gnd), .vdd(vdd), .A(_7067__bF_buf4), .B(micro_hash_ucr_2_Wx_204_), .Y(_7252_) );
INVX1 INVX1_517 ( .gnd(gnd), .vdd(vdd), .A(_7252_), .Y(_7253_) );
AOI21X1 AOI21X1_1234 ( .gnd(gnd), .vdd(vdd), .A(_6997_), .B(_6996_), .C(_6998_), .Y(_7254_) );
NAND2X1 NAND2X1_935 ( .gnd(gnd), .vdd(vdd), .A(_7253_), .B(_7254_), .Y(_7255_) );
NOR2X1 NOR2X1_1253 ( .gnd(gnd), .vdd(vdd), .A(_7253_), .B(_7254_), .Y(_7256_) );
NOR2X1 NOR2X1_1254 ( .gnd(gnd), .vdd(vdd), .A(_5085__bF_buf0), .B(_7256_), .Y(_7257_) );
AOI21X1 AOI21X1_1235 ( .gnd(gnd), .vdd(vdd), .A(_7255_), .B(_7257_), .C(micro_hash_ucr_2_pipe60_bF_buf1), .Y(_7258_) );
OAI21X1 OAI21X1_2021 ( .gnd(gnd), .vdd(vdd), .A(_7251_), .B(micro_hash_ucr_2_pipe58_bF_buf4), .C(_7258_), .Y(_7259_) );
XOR2X1 XOR2X1_125 ( .gnd(gnd), .vdd(vdd), .A(_7067__bF_buf3), .B(micro_hash_ucr_2_Wx_212_), .Y(_7260_) );
AOI21X1 AOI21X1_1236 ( .gnd(gnd), .vdd(vdd), .A(_7006_), .B(_7005_), .C(_7007_), .Y(_7261_) );
AND2X2 AND2X2_478 ( .gnd(gnd), .vdd(vdd), .A(_7261_), .B(_7260_), .Y(_7262_) );
NOR2X1 NOR2X1_1255 ( .gnd(gnd), .vdd(vdd), .A(_7260_), .B(_7261_), .Y(_7263_) );
OAI21X1 OAI21X1_2022 ( .gnd(gnd), .vdd(vdd), .A(_7262_), .B(_7263_), .C(micro_hash_ucr_2_pipe60_bF_buf0), .Y(_7264_) );
NAND3X1 NAND3X1_319 ( .gnd(gnd), .vdd(vdd), .A(_5081__bF_buf0), .B(_7264_), .C(_7259_), .Y(_7265_) );
XNOR2X1 XNOR2X1_283 ( .gnd(gnd), .vdd(vdd), .A(_7067__bF_buf2), .B(micro_hash_ucr_2_Wx_220_), .Y(_7266_) );
INVX1 INVX1_518 ( .gnd(gnd), .vdd(vdd), .A(_7266_), .Y(_7267_) );
AOI21X1 AOI21X1_1237 ( .gnd(gnd), .vdd(vdd), .A(_7014_), .B(_7013_), .C(_7016_), .Y(_7268_) );
NOR2X1 NOR2X1_1256 ( .gnd(gnd), .vdd(vdd), .A(_7268_), .B(_7267_), .Y(_7269_) );
NAND2X1 NAND2X1_936 ( .gnd(gnd), .vdd(vdd), .A(_7268_), .B(_7267_), .Y(_7270_) );
NAND2X1 NAND2X1_937 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe62_bF_buf4), .B(_7270_), .Y(_7271_) );
OAI21X1 OAI21X1_2023 ( .gnd(gnd), .vdd(vdd), .A(_7269_), .B(_7271_), .C(_7265_), .Y(_7272_) );
XNOR2X1 XNOR2X1_284 ( .gnd(gnd), .vdd(vdd), .A(_7067__bF_buf1), .B(micro_hash_ucr_2_Wx_228_), .Y(_7273_) );
INVX2 INVX2_242 ( .gnd(gnd), .vdd(vdd), .A(_7273_), .Y(_7274_) );
AOI21X1 AOI21X1_1238 ( .gnd(gnd), .vdd(vdd), .A(_7024_), .B(_7022_), .C(_7025_), .Y(_7275_) );
AND2X2 AND2X2_479 ( .gnd(gnd), .vdd(vdd), .A(_7275_), .B(_7274_), .Y(_7276_) );
OAI21X1 OAI21X1_2024 ( .gnd(gnd), .vdd(vdd), .A(_7275_), .B(_7274_), .C(micro_hash_ucr_2_pipe64_bF_buf2), .Y(_7277_) );
OAI21X1 OAI21X1_2025 ( .gnd(gnd), .vdd(vdd), .A(_7276_), .B(_7277_), .C(_5074__bF_buf2), .Y(_7278_) );
AOI21X1 AOI21X1_1239 ( .gnd(gnd), .vdd(vdd), .A(_5079__bF_buf0), .B(_7272_), .C(_7278_), .Y(_7279_) );
XNOR2X1 XNOR2X1_285 ( .gnd(gnd), .vdd(vdd), .A(_7067__bF_buf0), .B(micro_hash_ucr_2_Wx_236_), .Y(_7280_) );
INVX1 INVX1_519 ( .gnd(gnd), .vdd(vdd), .A(_7280_), .Y(_7281_) );
AOI21X1 AOI21X1_1240 ( .gnd(gnd), .vdd(vdd), .A(_7033_), .B(_7031_), .C(_7034_), .Y(_7282_) );
NAND2X1 NAND2X1_938 ( .gnd(gnd), .vdd(vdd), .A(_7282_), .B(_7281_), .Y(_7283_) );
NOR2X1 NOR2X1_1257 ( .gnd(gnd), .vdd(vdd), .A(_7282_), .B(_7281_), .Y(_7284_) );
INVX1 INVX1_520 ( .gnd(gnd), .vdd(vdd), .A(_7284_), .Y(_7285_) );
AOI21X1 AOI21X1_1241 ( .gnd(gnd), .vdd(vdd), .A(_7283_), .B(_7285_), .C(_5074__bF_buf1), .Y(_7286_) );
OAI21X1 OAI21X1_2026 ( .gnd(gnd), .vdd(vdd), .A(_7279_), .B(_7286_), .C(_5075__bF_buf0), .Y(_7287_) );
XNOR2X1 XNOR2X1_286 ( .gnd(gnd), .vdd(vdd), .A(_7067__bF_buf5), .B(micro_hash_ucr_2_Wx_244_), .Y(_7288_) );
INVX1 INVX1_521 ( .gnd(gnd), .vdd(vdd), .A(_7288_), .Y(_7289_) );
AOI21X1 AOI21X1_1242 ( .gnd(gnd), .vdd(vdd), .A(_7043_), .B(_7041_), .C(_7045_), .Y(_7290_) );
AND2X2 AND2X2_480 ( .gnd(gnd), .vdd(vdd), .A(_7290_), .B(_7289_), .Y(_7291_) );
NOR2X1 NOR2X1_1258 ( .gnd(gnd), .vdd(vdd), .A(_7289_), .B(_7290_), .Y(_7292_) );
OAI21X1 OAI21X1_2027 ( .gnd(gnd), .vdd(vdd), .A(_7291_), .B(_7292_), .C(micro_hash_ucr_2_pipe68), .Y(_7293_) );
NAND2X1 NAND2X1_939 ( .gnd(gnd), .vdd(vdd), .A(_7293_), .B(_7287_), .Y(_7294_) );
XNOR2X1 XNOR2X1_287 ( .gnd(gnd), .vdd(vdd), .A(_7067__bF_buf4), .B(micro_hash_ucr_2_Wx_252_), .Y(_7295_) );
INVX2 INVX2_243 ( .gnd(gnd), .vdd(vdd), .A(_7295_), .Y(_7296_) );
AOI21X1 AOI21X1_1243 ( .gnd(gnd), .vdd(vdd), .A(_7052_), .B(_7050_), .C(_7054_), .Y(_7297_) );
AOI21X1 AOI21X1_1244 ( .gnd(gnd), .vdd(vdd), .A(_7296_), .B(_7297_), .C(_4594__bF_buf12), .Y(_7298_) );
OAI21X1 OAI21X1_2028 ( .gnd(gnd), .vdd(vdd), .A(_7296_), .B(_7297_), .C(_7298_), .Y(_7299_) );
AOI22X1 AOI22X1_57 ( .gnd(gnd), .vdd(vdd), .A(_6147_), .B(_7299_), .C(_7294_), .D(_5073__bF_buf0), .Y(_4493__4_) );
INVX1 INVX1_522 ( .gnd(gnd), .vdd(vdd), .A(_4563_), .Y(_7300_) );
INVX8 INVX8_190 ( .gnd(gnd), .vdd(vdd), .A(_7067__bF_buf3), .Y(_7301_) );
AOI21X1 AOI21X1_1245 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_220_), .B(_7301__bF_buf3), .C(_7269_), .Y(_7302_) );
INVX1 INVX1_523 ( .gnd(gnd), .vdd(vdd), .A(_7062_), .Y(_7303_) );
OAI21X1 OAI21X1_2029 ( .gnd(gnd), .vdd(vdd), .A(_7058_), .B(_7064_), .C(_7303_), .Y(_7304_) );
INVX2 INVX2_244 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_x_5_), .Y(_7305_) );
NAND2X1 NAND2X1_940 ( .gnd(gnd), .vdd(vdd), .A(_6030_), .B(_7305_), .Y(_7306_) );
NOR2X1 NOR2X1_1259 ( .gnd(gnd), .vdd(vdd), .A(_6030_), .B(_7305_), .Y(_7307_) );
INVX1 INVX1_524 ( .gnd(gnd), .vdd(vdd), .A(_7307_), .Y(_7308_) );
AND2X2 AND2X2_481 ( .gnd(gnd), .vdd(vdd), .A(_7308_), .B(_7306_), .Y(_7309_) );
NAND2X1 NAND2X1_941 ( .gnd(gnd), .vdd(vdd), .A(_7309_), .B(_7304_), .Y(_7310_) );
INVX8 INVX8_191 ( .gnd(gnd), .vdd(vdd), .A(_7310_), .Y(_7311_) );
NOR2X1 NOR2X1_1260 ( .gnd(gnd), .vdd(vdd), .A(_7309_), .B(_7304_), .Y(_7312_) );
OAI21X1 OAI21X1_2030 ( .gnd(gnd), .vdd(vdd), .A(_7311__bF_buf3), .B(_7312_), .C(_4744_), .Y(_7313_) );
INVX1 INVX1_525 ( .gnd(gnd), .vdd(vdd), .A(_7313_), .Y(_7314_) );
NOR2X1 NOR2X1_1261 ( .gnd(gnd), .vdd(vdd), .A(_7312_), .B(_7311__bF_buf2), .Y(_7315_) );
INVX8 INVX8_192 ( .gnd(gnd), .vdd(vdd), .A(_7315__bF_buf5), .Y(_7316_) );
NOR2X1 NOR2X1_1262 ( .gnd(gnd), .vdd(vdd), .A(_4744_), .B(_7316__bF_buf3), .Y(_7317_) );
NOR2X1 NOR2X1_1263 ( .gnd(gnd), .vdd(vdd), .A(_7314_), .B(_7317_), .Y(_7318_) );
XNOR2X1 XNOR2X1_288 ( .gnd(gnd), .vdd(vdd), .A(_7302_), .B(_7318_), .Y(_7319_) );
AOI21X1 AOI21X1_1246 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_188_), .B(_7301__bF_buf2), .C(_7242_), .Y(_7320_) );
OAI21X1 OAI21X1_2031 ( .gnd(gnd), .vdd(vdd), .A(_7311__bF_buf1), .B(_7312_), .C(_4859_), .Y(_7321_) );
INVX1 INVX1_526 ( .gnd(gnd), .vdd(vdd), .A(_7321_), .Y(_7322_) );
NOR2X1 NOR2X1_1264 ( .gnd(gnd), .vdd(vdd), .A(_4859_), .B(_7316__bF_buf2), .Y(_7323_) );
NOR2X1 NOR2X1_1265 ( .gnd(gnd), .vdd(vdd), .A(_7322_), .B(_7323_), .Y(_7324_) );
XNOR2X1 XNOR2X1_289 ( .gnd(gnd), .vdd(vdd), .A(_7320_), .B(_7324_), .Y(_7325_) );
AOI21X1 AOI21X1_1247 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_4_), .B(_7301__bF_buf1), .C(_7072_), .Y(_7326_) );
XNOR2X1 XNOR2X1_290 ( .gnd(gnd), .vdd(vdd), .A(_7315__bF_buf4), .B(micro_hash_ucr_2_Wx_5_), .Y(_7327_) );
XNOR2X1 XNOR2X1_291 ( .gnd(gnd), .vdd(vdd), .A(_7326_), .B(_7327_), .Y(_7328_) );
NOR2X1 NOR2X1_1266 ( .gnd(gnd), .vdd(vdd), .A(_8668_), .B(_5134_), .Y(_7329_) );
OAI21X1 OAI21X1_2032 ( .gnd(gnd), .vdd(vdd), .A(_8669_), .B(micro_hash_ucr_2_pipe6), .C(_5135_), .Y(_7330_) );
OAI21X1 OAI21X1_2033 ( .gnd(gnd), .vdd(vdd), .A(_7330_), .B(_7329_), .C(_5133_), .Y(_7331_) );
AOI21X1 AOI21X1_1248 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe8), .B(_7328_), .C(_7331_), .Y(_7332_) );
INVX1 INVX1_527 ( .gnd(gnd), .vdd(vdd), .A(_7076_), .Y(_7333_) );
NOR2X1 NOR2X1_1267 ( .gnd(gnd), .vdd(vdd), .A(_7074_), .B(_7333_), .Y(_7334_) );
AOI21X1 AOI21X1_1249 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_12_), .B(_7301__bF_buf0), .C(_7334_), .Y(_7335_) );
NOR2X1 NOR2X1_1268 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_13_), .B(_7315__bF_buf3), .Y(_7336_) );
INVX1 INVX1_528 ( .gnd(gnd), .vdd(vdd), .A(_7336_), .Y(_7337_) );
NAND2X1 NAND2X1_942 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_13_), .B(_7315__bF_buf2), .Y(_7338_) );
NAND2X1 NAND2X1_943 ( .gnd(gnd), .vdd(vdd), .A(_7338_), .B(_7337_), .Y(_7339_) );
XNOR2X1 XNOR2X1_292 ( .gnd(gnd), .vdd(vdd), .A(_7335_), .B(_7339_), .Y(_7340_) );
OAI21X1 OAI21X1_2034 ( .gnd(gnd), .vdd(vdd), .A(_7340_), .B(_5133_), .C(_5128_), .Y(_7341_) );
OAI21X1 OAI21X1_2035 ( .gnd(gnd), .vdd(vdd), .A(_7082_), .B(_7067__bF_buf2), .C(_7087_), .Y(_7342_) );
NOR2X1 NOR2X1_1269 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_21_), .B(_7315__bF_buf1), .Y(_7343_) );
INVX1 INVX1_529 ( .gnd(gnd), .vdd(vdd), .A(_7343_), .Y(_7344_) );
NAND2X1 NAND2X1_944 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_21_), .B(_7315__bF_buf0), .Y(_7345_) );
NAND2X1 NAND2X1_945 ( .gnd(gnd), .vdd(vdd), .A(_7345_), .B(_7344_), .Y(_7346_) );
AOI21X1 AOI21X1_1250 ( .gnd(gnd), .vdd(vdd), .A(_7346_), .B(_7342_), .C(_5128_), .Y(_7347_) );
OAI21X1 OAI21X1_2036 ( .gnd(gnd), .vdd(vdd), .A(_7342_), .B(_7346_), .C(_7347_), .Y(_7348_) );
OAI21X1 OAI21X1_2037 ( .gnd(gnd), .vdd(vdd), .A(_7332_), .B(_7341_), .C(_7348_), .Y(_7349_) );
NAND2X1 NAND2X1_946 ( .gnd(gnd), .vdd(vdd), .A(_5129_), .B(_7349_), .Y(_7350_) );
AOI21X1 AOI21X1_1251 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_28_), .B(_7301__bF_buf3), .C(_7092_), .Y(_7351_) );
NOR2X1 NOR2X1_1270 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_29_), .B(_7315__bF_buf5), .Y(_7352_) );
INVX1 INVX1_530 ( .gnd(gnd), .vdd(vdd), .A(_7352_), .Y(_7353_) );
NAND2X1 NAND2X1_947 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_29_), .B(_7315__bF_buf4), .Y(_7354_) );
NAND2X1 NAND2X1_948 ( .gnd(gnd), .vdd(vdd), .A(_7354_), .B(_7353_), .Y(_7355_) );
XOR2X1 XOR2X1_126 ( .gnd(gnd), .vdd(vdd), .A(_7355_), .B(_7351_), .Y(_7356_) );
OAI21X1 OAI21X1_2038 ( .gnd(gnd), .vdd(vdd), .A(_5129_), .B(_7356_), .C(_7350_), .Y(_7357_) );
NAND2X1 NAND2X1_949 ( .gnd(gnd), .vdd(vdd), .A(_5127__bF_buf1), .B(_7357_), .Y(_7358_) );
AOI21X1 AOI21X1_1252 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_36_), .B(_7301__bF_buf2), .C(_7100_), .Y(_7359_) );
INVX2 INVX2_245 ( .gnd(gnd), .vdd(vdd), .A(_7359_), .Y(_7360_) );
INVX1 INVX1_531 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_37_), .Y(_7361_) );
OAI21X1 OAI21X1_2039 ( .gnd(gnd), .vdd(vdd), .A(_7311__bF_buf0), .B(_7312_), .C(_7361_), .Y(_7362_) );
NOR2X1 NOR2X1_1271 ( .gnd(gnd), .vdd(vdd), .A(_7361_), .B(_7316__bF_buf1), .Y(_7363_) );
INVX1 INVX1_532 ( .gnd(gnd), .vdd(vdd), .A(_7363_), .Y(_7364_) );
NAND2X1 NAND2X1_950 ( .gnd(gnd), .vdd(vdd), .A(_7362_), .B(_7364_), .Y(_7365_) );
AOI21X1 AOI21X1_1253 ( .gnd(gnd), .vdd(vdd), .A(_7365_), .B(_7360_), .C(_5127__bF_buf0), .Y(_7366_) );
OAI21X1 OAI21X1_2040 ( .gnd(gnd), .vdd(vdd), .A(_7360_), .B(_7365_), .C(_7366_), .Y(_7367_) );
AND2X2 AND2X2_482 ( .gnd(gnd), .vdd(vdd), .A(_7367_), .B(_5122__bF_buf3), .Y(_7368_) );
AOI21X1 AOI21X1_1254 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_44_), .B(_7301__bF_buf1), .C(_7106_), .Y(_7369_) );
NOR2X1 NOR2X1_1272 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_45_), .B(_7315__bF_buf3), .Y(_7370_) );
INVX1 INVX1_533 ( .gnd(gnd), .vdd(vdd), .A(_7370_), .Y(_7371_) );
NAND2X1 NAND2X1_951 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_45_), .B(_7315__bF_buf2), .Y(_7372_) );
NAND2X1 NAND2X1_952 ( .gnd(gnd), .vdd(vdd), .A(_7372_), .B(_7371_), .Y(_7373_) );
AND2X2 AND2X2_483 ( .gnd(gnd), .vdd(vdd), .A(_7369_), .B(_7373_), .Y(_7374_) );
OAI21X1 OAI21X1_2041 ( .gnd(gnd), .vdd(vdd), .A(_7369_), .B(_7373_), .C(micro_hash_ucr_2_pipe18_bF_buf1), .Y(_7375_) );
OAI21X1 OAI21X1_2042 ( .gnd(gnd), .vdd(vdd), .A(_7374_), .B(_7375_), .C(_5123__bF_buf3), .Y(_7376_) );
AOI21X1 AOI21X1_1255 ( .gnd(gnd), .vdd(vdd), .A(_7368_), .B(_7358_), .C(_7376_), .Y(_7377_) );
AOI21X1 AOI21X1_1256 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_52_), .B(_7301__bF_buf0), .C(_7114_), .Y(_7378_) );
NOR2X1 NOR2X1_1273 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_53_), .B(_7315__bF_buf1), .Y(_7379_) );
INVX1 INVX1_534 ( .gnd(gnd), .vdd(vdd), .A(_7379_), .Y(_7380_) );
NAND2X1 NAND2X1_953 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_53_), .B(_7315__bF_buf0), .Y(_7381_) );
NAND2X1 NAND2X1_954 ( .gnd(gnd), .vdd(vdd), .A(_7381_), .B(_7380_), .Y(_7382_) );
XOR2X1 XOR2X1_127 ( .gnd(gnd), .vdd(vdd), .A(_7378_), .B(_7382_), .Y(_7383_) );
OAI21X1 OAI21X1_2043 ( .gnd(gnd), .vdd(vdd), .A(_7383_), .B(_5123__bF_buf2), .C(_5121__bF_buf2), .Y(_7384_) );
OAI21X1 OAI21X1_2044 ( .gnd(gnd), .vdd(vdd), .A(_5016_), .B(_7067__bF_buf1), .C(_7123_), .Y(_7385_) );
XNOR2X1 XNOR2X1_293 ( .gnd(gnd), .vdd(vdd), .A(_7315__bF_buf5), .B(micro_hash_ucr_2_Wx_61_), .Y(_7386_) );
XNOR2X1 XNOR2X1_294 ( .gnd(gnd), .vdd(vdd), .A(_7385_), .B(_7386_), .Y(_7387_) );
AOI21X1 AOI21X1_1257 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe22_bF_buf2), .B(_7387_), .C(micro_hash_ucr_2_pipe24_bF_buf2), .Y(_7388_) );
OAI21X1 OAI21X1_2045 ( .gnd(gnd), .vdd(vdd), .A(_7377_), .B(_7384_), .C(_7388_), .Y(_7389_) );
INVX1 INVX1_535 ( .gnd(gnd), .vdd(vdd), .A(_7128_), .Y(_7390_) );
NAND2X1 NAND2X1_955 ( .gnd(gnd), .vdd(vdd), .A(_7127_), .B(_7390_), .Y(_7391_) );
OAI21X1 OAI21X1_2046 ( .gnd(gnd), .vdd(vdd), .A(_5062_), .B(_7067__bF_buf0), .C(_7391_), .Y(_7392_) );
OAI21X1 OAI21X1_2047 ( .gnd(gnd), .vdd(vdd), .A(_7311__bF_buf3), .B(_7312_), .C(_5065_), .Y(_7393_) );
NOR2X1 NOR2X1_1274 ( .gnd(gnd), .vdd(vdd), .A(_5065_), .B(_7316__bF_buf0), .Y(_7394_) );
INVX1 INVX1_536 ( .gnd(gnd), .vdd(vdd), .A(_7394_), .Y(_7395_) );
NAND2X1 NAND2X1_956 ( .gnd(gnd), .vdd(vdd), .A(_7393_), .B(_7395_), .Y(_7396_) );
AOI21X1 AOI21X1_1258 ( .gnd(gnd), .vdd(vdd), .A(_7392_), .B(_7396_), .C(_5116__bF_buf3), .Y(_7397_) );
OAI21X1 OAI21X1_2048 ( .gnd(gnd), .vdd(vdd), .A(_7392_), .B(_7396_), .C(_7397_), .Y(_7398_) );
AND2X2 AND2X2_484 ( .gnd(gnd), .vdd(vdd), .A(_7398_), .B(_5117__bF_buf4), .Y(_7399_) );
AOI21X1 AOI21X1_1259 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_76_), .B(_7301__bF_buf3), .C(_7133_), .Y(_7400_) );
OAI21X1 OAI21X1_2049 ( .gnd(gnd), .vdd(vdd), .A(_7311__bF_buf2), .B(_7312_), .C(_5041_), .Y(_7401_) );
NAND2X1 NAND2X1_957 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_77_), .B(_7315__bF_buf4), .Y(_7402_) );
NAND2X1 NAND2X1_958 ( .gnd(gnd), .vdd(vdd), .A(_7401_), .B(_7402_), .Y(_7403_) );
AND2X2 AND2X2_485 ( .gnd(gnd), .vdd(vdd), .A(_7400_), .B(_7403_), .Y(_7404_) );
OAI21X1 OAI21X1_2050 ( .gnd(gnd), .vdd(vdd), .A(_7400_), .B(_7403_), .C(micro_hash_ucr_2_pipe26_bF_buf2), .Y(_7405_) );
OAI21X1 OAI21X1_2051 ( .gnd(gnd), .vdd(vdd), .A(_7404_), .B(_7405_), .C(_5115__bF_buf1), .Y(_7406_) );
AOI21X1 AOI21X1_1260 ( .gnd(gnd), .vdd(vdd), .A(_7399_), .B(_7389_), .C(_7406_), .Y(_7407_) );
OAI21X1 OAI21X1_2052 ( .gnd(gnd), .vdd(vdd), .A(_4947_), .B(_7067__bF_buf5), .C(_7142_), .Y(_7408_) );
XNOR2X1 XNOR2X1_295 ( .gnd(gnd), .vdd(vdd), .A(_7315__bF_buf3), .B(micro_hash_ucr_2_Wx_85_), .Y(_7409_) );
XNOR2X1 XNOR2X1_296 ( .gnd(gnd), .vdd(vdd), .A(_7408_), .B(_7409_), .Y(_7410_) );
OAI21X1 OAI21X1_2053 ( .gnd(gnd), .vdd(vdd), .A(_7410_), .B(_5115__bF_buf0), .C(_5110__bF_buf3), .Y(_7411_) );
OAI21X1 OAI21X1_2054 ( .gnd(gnd), .vdd(vdd), .A(_4991_), .B(_7067__bF_buf4), .C(_7149_), .Y(_7412_) );
OAI21X1 OAI21X1_2055 ( .gnd(gnd), .vdd(vdd), .A(_7311__bF_buf1), .B(_7312_), .C(_4994_), .Y(_7413_) );
INVX1 INVX1_537 ( .gnd(gnd), .vdd(vdd), .A(_7413_), .Y(_7414_) );
NOR2X1 NOR2X1_1275 ( .gnd(gnd), .vdd(vdd), .A(_4994_), .B(_7316__bF_buf3), .Y(_7415_) );
NOR2X1 NOR2X1_1276 ( .gnd(gnd), .vdd(vdd), .A(_7414_), .B(_7415_), .Y(_7416_) );
XOR2X1 XOR2X1_128 ( .gnd(gnd), .vdd(vdd), .A(_7412_), .B(_7416_), .Y(_7417_) );
AOI21X1 AOI21X1_1261 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe30_bF_buf3), .B(_7417_), .C(micro_hash_ucr_2_pipe32_bF_buf3), .Y(_7418_) );
OAI21X1 OAI21X1_2056 ( .gnd(gnd), .vdd(vdd), .A(_7407_), .B(_7411_), .C(_7418_), .Y(_7419_) );
AOI21X1 AOI21X1_1262 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_100_), .B(_7301__bF_buf2), .C(_7157_), .Y(_7420_) );
XNOR2X1 XNOR2X1_297 ( .gnd(gnd), .vdd(vdd), .A(_7315__bF_buf2), .B(micro_hash_ucr_2_Wx_101_), .Y(_7421_) );
XNOR2X1 XNOR2X1_298 ( .gnd(gnd), .vdd(vdd), .A(_7420_), .B(_7421_), .Y(_7422_) );
AOI21X1 AOI21X1_1263 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe32_bF_buf2), .B(_7422_), .C(micro_hash_ucr_2_pipe34_bF_buf1), .Y(_7423_) );
OAI21X1 OAI21X1_2057 ( .gnd(gnd), .vdd(vdd), .A(_4881_), .B(_7067__bF_buf3), .C(_7165_), .Y(_7424_) );
OAI21X1 OAI21X1_2058 ( .gnd(gnd), .vdd(vdd), .A(_7311__bF_buf0), .B(_7312_), .C(_4884_), .Y(_7425_) );
NOR2X1 NOR2X1_1277 ( .gnd(gnd), .vdd(vdd), .A(_4884_), .B(_7316__bF_buf2), .Y(_7426_) );
INVX1 INVX1_538 ( .gnd(gnd), .vdd(vdd), .A(_7426_), .Y(_7427_) );
NAND2X1 NAND2X1_959 ( .gnd(gnd), .vdd(vdd), .A(_7425_), .B(_7427_), .Y(_7428_) );
XOR2X1 XOR2X1_129 ( .gnd(gnd), .vdd(vdd), .A(_7424_), .B(_7428_), .Y(_7429_) );
OAI21X1 OAI21X1_2059 ( .gnd(gnd), .vdd(vdd), .A(_7429_), .B(_5109__bF_buf1), .C(_5104__bF_buf1), .Y(_7430_) );
AOI21X1 AOI21X1_1264 ( .gnd(gnd), .vdd(vdd), .A(_7423_), .B(_7419_), .C(_7430_), .Y(_7431_) );
OAI21X1 OAI21X1_2060 ( .gnd(gnd), .vdd(vdd), .A(_4925_), .B(_7067__bF_buf2), .C(_7172_), .Y(_7432_) );
OAI21X1 OAI21X1_2061 ( .gnd(gnd), .vdd(vdd), .A(_7311__bF_buf3), .B(_7312_), .C(_4928_), .Y(_7433_) );
NOR2X1 NOR2X1_1278 ( .gnd(gnd), .vdd(vdd), .A(_4928_), .B(_7316__bF_buf1), .Y(_7434_) );
INVX1 INVX1_539 ( .gnd(gnd), .vdd(vdd), .A(_7434_), .Y(_7435_) );
NAND2X1 NAND2X1_960 ( .gnd(gnd), .vdd(vdd), .A(_7433_), .B(_7435_), .Y(_7436_) );
XNOR2X1 XNOR2X1_299 ( .gnd(gnd), .vdd(vdd), .A(_7432_), .B(_7436_), .Y(_7437_) );
OAI21X1 OAI21X1_2062 ( .gnd(gnd), .vdd(vdd), .A(_7437_), .B(_5104__bF_buf0), .C(_5105__bF_buf4), .Y(_7438_) );
OAI21X1 OAI21X1_2063 ( .gnd(gnd), .vdd(vdd), .A(_4768_), .B(_7067__bF_buf1), .C(_7180_), .Y(_7439_) );
XNOR2X1 XNOR2X1_300 ( .gnd(gnd), .vdd(vdd), .A(_7315__bF_buf1), .B(micro_hash_ucr_2_Wx_125_), .Y(_7440_) );
XNOR2X1 XNOR2X1_301 ( .gnd(gnd), .vdd(vdd), .A(_7439_), .B(_7440_), .Y(_7441_) );
AOI21X1 AOI21X1_1265 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe38_bF_buf2), .B(_7441_), .C(micro_hash_ucr_2_pipe40_bF_buf1), .Y(_7442_) );
OAI21X1 OAI21X1_2064 ( .gnd(gnd), .vdd(vdd), .A(_7431_), .B(_7438_), .C(_7442_), .Y(_7443_) );
OAI21X1 OAI21X1_2065 ( .gnd(gnd), .vdd(vdd), .A(_4797_), .B(_7067__bF_buf0), .C(_7190_), .Y(_7444_) );
OAI21X1 OAI21X1_2066 ( .gnd(gnd), .vdd(vdd), .A(_7311__bF_buf2), .B(_7312_), .C(_4801_), .Y(_7445_) );
NOR2X1 NOR2X1_1279 ( .gnd(gnd), .vdd(vdd), .A(_4801_), .B(_7316__bF_buf0), .Y(_7446_) );
INVX1 INVX1_540 ( .gnd(gnd), .vdd(vdd), .A(_7446_), .Y(_7447_) );
NAND2X1 NAND2X1_961 ( .gnd(gnd), .vdd(vdd), .A(_7445_), .B(_7447_), .Y(_7448_) );
AOI21X1 AOI21X1_1266 ( .gnd(gnd), .vdd(vdd), .A(_7448_), .B(_7444_), .C(_5103__bF_buf1), .Y(_7449_) );
OAI21X1 OAI21X1_2067 ( .gnd(gnd), .vdd(vdd), .A(_7444_), .B(_7448_), .C(_7449_), .Y(_7450_) );
AND2X2 AND2X2_486 ( .gnd(gnd), .vdd(vdd), .A(_7450_), .B(_5098__bF_buf1), .Y(_7451_) );
AOI21X1 AOI21X1_1267 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_140_), .B(_7301__bF_buf1), .C(_7197_), .Y(_7452_) );
OAI21X1 OAI21X1_2068 ( .gnd(gnd), .vdd(vdd), .A(_7311__bF_buf1), .B(_7312_), .C(_4995_), .Y(_7453_) );
NAND2X1 NAND2X1_962 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_141_), .B(_7315__bF_buf0), .Y(_7454_) );
NAND2X1 NAND2X1_963 ( .gnd(gnd), .vdd(vdd), .A(_7453_), .B(_7454_), .Y(_7455_) );
AND2X2 AND2X2_487 ( .gnd(gnd), .vdd(vdd), .A(_7452_), .B(_7455_), .Y(_7456_) );
OAI21X1 OAI21X1_2069 ( .gnd(gnd), .vdd(vdd), .A(_7452_), .B(_7455_), .C(micro_hash_ucr_2_pipe42_bF_buf0), .Y(_7457_) );
OAI21X1 OAI21X1_2070 ( .gnd(gnd), .vdd(vdd), .A(_7456_), .B(_7457_), .C(_5099__bF_buf2), .Y(_7458_) );
AOI21X1 AOI21X1_1268 ( .gnd(gnd), .vdd(vdd), .A(_7451_), .B(_7443_), .C(_7458_), .Y(_7459_) );
OAI21X1 OAI21X1_2071 ( .gnd(gnd), .vdd(vdd), .A(_4827_), .B(_7067__bF_buf5), .C(_7204_), .Y(_7460_) );
OAI21X1 OAI21X1_2072 ( .gnd(gnd), .vdd(vdd), .A(_7311__bF_buf0), .B(_7312_), .C(_4830_), .Y(_7461_) );
NOR2X1 NOR2X1_1280 ( .gnd(gnd), .vdd(vdd), .A(_4830_), .B(_7316__bF_buf3), .Y(_7462_) );
INVX1 INVX1_541 ( .gnd(gnd), .vdd(vdd), .A(_7462_), .Y(_7463_) );
NAND2X1 NAND2X1_964 ( .gnd(gnd), .vdd(vdd), .A(_7461_), .B(_7463_), .Y(_7464_) );
AOI21X1 AOI21X1_1269 ( .gnd(gnd), .vdd(vdd), .A(_7464_), .B(_7460_), .C(_5099__bF_buf1), .Y(_7465_) );
OAI21X1 OAI21X1_2073 ( .gnd(gnd), .vdd(vdd), .A(_7460_), .B(_7464_), .C(_7465_), .Y(_7466_) );
NAND2X1 NAND2X1_965 ( .gnd(gnd), .vdd(vdd), .A(_5097__bF_buf0), .B(_7466_), .Y(_7467_) );
OAI21X1 OAI21X1_2074 ( .gnd(gnd), .vdd(vdd), .A(_4713_), .B(_7067__bF_buf4), .C(_7214_), .Y(_7468_) );
XNOR2X1 XNOR2X1_302 ( .gnd(gnd), .vdd(vdd), .A(_7315__bF_buf5), .B(micro_hash_ucr_2_Wx_157_), .Y(_7469_) );
XNOR2X1 XNOR2X1_303 ( .gnd(gnd), .vdd(vdd), .A(_7468_), .B(_7469_), .Y(_7470_) );
AOI21X1 AOI21X1_1270 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe46_bF_buf2), .B(_7470_), .C(micro_hash_ucr_2_pipe48_bF_buf4), .Y(_7471_) );
OAI21X1 OAI21X1_2075 ( .gnd(gnd), .vdd(vdd), .A(_7459_), .B(_7467_), .C(_7471_), .Y(_7472_) );
AOI21X1 AOI21X1_1271 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_164_), .B(_7301__bF_buf0), .C(_7221_), .Y(_7473_) );
OAI21X1 OAI21X1_2076 ( .gnd(gnd), .vdd(vdd), .A(_7311__bF_buf3), .B(_7312_), .C(_4771_), .Y(_7474_) );
NAND2X1 NAND2X1_966 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_165_), .B(_7315__bF_buf4), .Y(_7475_) );
NAND2X1 NAND2X1_967 ( .gnd(gnd), .vdd(vdd), .A(_7474_), .B(_7475_), .Y(_7476_) );
XNOR2X1 XNOR2X1_304 ( .gnd(gnd), .vdd(vdd), .A(_7473_), .B(_7476_), .Y(_7477_) );
AOI21X1 AOI21X1_1272 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe48_bF_buf3), .B(_7477_), .C(micro_hash_ucr_2_pipe50_bF_buf2), .Y(_7478_) );
OAI21X1 OAI21X1_2077 ( .gnd(gnd), .vdd(vdd), .A(_4740_), .B(_7067__bF_buf3), .C(_7227_), .Y(_7479_) );
OAI21X1 OAI21X1_2078 ( .gnd(gnd), .vdd(vdd), .A(_7311__bF_buf2), .B(_7312_), .C(_4743_), .Y(_7480_) );
NOR2X1 NOR2X1_1281 ( .gnd(gnd), .vdd(vdd), .A(_4743_), .B(_7316__bF_buf2), .Y(_7481_) );
INVX1 INVX1_542 ( .gnd(gnd), .vdd(vdd), .A(_7481_), .Y(_7482_) );
NAND2X1 NAND2X1_968 ( .gnd(gnd), .vdd(vdd), .A(_7480_), .B(_7482_), .Y(_7483_) );
XOR2X1 XOR2X1_130 ( .gnd(gnd), .vdd(vdd), .A(_7483_), .B(_7479_), .Y(_7484_) );
OAI21X1 OAI21X1_2079 ( .gnd(gnd), .vdd(vdd), .A(_7484_), .B(_5093__bF_buf4), .C(_5091__bF_buf1), .Y(_7485_) );
AOI21X1 AOI21X1_1273 ( .gnd(gnd), .vdd(vdd), .A(_7478_), .B(_7472_), .C(_7485_), .Y(_7486_) );
AOI21X1 AOI21X1_1274 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_180_), .B(_7301__bF_buf3), .C(_7234_), .Y(_7487_) );
NOR2X1 NOR2X1_1282 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_181_), .B(_7315__bF_buf3), .Y(_7488_) );
NOR2X1 NOR2X1_1283 ( .gnd(gnd), .vdd(vdd), .A(_4802_), .B(_7316__bF_buf1), .Y(_7489_) );
NOR2X1 NOR2X1_1284 ( .gnd(gnd), .vdd(vdd), .A(_7488_), .B(_7489_), .Y(_7490_) );
OAI21X1 OAI21X1_2080 ( .gnd(gnd), .vdd(vdd), .A(_7490_), .B(_7487_), .C(micro_hash_ucr_2_pipe52_bF_buf0), .Y(_7491_) );
AOI21X1 AOI21X1_1275 ( .gnd(gnd), .vdd(vdd), .A(_7487_), .B(_7490_), .C(_7491_), .Y(_7492_) );
OAI21X1 OAI21X1_2081 ( .gnd(gnd), .vdd(vdd), .A(_7486_), .B(_7492_), .C(_5086__bF_buf1), .Y(_7493_) );
OAI21X1 OAI21X1_2082 ( .gnd(gnd), .vdd(vdd), .A(_5086__bF_buf0), .B(_7325_), .C(_7493_), .Y(_7494_) );
NAND2X1 NAND2X1_969 ( .gnd(gnd), .vdd(vdd), .A(_5087__bF_buf0), .B(_7494_), .Y(_7495_) );
AOI21X1 AOI21X1_1276 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_196_), .B(_7301__bF_buf2), .C(_7248_), .Y(_7496_) );
NOR2X1 NOR2X1_1285 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_197_), .B(_7315__bF_buf2), .Y(_7497_) );
INVX1 INVX1_543 ( .gnd(gnd), .vdd(vdd), .A(_7497_), .Y(_7498_) );
NAND2X1 NAND2X1_970 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_197_), .B(_7315__bF_buf1), .Y(_7499_) );
NAND2X1 NAND2X1_971 ( .gnd(gnd), .vdd(vdd), .A(_7499_), .B(_7498_), .Y(_7500_) );
XNOR2X1 XNOR2X1_305 ( .gnd(gnd), .vdd(vdd), .A(_7496_), .B(_7500_), .Y(_7501_) );
AOI21X1 AOI21X1_1277 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe56_bF_buf1), .B(_7501_), .C(micro_hash_ucr_2_pipe58_bF_buf3), .Y(_7502_) );
AOI21X1 AOI21X1_1278 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_204_), .B(_7301__bF_buf1), .C(_7256_), .Y(_7503_) );
NOR2X1 NOR2X1_1286 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_205_), .B(_7315__bF_buf0), .Y(_7504_) );
INVX1 INVX1_544 ( .gnd(gnd), .vdd(vdd), .A(_7504_), .Y(_7505_) );
NAND2X1 NAND2X1_972 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_205_), .B(_7315__bF_buf5), .Y(_7506_) );
NAND2X1 NAND2X1_973 ( .gnd(gnd), .vdd(vdd), .A(_7506_), .B(_7505_), .Y(_7507_) );
AND2X2 AND2X2_488 ( .gnd(gnd), .vdd(vdd), .A(_7503_), .B(_7507_), .Y(_7508_) );
OAI21X1 OAI21X1_2083 ( .gnd(gnd), .vdd(vdd), .A(_7503_), .B(_7507_), .C(micro_hash_ucr_2_pipe58_bF_buf2), .Y(_7509_) );
OAI21X1 OAI21X1_2084 ( .gnd(gnd), .vdd(vdd), .A(_7508_), .B(_7509_), .C(_5080__bF_buf2), .Y(_7510_) );
AOI21X1 AOI21X1_1279 ( .gnd(gnd), .vdd(vdd), .A(_7502_), .B(_7495_), .C(_7510_), .Y(_7511_) );
AOI21X1 AOI21X1_1280 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_212_), .B(_7301__bF_buf0), .C(_7263_), .Y(_7512_) );
NOR2X1 NOR2X1_1287 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_213_), .B(_7315__bF_buf4), .Y(_7513_) );
NAND2X1 NAND2X1_974 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_213_), .B(_7315__bF_buf3), .Y(_7514_) );
INVX1 INVX1_545 ( .gnd(gnd), .vdd(vdd), .A(_7514_), .Y(_7515_) );
NOR2X1 NOR2X1_1288 ( .gnd(gnd), .vdd(vdd), .A(_7513_), .B(_7515_), .Y(_7516_) );
OAI21X1 OAI21X1_2085 ( .gnd(gnd), .vdd(vdd), .A(_7512_), .B(_7516_), .C(micro_hash_ucr_2_pipe60_bF_buf4), .Y(_7517_) );
AOI21X1 AOI21X1_1281 ( .gnd(gnd), .vdd(vdd), .A(_7512_), .B(_7516_), .C(_7517_), .Y(_7518_) );
OAI21X1 OAI21X1_2086 ( .gnd(gnd), .vdd(vdd), .A(_7511_), .B(_7518_), .C(_5081__bF_buf3), .Y(_7519_) );
OAI21X1 OAI21X1_2087 ( .gnd(gnd), .vdd(vdd), .A(_5081__bF_buf2), .B(_7319_), .C(_7519_), .Y(_7520_) );
NAND2X1 NAND2X1_975 ( .gnd(gnd), .vdd(vdd), .A(_5079__bF_buf4), .B(_7520_), .Y(_7521_) );
NOR2X1 NOR2X1_1289 ( .gnd(gnd), .vdd(vdd), .A(_7274_), .B(_7275_), .Y(_7522_) );
AOI21X1 AOI21X1_1282 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_228_), .B(_7301__bF_buf3), .C(_7522_), .Y(_7523_) );
NOR2X1 NOR2X1_1290 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_229_), .B(_7315__bF_buf2), .Y(_7524_) );
INVX1 INVX1_546 ( .gnd(gnd), .vdd(vdd), .A(_7524_), .Y(_7525_) );
NAND2X1 NAND2X1_976 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_229_), .B(_7315__bF_buf1), .Y(_7526_) );
NAND2X1 NAND2X1_977 ( .gnd(gnd), .vdd(vdd), .A(_7526_), .B(_7525_), .Y(_7527_) );
XNOR2X1 XNOR2X1_306 ( .gnd(gnd), .vdd(vdd), .A(_7523_), .B(_7527_), .Y(_7528_) );
AOI21X1 AOI21X1_1283 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe64_bF_buf1), .B(_7528_), .C(micro_hash_ucr_2_pipe66_bF_buf1), .Y(_7529_) );
AOI21X1 AOI21X1_1284 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_236_), .B(_7301__bF_buf2), .C(_7284_), .Y(_7530_) );
NOR2X1 NOR2X1_1291 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_237_), .B(_7315__bF_buf0), .Y(_7531_) );
INVX1 INVX1_547 ( .gnd(gnd), .vdd(vdd), .A(_7531_), .Y(_7532_) );
NAND2X1 NAND2X1_978 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_237_), .B(_7315__bF_buf5), .Y(_7533_) );
NAND2X1 NAND2X1_979 ( .gnd(gnd), .vdd(vdd), .A(_7533_), .B(_7532_), .Y(_7534_) );
AND2X2 AND2X2_489 ( .gnd(gnd), .vdd(vdd), .A(_7530_), .B(_7534_), .Y(_7535_) );
OAI21X1 OAI21X1_2088 ( .gnd(gnd), .vdd(vdd), .A(_7530_), .B(_7534_), .C(micro_hash_ucr_2_pipe66_bF_buf0), .Y(_7536_) );
OAI21X1 OAI21X1_2089 ( .gnd(gnd), .vdd(vdd), .A(_7535_), .B(_7536_), .C(_5075__bF_buf4), .Y(_7537_) );
AOI21X1 AOI21X1_1285 ( .gnd(gnd), .vdd(vdd), .A(_7529_), .B(_7521_), .C(_7537_), .Y(_7538_) );
AOI21X1 AOI21X1_1286 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_244_), .B(_7301__bF_buf1), .C(_7292_), .Y(_7539_) );
INVX1 INVX1_548 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_245_), .Y(_7540_) );
OAI21X1 OAI21X1_2090 ( .gnd(gnd), .vdd(vdd), .A(_7311__bF_buf1), .B(_7312_), .C(_7540_), .Y(_7541_) );
INVX1 INVX1_549 ( .gnd(gnd), .vdd(vdd), .A(_7541_), .Y(_7542_) );
NOR2X1 NOR2X1_1292 ( .gnd(gnd), .vdd(vdd), .A(_7540_), .B(_7316__bF_buf0), .Y(_7543_) );
NOR2X1 NOR2X1_1293 ( .gnd(gnd), .vdd(vdd), .A(_7542_), .B(_7543_), .Y(_7544_) );
AND2X2 AND2X2_490 ( .gnd(gnd), .vdd(vdd), .A(_7539_), .B(_7544_), .Y(_7545_) );
OAI21X1 OAI21X1_2091 ( .gnd(gnd), .vdd(vdd), .A(_7539_), .B(_7544_), .C(micro_hash_ucr_2_pipe68), .Y(_7546_) );
OAI21X1 OAI21X1_2092 ( .gnd(gnd), .vdd(vdd), .A(_7545_), .B(_7546_), .C(_6146_), .Y(_7547_) );
NAND2X1 NAND2X1_980 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_252_), .B(_7301__bF_buf0), .Y(_7548_) );
OAI21X1 OAI21X1_2093 ( .gnd(gnd), .vdd(vdd), .A(_7297_), .B(_7296_), .C(_7548_), .Y(_7549_) );
INVX1 INVX1_550 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_253_), .Y(_7550_) );
OAI21X1 OAI21X1_2094 ( .gnd(gnd), .vdd(vdd), .A(_7311__bF_buf0), .B(_7312_), .C(_7550_), .Y(_7551_) );
NOR2X1 NOR2X1_1294 ( .gnd(gnd), .vdd(vdd), .A(_7550_), .B(_7316__bF_buf3), .Y(_7552_) );
INVX1 INVX1_551 ( .gnd(gnd), .vdd(vdd), .A(_7552_), .Y(_7553_) );
NAND2X1 NAND2X1_981 ( .gnd(gnd), .vdd(vdd), .A(_7551_), .B(_7553_), .Y(_7554_) );
XOR2X1 XOR2X1_131 ( .gnd(gnd), .vdd(vdd), .A(_7554_), .B(_7549_), .Y(_7555_) );
OAI22X1 OAI22X1_101 ( .gnd(gnd), .vdd(vdd), .A(_7300_), .B(_7555_), .C(_7538_), .D(_7547_), .Y(_4493__5_) );
OAI21X1 OAI21X1_2095 ( .gnd(gnd), .vdd(vdd), .A(_6030_), .B(_7305_), .C(_7310_), .Y(_7556_) );
XOR2X1 XOR2X1_132 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_k_6_), .B(micro_hash_ucr_2_x_6_), .Y(_7557_) );
NOR2X1 NOR2X1_1295 ( .gnd(gnd), .vdd(vdd), .A(_7557_), .B(_7556_), .Y(_7558_) );
OAI21X1 OAI21X1_2096 ( .gnd(gnd), .vdd(vdd), .A(_7311__bF_buf3), .B(_7307_), .C(_7557_), .Y(_7559_) );
INVX2 INVX2_246 ( .gnd(gnd), .vdd(vdd), .A(_7559_), .Y(_7560_) );
NOR2X1 NOR2X1_1296 ( .gnd(gnd), .vdd(vdd), .A(_7558_), .B(_7560_), .Y(_7561_) );
INVX8 INVX8_193 ( .gnd(gnd), .vdd(vdd), .A(_7561__bF_buf4), .Y(_7562_) );
NOR2X1 NOR2X1_1297 ( .gnd(gnd), .vdd(vdd), .A(_4806_), .B(_7562__bF_buf4), .Y(_7563_) );
INVX1 INVX1_552 ( .gnd(gnd), .vdd(vdd), .A(_7563_), .Y(_7564_) );
OAI21X1 OAI21X1_2097 ( .gnd(gnd), .vdd(vdd), .A(_7560_), .B(_7558_), .C(_4806_), .Y(_7565_) );
NAND2X1 NAND2X1_982 ( .gnd(gnd), .vdd(vdd), .A(_7565_), .B(_7564_), .Y(_7566_) );
INVX1 INVX1_553 ( .gnd(gnd), .vdd(vdd), .A(_7489_), .Y(_7567_) );
OAI21X1 OAI21X1_2098 ( .gnd(gnd), .vdd(vdd), .A(_7487_), .B(_7488_), .C(_7567_), .Y(_7568_) );
XOR2X1 XOR2X1_133 ( .gnd(gnd), .vdd(vdd), .A(_7566_), .B(_7568_), .Y(_7569_) );
XOR2X1 XOR2X1_134 ( .gnd(gnd), .vdd(vdd), .A(_7561__bF_buf3), .B(micro_hash_ucr_2_Wx_14_), .Y(_7570_) );
OAI21X1 OAI21X1_2099 ( .gnd(gnd), .vdd(vdd), .A(_7335_), .B(_7336_), .C(_7338_), .Y(_7571_) );
XNOR2X1 XNOR2X1_307 ( .gnd(gnd), .vdd(vdd), .A(_7571_), .B(_7570_), .Y(_7572_) );
XNOR2X1 XNOR2X1_308 ( .gnd(gnd), .vdd(vdd), .A(_7561__bF_buf2), .B(micro_hash_ucr_2_Wx_6_), .Y(_7573_) );
INVX1 INVX1_554 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_5_), .Y(_7574_) );
OAI21X1 OAI21X1_2100 ( .gnd(gnd), .vdd(vdd), .A(_7574_), .B(_7316__bF_buf2), .C(_7326_), .Y(_7575_) );
OAI21X1 OAI21X1_2101 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_5_), .B(_7315__bF_buf4), .C(_7575_), .Y(_7576_) );
OAI21X1 OAI21X1_2102 ( .gnd(gnd), .vdd(vdd), .A(_7576_), .B(_7573_), .C(micro_hash_ucr_2_pipe8), .Y(_7577_) );
AOI21X1 AOI21X1_1287 ( .gnd(gnd), .vdd(vdd), .A(_7573_), .B(_7576_), .C(_7577_), .Y(_7578_) );
NAND2X1 NAND2X1_983 ( .gnd(gnd), .vdd(vdd), .A(H_2_22_), .B(micro_hash_ucr_2_pipe6), .Y(_7579_) );
OAI21X1 OAI21X1_2103 ( .gnd(gnd), .vdd(vdd), .A(_8681_), .B(micro_hash_ucr_2_pipe6), .C(_7579_), .Y(_7580_) );
AOI21X1 AOI21X1_1288 ( .gnd(gnd), .vdd(vdd), .A(_5135_), .B(_7580_), .C(_7578_), .Y(_7581_) );
MUX2X1 MUX2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_7581_), .B(_7572_), .S(_5133_), .Y(_7582_) );
INVX1 INVX1_555 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_22_), .Y(_7583_) );
NOR2X1 NOR2X1_1298 ( .gnd(gnd), .vdd(vdd), .A(_7583_), .B(_7562__bF_buf3), .Y(_7584_) );
NOR2X1 NOR2X1_1299 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_22_), .B(_7561__bF_buf1), .Y(_7585_) );
NOR2X1 NOR2X1_1300 ( .gnd(gnd), .vdd(vdd), .A(_7585_), .B(_7584_), .Y(_7586_) );
INVX1 INVX1_556 ( .gnd(gnd), .vdd(vdd), .A(_7342_), .Y(_7587_) );
OAI21X1 OAI21X1_2104 ( .gnd(gnd), .vdd(vdd), .A(_7587_), .B(_7343_), .C(_7345_), .Y(_7588_) );
XOR2X1 XOR2X1_135 ( .gnd(gnd), .vdd(vdd), .A(_7588_), .B(_7586_), .Y(_7589_) );
MUX2X1 MUX2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_7582_), .B(_7589_), .S(_5128_), .Y(_7590_) );
INVX2 INVX2_247 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_30_), .Y(_7591_) );
XNOR2X1 XNOR2X1_309 ( .gnd(gnd), .vdd(vdd), .A(_7561__bF_buf0), .B(_7591_), .Y(_7592_) );
OAI21X1 OAI21X1_2105 ( .gnd(gnd), .vdd(vdd), .A(_7351_), .B(_7352_), .C(_7354_), .Y(_7593_) );
XNOR2X1 XNOR2X1_310 ( .gnd(gnd), .vdd(vdd), .A(_7592_), .B(_7593_), .Y(_7594_) );
MUX2X1 MUX2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_7590_), .B(_7594_), .S(_5129_), .Y(_7595_) );
NAND2X1 NAND2X1_984 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_38_), .B(_7561__bF_buf4), .Y(_7596_) );
INVX1 INVX1_557 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_38_), .Y(_7597_) );
OAI21X1 OAI21X1_2106 ( .gnd(gnd), .vdd(vdd), .A(_7560_), .B(_7558_), .C(_7597_), .Y(_7598_) );
AND2X2 AND2X2_491 ( .gnd(gnd), .vdd(vdd), .A(_7596_), .B(_7598_), .Y(_7599_) );
AOI21X1 AOI21X1_1289 ( .gnd(gnd), .vdd(vdd), .A(_7362_), .B(_7360_), .C(_7363_), .Y(_7600_) );
XNOR2X1 XNOR2X1_311 ( .gnd(gnd), .vdd(vdd), .A(_7600_), .B(_7599_), .Y(_7601_) );
MUX2X1 MUX2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_7595_), .B(_7601_), .S(_5127__bF_buf3), .Y(_7602_) );
INVX2 INVX2_248 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_46_), .Y(_7603_) );
XNOR2X1 XNOR2X1_312 ( .gnd(gnd), .vdd(vdd), .A(_7561__bF_buf3), .B(_7603_), .Y(_7604_) );
OAI21X1 OAI21X1_2107 ( .gnd(gnd), .vdd(vdd), .A(_7369_), .B(_7370_), .C(_7372_), .Y(_7605_) );
OR2X2 OR2X2_56 ( .gnd(gnd), .vdd(vdd), .A(_7605_), .B(_7604_), .Y(_7606_) );
NAND2X1 NAND2X1_985 ( .gnd(gnd), .vdd(vdd), .A(_7604_), .B(_7605_), .Y(_7607_) );
NAND3X1 NAND3X1_320 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe18_bF_buf0), .B(_7607_), .C(_7606_), .Y(_7608_) );
OAI21X1 OAI21X1_2108 ( .gnd(gnd), .vdd(vdd), .A(_7602_), .B(micro_hash_ucr_2_pipe18_bF_buf4), .C(_7608_), .Y(_7609_) );
INVX2 INVX2_249 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_54_), .Y(_7610_) );
XNOR2X1 XNOR2X1_313 ( .gnd(gnd), .vdd(vdd), .A(_7561__bF_buf2), .B(_7610_), .Y(_7611_) );
OAI21X1 OAI21X1_2109 ( .gnd(gnd), .vdd(vdd), .A(_7378_), .B(_7379_), .C(_7381_), .Y(_7612_) );
OAI21X1 OAI21X1_2110 ( .gnd(gnd), .vdd(vdd), .A(_7612_), .B(_7611_), .C(micro_hash_ucr_2_pipe20_bF_buf2), .Y(_7613_) );
AOI21X1 AOI21X1_1290 ( .gnd(gnd), .vdd(vdd), .A(_7611_), .B(_7612_), .C(_7613_), .Y(_7614_) );
AOI21X1 AOI21X1_1291 ( .gnd(gnd), .vdd(vdd), .A(_5123__bF_buf1), .B(_7609_), .C(_7614_), .Y(_7615_) );
NAND2X1 NAND2X1_986 ( .gnd(gnd), .vdd(vdd), .A(_5121__bF_buf1), .B(_7615_), .Y(_7616_) );
XNOR2X1 XNOR2X1_314 ( .gnd(gnd), .vdd(vdd), .A(_7561__bF_buf1), .B(_5022_), .Y(_7617_) );
OAI21X1 OAI21X1_2111 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_61_), .B(_7315__bF_buf3), .C(_7385_), .Y(_7618_) );
OAI21X1 OAI21X1_2112 ( .gnd(gnd), .vdd(vdd), .A(_5019_), .B(_7316__bF_buf1), .C(_7618_), .Y(_7619_) );
XOR2X1 XOR2X1_136 ( .gnd(gnd), .vdd(vdd), .A(_7619_), .B(_7617_), .Y(_7620_) );
OAI21X1 OAI21X1_2113 ( .gnd(gnd), .vdd(vdd), .A(_5121__bF_buf0), .B(_7620_), .C(_7616_), .Y(_7621_) );
XNOR2X1 XNOR2X1_315 ( .gnd(gnd), .vdd(vdd), .A(_7561__bF_buf0), .B(_4887_), .Y(_7622_) );
INVX1 INVX1_558 ( .gnd(gnd), .vdd(vdd), .A(_7622_), .Y(_7623_) );
AOI21X1 AOI21X1_1292 ( .gnd(gnd), .vdd(vdd), .A(_7393_), .B(_7392_), .C(_7394_), .Y(_7624_) );
OR2X2 OR2X2_57 ( .gnd(gnd), .vdd(vdd), .A(_7623_), .B(_7624_), .Y(_7625_) );
NAND2X1 NAND2X1_987 ( .gnd(gnd), .vdd(vdd), .A(_7624_), .B(_7623_), .Y(_7626_) );
NAND3X1 NAND3X1_321 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe24_bF_buf1), .B(_7626_), .C(_7625_), .Y(_7627_) );
OAI21X1 OAI21X1_2114 ( .gnd(gnd), .vdd(vdd), .A(_7621_), .B(micro_hash_ucr_2_pipe24_bF_buf0), .C(_7627_), .Y(_7628_) );
XNOR2X1 XNOR2X1_316 ( .gnd(gnd), .vdd(vdd), .A(_7561__bF_buf4), .B(_5044_), .Y(_7629_) );
INVX1 INVX1_559 ( .gnd(gnd), .vdd(vdd), .A(_7401_), .Y(_7630_) );
OAI21X1 OAI21X1_2115 ( .gnd(gnd), .vdd(vdd), .A(_7400_), .B(_7630_), .C(_7402_), .Y(_7631_) );
NOR2X1 NOR2X1_1301 ( .gnd(gnd), .vdd(vdd), .A(_7629_), .B(_7631_), .Y(_7632_) );
NAND2X1 NAND2X1_988 ( .gnd(gnd), .vdd(vdd), .A(_7629_), .B(_7631_), .Y(_7633_) );
NAND2X1 NAND2X1_989 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe26_bF_buf1), .B(_7633_), .Y(_7634_) );
OAI21X1 OAI21X1_2116 ( .gnd(gnd), .vdd(vdd), .A(_7634_), .B(_7632_), .C(_5115__bF_buf4), .Y(_7635_) );
AOI21X1 AOI21X1_1293 ( .gnd(gnd), .vdd(vdd), .A(_5117__bF_buf3), .B(_7628_), .C(_7635_), .Y(_7636_) );
XNOR2X1 XNOR2X1_317 ( .gnd(gnd), .vdd(vdd), .A(_7561__bF_buf3), .B(_4953_), .Y(_7637_) );
OAI21X1 OAI21X1_2117 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_85_), .B(_7315__bF_buf2), .C(_7408_), .Y(_7638_) );
OAI21X1 OAI21X1_2118 ( .gnd(gnd), .vdd(vdd), .A(_4950_), .B(_7316__bF_buf0), .C(_7638_), .Y(_7639_) );
XOR2X1 XOR2X1_137 ( .gnd(gnd), .vdd(vdd), .A(_7639_), .B(_7637_), .Y(_7640_) );
OAI21X1 OAI21X1_2119 ( .gnd(gnd), .vdd(vdd), .A(_7640_), .B(_5115__bF_buf3), .C(_5110__bF_buf2), .Y(_7641_) );
XNOR2X1 XNOR2X1_318 ( .gnd(gnd), .vdd(vdd), .A(_7561__bF_buf2), .B(_4998_), .Y(_7642_) );
INVX1 INVX1_560 ( .gnd(gnd), .vdd(vdd), .A(_7642_), .Y(_7643_) );
AOI21X1 AOI21X1_1294 ( .gnd(gnd), .vdd(vdd), .A(_7413_), .B(_7412_), .C(_7415_), .Y(_7644_) );
OR2X2 OR2X2_58 ( .gnd(gnd), .vdd(vdd), .A(_7644_), .B(_7643_), .Y(_7645_) );
NAND2X1 NAND2X1_990 ( .gnd(gnd), .vdd(vdd), .A(_7643_), .B(_7644_), .Y(_7646_) );
NAND2X1 NAND2X1_991 ( .gnd(gnd), .vdd(vdd), .A(_7646_), .B(_7645_), .Y(_7647_) );
OAI22X1 OAI22X1_102 ( .gnd(gnd), .vdd(vdd), .A(_5110__bF_buf1), .B(_7647_), .C(_7636_), .D(_7641_), .Y(_7648_) );
XNOR2X1 XNOR2X1_319 ( .gnd(gnd), .vdd(vdd), .A(_7561__bF_buf1), .B(micro_hash_ucr_2_Wx_102_), .Y(_7649_) );
OAI21X1 OAI21X1_2120 ( .gnd(gnd), .vdd(vdd), .A(_4858_), .B(_7316__bF_buf3), .C(_7420_), .Y(_7650_) );
OAI21X1 OAI21X1_2121 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_101_), .B(_7315__bF_buf1), .C(_7650_), .Y(_7651_) );
NAND2X1 NAND2X1_992 ( .gnd(gnd), .vdd(vdd), .A(_7649_), .B(_7651_), .Y(_7652_) );
OR2X2 OR2X2_59 ( .gnd(gnd), .vdd(vdd), .A(_7651_), .B(_7649_), .Y(_7653_) );
NAND2X1 NAND2X1_993 ( .gnd(gnd), .vdd(vdd), .A(_7652_), .B(_7653_), .Y(_7654_) );
OAI21X1 OAI21X1_2122 ( .gnd(gnd), .vdd(vdd), .A(_7654_), .B(_5111__bF_buf4), .C(_5109__bF_buf0), .Y(_7655_) );
AOI21X1 AOI21X1_1295 ( .gnd(gnd), .vdd(vdd), .A(_5111__bF_buf3), .B(_7648_), .C(_7655_), .Y(_7656_) );
XNOR2X1 XNOR2X1_320 ( .gnd(gnd), .vdd(vdd), .A(_7561__bF_buf0), .B(micro_hash_ucr_2_Wx_110_), .Y(_7657_) );
AOI21X1 AOI21X1_1296 ( .gnd(gnd), .vdd(vdd), .A(_7425_), .B(_7424_), .C(_7426_), .Y(_7658_) );
XOR2X1 XOR2X1_138 ( .gnd(gnd), .vdd(vdd), .A(_7658_), .B(_7657_), .Y(_7659_) );
OAI21X1 OAI21X1_2123 ( .gnd(gnd), .vdd(vdd), .A(_7659_), .B(_5109__bF_buf4), .C(_5104__bF_buf4), .Y(_7660_) );
NOR2X1 NOR2X1_1302 ( .gnd(gnd), .vdd(vdd), .A(_7660_), .B(_7656_), .Y(_7661_) );
XNOR2X1 XNOR2X1_321 ( .gnd(gnd), .vdd(vdd), .A(_7561__bF_buf4), .B(micro_hash_ucr_2_Wx_118_), .Y(_7662_) );
AOI21X1 AOI21X1_1297 ( .gnd(gnd), .vdd(vdd), .A(_7433_), .B(_7432_), .C(_7434_), .Y(_7663_) );
OR2X2 OR2X2_60 ( .gnd(gnd), .vdd(vdd), .A(_7663_), .B(_7662_), .Y(_7664_) );
AOI21X1 AOI21X1_1298 ( .gnd(gnd), .vdd(vdd), .A(_7662_), .B(_7663_), .C(_5104__bF_buf3), .Y(_7665_) );
AND2X2 AND2X2_492 ( .gnd(gnd), .vdd(vdd), .A(_7664_), .B(_7665_), .Y(_7666_) );
OAI21X1 OAI21X1_2124 ( .gnd(gnd), .vdd(vdd), .A(_7661_), .B(_7666_), .C(_5105__bF_buf3), .Y(_7667_) );
XNOR2X1 XNOR2X1_322 ( .gnd(gnd), .vdd(vdd), .A(_7561__bF_buf3), .B(_4909_), .Y(_7668_) );
OAI21X1 OAI21X1_2125 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_125_), .B(_7315__bF_buf0), .C(_7439_), .Y(_7669_) );
OAI21X1 OAI21X1_2126 ( .gnd(gnd), .vdd(vdd), .A(_4906_), .B(_7316__bF_buf2), .C(_7669_), .Y(_7670_) );
OR2X2 OR2X2_61 ( .gnd(gnd), .vdd(vdd), .A(_7670_), .B(_7668_), .Y(_7671_) );
NAND2X1 NAND2X1_994 ( .gnd(gnd), .vdd(vdd), .A(_7668_), .B(_7670_), .Y(_7672_) );
NAND3X1 NAND3X1_322 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe38_bF_buf1), .B(_7672_), .C(_7671_), .Y(_7673_) );
AOI21X1 AOI21X1_1299 ( .gnd(gnd), .vdd(vdd), .A(_7673_), .B(_7667_), .C(micro_hash_ucr_2_pipe40_bF_buf0), .Y(_7674_) );
XNOR2X1 XNOR2X1_323 ( .gnd(gnd), .vdd(vdd), .A(_7561__bF_buf2), .B(_4805_), .Y(_7675_) );
AOI21X1 AOI21X1_1300 ( .gnd(gnd), .vdd(vdd), .A(_7445_), .B(_7444_), .C(_7446_), .Y(_7676_) );
INVX1 INVX1_561 ( .gnd(gnd), .vdd(vdd), .A(_7676_), .Y(_7677_) );
NOR2X1 NOR2X1_1303 ( .gnd(gnd), .vdd(vdd), .A(_7675_), .B(_7677_), .Y(_7678_) );
NAND2X1 NAND2X1_995 ( .gnd(gnd), .vdd(vdd), .A(_7675_), .B(_7677_), .Y(_7679_) );
NAND2X1 NAND2X1_996 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe40_bF_buf4), .B(_7679_), .Y(_7680_) );
OAI21X1 OAI21X1_2127 ( .gnd(gnd), .vdd(vdd), .A(_7680_), .B(_7678_), .C(_5098__bF_buf0), .Y(_7681_) );
XNOR2X1 XNOR2X1_324 ( .gnd(gnd), .vdd(vdd), .A(_7561__bF_buf1), .B(_4999_), .Y(_7682_) );
INVX1 INVX1_562 ( .gnd(gnd), .vdd(vdd), .A(_7453_), .Y(_7683_) );
OAI21X1 OAI21X1_2128 ( .gnd(gnd), .vdd(vdd), .A(_7452_), .B(_7683_), .C(_7454_), .Y(_7684_) );
XOR2X1 XOR2X1_139 ( .gnd(gnd), .vdd(vdd), .A(_7684_), .B(_7682_), .Y(_7685_) );
OAI22X1 OAI22X1_103 ( .gnd(gnd), .vdd(vdd), .A(_5098__bF_buf4), .B(_7685_), .C(_7674_), .D(_7681_), .Y(_7686_) );
XNOR2X1 XNOR2X1_325 ( .gnd(gnd), .vdd(vdd), .A(_7561__bF_buf0), .B(_4833_), .Y(_7687_) );
INVX1 INVX1_563 ( .gnd(gnd), .vdd(vdd), .A(_7687_), .Y(_7688_) );
AOI21X1 AOI21X1_1301 ( .gnd(gnd), .vdd(vdd), .A(_7461_), .B(_7460_), .C(_7462_), .Y(_7689_) );
OR2X2 OR2X2_62 ( .gnd(gnd), .vdd(vdd), .A(_7689_), .B(_7688_), .Y(_7690_) );
NAND2X1 NAND2X1_997 ( .gnd(gnd), .vdd(vdd), .A(_7688_), .B(_7689_), .Y(_7691_) );
AOI21X1 AOI21X1_1302 ( .gnd(gnd), .vdd(vdd), .A(_7691_), .B(_7690_), .C(_5099__bF_buf0), .Y(_7692_) );
AOI21X1 AOI21X1_1303 ( .gnd(gnd), .vdd(vdd), .A(_5099__bF_buf4), .B(_7686_), .C(_7692_), .Y(_7693_) );
XNOR2X1 XNOR2X1_326 ( .gnd(gnd), .vdd(vdd), .A(_7561__bF_buf4), .B(_4719_), .Y(_7694_) );
OAI21X1 OAI21X1_2129 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_157_), .B(_7315__bF_buf5), .C(_7468_), .Y(_7695_) );
OAI21X1 OAI21X1_2130 ( .gnd(gnd), .vdd(vdd), .A(_4716_), .B(_7316__bF_buf1), .C(_7695_), .Y(_7696_) );
NOR2X1 NOR2X1_1304 ( .gnd(gnd), .vdd(vdd), .A(_7694_), .B(_7696_), .Y(_7697_) );
NAND2X1 NAND2X1_998 ( .gnd(gnd), .vdd(vdd), .A(_7694_), .B(_7696_), .Y(_7698_) );
NAND2X1 NAND2X1_999 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe46_bF_buf1), .B(_7698_), .Y(_7699_) );
OAI21X1 OAI21X1_2131 ( .gnd(gnd), .vdd(vdd), .A(_7699_), .B(_7697_), .C(_5092__bF_buf1), .Y(_7700_) );
AOI21X1 AOI21X1_1304 ( .gnd(gnd), .vdd(vdd), .A(_5097__bF_buf3), .B(_7693_), .C(_7700_), .Y(_7701_) );
XNOR2X1 XNOR2X1_327 ( .gnd(gnd), .vdd(vdd), .A(_7561__bF_buf3), .B(_4774_), .Y(_7702_) );
INVX1 INVX1_564 ( .gnd(gnd), .vdd(vdd), .A(_7474_), .Y(_7703_) );
OAI21X1 OAI21X1_2132 ( .gnd(gnd), .vdd(vdd), .A(_7473_), .B(_7703_), .C(_7475_), .Y(_7704_) );
XOR2X1 XOR2X1_140 ( .gnd(gnd), .vdd(vdd), .A(_7704_), .B(_7702_), .Y(_7705_) );
OAI21X1 OAI21X1_2133 ( .gnd(gnd), .vdd(vdd), .A(_7705_), .B(_5092__bF_buf0), .C(_5093__bF_buf3), .Y(_7706_) );
NOR2X1 NOR2X1_1305 ( .gnd(gnd), .vdd(vdd), .A(_7706_), .B(_7701_), .Y(_7707_) );
XNOR2X1 XNOR2X1_328 ( .gnd(gnd), .vdd(vdd), .A(_7561__bF_buf2), .B(micro_hash_ucr_2_Wx_174_), .Y(_7708_) );
AOI21X1 AOI21X1_1305 ( .gnd(gnd), .vdd(vdd), .A(_7480_), .B(_7479_), .C(_7481_), .Y(_7709_) );
OR2X2 OR2X2_63 ( .gnd(gnd), .vdd(vdd), .A(_7709_), .B(_7708_), .Y(_7710_) );
AOI21X1 AOI21X1_1306 ( .gnd(gnd), .vdd(vdd), .A(_7708_), .B(_7709_), .C(_5093__bF_buf2), .Y(_7711_) );
AND2X2 AND2X2_493 ( .gnd(gnd), .vdd(vdd), .A(_7710_), .B(_7711_), .Y(_7712_) );
OAI21X1 OAI21X1_2134 ( .gnd(gnd), .vdd(vdd), .A(_7707_), .B(_7712_), .C(_5091__bF_buf0), .Y(_7713_) );
OAI21X1 OAI21X1_2135 ( .gnd(gnd), .vdd(vdd), .A(_5091__bF_buf4), .B(_7569_), .C(_7713_), .Y(_7714_) );
XNOR2X1 XNOR2X1_329 ( .gnd(gnd), .vdd(vdd), .A(_7561__bF_buf1), .B(_4863_), .Y(_7715_) );
INVX1 INVX1_565 ( .gnd(gnd), .vdd(vdd), .A(_7323_), .Y(_7716_) );
OAI21X1 OAI21X1_2136 ( .gnd(gnd), .vdd(vdd), .A(_7320_), .B(_7322_), .C(_7716_), .Y(_7717_) );
NAND2X1 NAND2X1_1000 ( .gnd(gnd), .vdd(vdd), .A(_7715_), .B(_7717_), .Y(_7718_) );
INVX1 INVX1_566 ( .gnd(gnd), .vdd(vdd), .A(_7718_), .Y(_7719_) );
OAI21X1 OAI21X1_2137 ( .gnd(gnd), .vdd(vdd), .A(_7717_), .B(_7715_), .C(micro_hash_ucr_2_pipe54_bF_buf1), .Y(_7720_) );
OAI21X1 OAI21X1_2138 ( .gnd(gnd), .vdd(vdd), .A(_7719_), .B(_7720_), .C(_5087__bF_buf4), .Y(_7721_) );
AOI21X1 AOI21X1_1307 ( .gnd(gnd), .vdd(vdd), .A(_5086__bF_buf3), .B(_7714_), .C(_7721_), .Y(_7722_) );
NOR2X1 NOR2X1_1306 ( .gnd(gnd), .vdd(vdd), .A(_4834_), .B(_7562__bF_buf2), .Y(_7723_) );
INVX1 INVX1_567 ( .gnd(gnd), .vdd(vdd), .A(_7723_), .Y(_7724_) );
OAI21X1 OAI21X1_2139 ( .gnd(gnd), .vdd(vdd), .A(_7560_), .B(_7558_), .C(_4834_), .Y(_7725_) );
NAND2X1 NAND2X1_1001 ( .gnd(gnd), .vdd(vdd), .A(_7725_), .B(_7724_), .Y(_7726_) );
OAI21X1 OAI21X1_2140 ( .gnd(gnd), .vdd(vdd), .A(_7496_), .B(_7497_), .C(_7499_), .Y(_7727_) );
XNOR2X1 XNOR2X1_330 ( .gnd(gnd), .vdd(vdd), .A(_7726_), .B(_7727_), .Y(_7728_) );
OAI21X1 OAI21X1_2141 ( .gnd(gnd), .vdd(vdd), .A(_7728_), .B(_5087__bF_buf3), .C(_5085__bF_buf3), .Y(_7729_) );
XNOR2X1 XNOR2X1_331 ( .gnd(gnd), .vdd(vdd), .A(_7561__bF_buf0), .B(_4720_), .Y(_7730_) );
OAI21X1 OAI21X1_2142 ( .gnd(gnd), .vdd(vdd), .A(_7503_), .B(_7504_), .C(_7506_), .Y(_7731_) );
XOR2X1 XOR2X1_141 ( .gnd(gnd), .vdd(vdd), .A(_7731_), .B(_7730_), .Y(_7732_) );
AOI21X1 AOI21X1_1308 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe58_bF_buf1), .B(_7732_), .C(micro_hash_ucr_2_pipe60_bF_buf3), .Y(_7733_) );
OAI21X1 OAI21X1_2143 ( .gnd(gnd), .vdd(vdd), .A(_7722_), .B(_7729_), .C(_7733_), .Y(_7734_) );
XNOR2X1 XNOR2X1_332 ( .gnd(gnd), .vdd(vdd), .A(_7561__bF_buf4), .B(_4775_), .Y(_7735_) );
OAI21X1 OAI21X1_2144 ( .gnd(gnd), .vdd(vdd), .A(_7512_), .B(_7513_), .C(_7514_), .Y(_7736_) );
XNOR2X1 XNOR2X1_333 ( .gnd(gnd), .vdd(vdd), .A(_7736_), .B(_7735_), .Y(_7737_) );
AOI21X1 AOI21X1_1309 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe60_bF_buf2), .B(_7737_), .C(micro_hash_ucr_2_pipe62_bF_buf3), .Y(_7738_) );
XNOR2X1 XNOR2X1_334 ( .gnd(gnd), .vdd(vdd), .A(_7561__bF_buf3), .B(_4748_), .Y(_7739_) );
INVX1 INVX1_568 ( .gnd(gnd), .vdd(vdd), .A(_7317_), .Y(_7740_) );
OAI21X1 OAI21X1_2145 ( .gnd(gnd), .vdd(vdd), .A(_7302_), .B(_7314_), .C(_7740_), .Y(_7741_) );
NAND2X1 NAND2X1_1002 ( .gnd(gnd), .vdd(vdd), .A(_7739_), .B(_7741_), .Y(_7742_) );
NOR2X1 NOR2X1_1307 ( .gnd(gnd), .vdd(vdd), .A(_7739_), .B(_7741_), .Y(_7743_) );
NOR2X1 NOR2X1_1308 ( .gnd(gnd), .vdd(vdd), .A(_5081__bF_buf1), .B(_7743_), .Y(_7744_) );
AOI22X1 AOI22X1_58 ( .gnd(gnd), .vdd(vdd), .A(_7742_), .B(_7744_), .C(_7734_), .D(_7738_), .Y(_7745_) );
INVX2 INVX2_250 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_230_), .Y(_7746_) );
XNOR2X1 XNOR2X1_335 ( .gnd(gnd), .vdd(vdd), .A(_7561__bF_buf2), .B(_7746_), .Y(_7747_) );
OAI21X1 OAI21X1_2146 ( .gnd(gnd), .vdd(vdd), .A(_7523_), .B(_7524_), .C(_7526_), .Y(_7748_) );
XOR2X1 XOR2X1_142 ( .gnd(gnd), .vdd(vdd), .A(_7748_), .B(_7747_), .Y(_7749_) );
AOI21X1 AOI21X1_1310 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe64_bF_buf0), .B(_7749_), .C(micro_hash_ucr_2_pipe66_bF_buf4), .Y(_7750_) );
OAI21X1 OAI21X1_2147 ( .gnd(gnd), .vdd(vdd), .A(_7745_), .B(micro_hash_ucr_2_pipe64_bF_buf4), .C(_7750_), .Y(_7751_) );
INVX2 INVX2_251 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_238_), .Y(_7752_) );
XNOR2X1 XNOR2X1_336 ( .gnd(gnd), .vdd(vdd), .A(_7561__bF_buf1), .B(_7752_), .Y(_7753_) );
OAI21X1 OAI21X1_2148 ( .gnd(gnd), .vdd(vdd), .A(_7530_), .B(_7531_), .C(_7533_), .Y(_7754_) );
NOR2X1 NOR2X1_1309 ( .gnd(gnd), .vdd(vdd), .A(_7753_), .B(_7754_), .Y(_7755_) );
NAND2X1 NAND2X1_1003 ( .gnd(gnd), .vdd(vdd), .A(_7753_), .B(_7754_), .Y(_7756_) );
INVX1 INVX1_569 ( .gnd(gnd), .vdd(vdd), .A(_7756_), .Y(_7757_) );
OAI21X1 OAI21X1_2149 ( .gnd(gnd), .vdd(vdd), .A(_7757_), .B(_7755_), .C(micro_hash_ucr_2_pipe66_bF_buf3), .Y(_7758_) );
NAND3X1 NAND3X1_323 ( .gnd(gnd), .vdd(vdd), .A(_5075__bF_buf3), .B(_7758_), .C(_7751_), .Y(_7759_) );
INVX2 INVX2_252 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_246_), .Y(_7760_) );
XNOR2X1 XNOR2X1_337 ( .gnd(gnd), .vdd(vdd), .A(_7561__bF_buf0), .B(_7760_), .Y(_7761_) );
INVX1 INVX1_570 ( .gnd(gnd), .vdd(vdd), .A(_7543_), .Y(_7762_) );
OAI21X1 OAI21X1_2150 ( .gnd(gnd), .vdd(vdd), .A(_7539_), .B(_7542_), .C(_7762_), .Y(_7763_) );
XOR2X1 XOR2X1_143 ( .gnd(gnd), .vdd(vdd), .A(_7763_), .B(_7761_), .Y(_7764_) );
AOI21X1 AOI21X1_1311 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe68), .B(_7764_), .C(micro_hash_ucr_2_pipe69), .Y(_7765_) );
XNOR2X1 XNOR2X1_338 ( .gnd(gnd), .vdd(vdd), .A(_7561__bF_buf4), .B(micro_hash_ucr_2_Wx_254_), .Y(_7766_) );
AOI21X1 AOI21X1_1312 ( .gnd(gnd), .vdd(vdd), .A(_7551_), .B(_7549_), .C(_7552_), .Y(_7767_) );
AND2X2 AND2X2_494 ( .gnd(gnd), .vdd(vdd), .A(_7767_), .B(_7766_), .Y(_7768_) );
NOR2X1 NOR2X1_1310 ( .gnd(gnd), .vdd(vdd), .A(_4594__bF_buf11), .B(_7768_), .Y(_7769_) );
OAI21X1 OAI21X1_2151 ( .gnd(gnd), .vdd(vdd), .A(_7766_), .B(_7767_), .C(_7769_), .Y(_7770_) );
AOI22X1 AOI22X1_59 ( .gnd(gnd), .vdd(vdd), .A(_6147_), .B(_7770_), .C(_7759_), .D(_7765_), .Y(_4493__6_) );
NAND2X1 NAND2X1_1004 ( .gnd(gnd), .vdd(vdd), .A(_7735_), .B(_7736_), .Y(_7771_) );
OAI21X1 OAI21X1_2152 ( .gnd(gnd), .vdd(vdd), .A(_4775_), .B(_7562__bF_buf1), .C(_7771_), .Y(_7772_) );
NAND2X1 NAND2X1_1005 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_k_6_), .B(micro_hash_ucr_2_x_6_), .Y(_7773_) );
NAND2X1 NAND2X1_1006 ( .gnd(gnd), .vdd(vdd), .A(_7773_), .B(_7559_), .Y(_7774_) );
XOR2X1 XOR2X1_144 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_k_7_), .B(micro_hash_ucr_2_x_7_), .Y(_7775_) );
XOR2X1 XOR2X1_145 ( .gnd(gnd), .vdd(vdd), .A(_7774_), .B(_7775_), .Y(_7776_) );
XNOR2X1 XNOR2X1_339 ( .gnd(gnd), .vdd(vdd), .A(_7776__bF_buf4), .B(micro_hash_ucr_2_Wx_215_), .Y(_7777_) );
XNOR2X1 XNOR2X1_340 ( .gnd(gnd), .vdd(vdd), .A(_7772_), .B(_7777_), .Y(_7778_) );
NAND2X1 NAND2X1_1007 ( .gnd(gnd), .vdd(vdd), .A(_7702_), .B(_7704_), .Y(_7779_) );
OAI21X1 OAI21X1_2153 ( .gnd(gnd), .vdd(vdd), .A(_4774_), .B(_7562__bF_buf0), .C(_7779_), .Y(_7780_) );
XNOR2X1 XNOR2X1_341 ( .gnd(gnd), .vdd(vdd), .A(_7776__bF_buf3), .B(micro_hash_ucr_2_Wx_167_), .Y(_7781_) );
XNOR2X1 XNOR2X1_342 ( .gnd(gnd), .vdd(vdd), .A(_7780_), .B(_7781_), .Y(_7782_) );
NAND2X1 NAND2X1_1008 ( .gnd(gnd), .vdd(vdd), .A(_7682_), .B(_7684_), .Y(_7783_) );
OAI21X1 OAI21X1_2154 ( .gnd(gnd), .vdd(vdd), .A(_4999_), .B(_7562__bF_buf4), .C(_7783_), .Y(_7784_) );
XNOR2X1 XNOR2X1_343 ( .gnd(gnd), .vdd(vdd), .A(_7776__bF_buf2), .B(micro_hash_ucr_2_Wx_143_), .Y(_7785_) );
XNOR2X1 XNOR2X1_344 ( .gnd(gnd), .vdd(vdd), .A(_7784_), .B(_7785_), .Y(_7786_) );
OAI21X1 OAI21X1_2155 ( .gnd(gnd), .vdd(vdd), .A(_4998_), .B(_7562__bF_buf3), .C(_7645_), .Y(_7787_) );
XNOR2X1 XNOR2X1_345 ( .gnd(gnd), .vdd(vdd), .A(_7776__bF_buf1), .B(micro_hash_ucr_2_Wx_95_), .Y(_7788_) );
XNOR2X1 XNOR2X1_346 ( .gnd(gnd), .vdd(vdd), .A(_7787_), .B(_7788_), .Y(_7789_) );
NAND2X1 NAND2X1_1009 ( .gnd(gnd), .vdd(vdd), .A(_7617_), .B(_7619_), .Y(_7790_) );
OAI21X1 OAI21X1_2156 ( .gnd(gnd), .vdd(vdd), .A(_5022_), .B(_7562__bF_buf2), .C(_7790_), .Y(_7791_) );
XNOR2X1 XNOR2X1_347 ( .gnd(gnd), .vdd(vdd), .A(_7776__bF_buf0), .B(micro_hash_ucr_2_Wx_63_), .Y(_7792_) );
XNOR2X1 XNOR2X1_348 ( .gnd(gnd), .vdd(vdd), .A(_7791_), .B(_7792_), .Y(_7793_) );
NAND2X1 NAND2X1_1010 ( .gnd(gnd), .vdd(vdd), .A(_7593_), .B(_7592_), .Y(_7794_) );
OAI21X1 OAI21X1_2157 ( .gnd(gnd), .vdd(vdd), .A(_7591_), .B(_7562__bF_buf1), .C(_7794_), .Y(_7795_) );
XOR2X1 XOR2X1_146 ( .gnd(gnd), .vdd(vdd), .A(_7776__bF_buf4), .B(micro_hash_ucr_2_Wx_31_), .Y(_7796_) );
XOR2X1 XOR2X1_147 ( .gnd(gnd), .vdd(vdd), .A(_7795_), .B(_7796_), .Y(_7797_) );
NAND2X1 NAND2X1_1011 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_6_), .B(_7561__bF_buf3), .Y(_7798_) );
OAI21X1 OAI21X1_2158 ( .gnd(gnd), .vdd(vdd), .A(_7576_), .B(_7573_), .C(_7798_), .Y(_7799_) );
XNOR2X1 XNOR2X1_349 ( .gnd(gnd), .vdd(vdd), .A(_7776__bF_buf3), .B(micro_hash_ucr_2_Wx_7_), .Y(_7800_) );
AND2X2 AND2X2_495 ( .gnd(gnd), .vdd(vdd), .A(_7799_), .B(_7800_), .Y(_7801_) );
OAI21X1 OAI21X1_2159 ( .gnd(gnd), .vdd(vdd), .A(_7799_), .B(_7800_), .C(micro_hash_ucr_2_pipe8), .Y(_7802_) );
INVX1 INVX1_571 ( .gnd(gnd), .vdd(vdd), .A(H_2_23_), .Y(_7803_) );
AOI21X1 AOI21X1_1313 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_7_), .B(_5134_), .C(micro_hash_ucr_2_pipe8), .Y(_7804_) );
OAI21X1 OAI21X1_2160 ( .gnd(gnd), .vdd(vdd), .A(_7803_), .B(_5134_), .C(_7804_), .Y(_7805_) );
OAI21X1 OAI21X1_2161 ( .gnd(gnd), .vdd(vdd), .A(_7801_), .B(_7802_), .C(_7805_), .Y(_7806_) );
AND2X2 AND2X2_496 ( .gnd(gnd), .vdd(vdd), .A(_7561__bF_buf2), .B(micro_hash_ucr_2_Wx_14_), .Y(_7807_) );
AOI21X1 AOI21X1_1314 ( .gnd(gnd), .vdd(vdd), .A(_7570_), .B(_7571_), .C(_7807_), .Y(_7808_) );
XNOR2X1 XNOR2X1_350 ( .gnd(gnd), .vdd(vdd), .A(_7776__bF_buf2), .B(micro_hash_ucr_2_Wx_15_), .Y(_7809_) );
AND2X2 AND2X2_497 ( .gnd(gnd), .vdd(vdd), .A(_7808_), .B(_7809_), .Y(_7810_) );
OAI21X1 OAI21X1_2162 ( .gnd(gnd), .vdd(vdd), .A(_7808_), .B(_7809_), .C(micro_hash_ucr_2_pipe10), .Y(_7811_) );
OAI22X1 OAI22X1_104 ( .gnd(gnd), .vdd(vdd), .A(_7810_), .B(_7811_), .C(_7806_), .D(micro_hash_ucr_2_pipe10), .Y(_7812_) );
AOI21X1 AOI21X1_1315 ( .gnd(gnd), .vdd(vdd), .A(_7586_), .B(_7588_), .C(_7584_), .Y(_7813_) );
XOR2X1 XOR2X1_148 ( .gnd(gnd), .vdd(vdd), .A(_7776__bF_buf1), .B(micro_hash_ucr_2_Wx_23_), .Y(_7814_) );
AOI21X1 AOI21X1_1316 ( .gnd(gnd), .vdd(vdd), .A(_7814_), .B(_7813_), .C(_5128_), .Y(_7815_) );
OAI21X1 OAI21X1_2163 ( .gnd(gnd), .vdd(vdd), .A(_7813_), .B(_7814_), .C(_7815_), .Y(_7816_) );
OAI21X1 OAI21X1_2164 ( .gnd(gnd), .vdd(vdd), .A(_7812_), .B(micro_hash_ucr_2_pipe12_bF_buf3), .C(_7816_), .Y(_7817_) );
NAND2X1 NAND2X1_1012 ( .gnd(gnd), .vdd(vdd), .A(_5129_), .B(_7817_), .Y(_7818_) );
OAI21X1 OAI21X1_2165 ( .gnd(gnd), .vdd(vdd), .A(_5129_), .B(_7797_), .C(_7818_), .Y(_7819_) );
INVX1 INVX1_572 ( .gnd(gnd), .vdd(vdd), .A(_7599_), .Y(_7820_) );
OAI21X1 OAI21X1_2166 ( .gnd(gnd), .vdd(vdd), .A(_7600_), .B(_7820_), .C(_7596_), .Y(_7821_) );
XOR2X1 XOR2X1_149 ( .gnd(gnd), .vdd(vdd), .A(_7776__bF_buf0), .B(micro_hash_ucr_2_Wx_39_), .Y(_7822_) );
AOI21X1 AOI21X1_1317 ( .gnd(gnd), .vdd(vdd), .A(_7822_), .B(_7821_), .C(_5127__bF_buf2), .Y(_7823_) );
OAI21X1 OAI21X1_2167 ( .gnd(gnd), .vdd(vdd), .A(_7821_), .B(_7822_), .C(_7823_), .Y(_7824_) );
OAI21X1 OAI21X1_2168 ( .gnd(gnd), .vdd(vdd), .A(_7819_), .B(micro_hash_ucr_2_pipe16_bF_buf4), .C(_7824_), .Y(_7825_) );
OAI21X1 OAI21X1_2169 ( .gnd(gnd), .vdd(vdd), .A(_7603_), .B(_7562__bF_buf0), .C(_7607_), .Y(_7826_) );
XOR2X1 XOR2X1_150 ( .gnd(gnd), .vdd(vdd), .A(_7776__bF_buf4), .B(micro_hash_ucr_2_Wx_47_), .Y(_7827_) );
XNOR2X1 XNOR2X1_351 ( .gnd(gnd), .vdd(vdd), .A(_7826_), .B(_7827_), .Y(_7828_) );
OAI21X1 OAI21X1_2170 ( .gnd(gnd), .vdd(vdd), .A(_7828_), .B(_5122__bF_buf2), .C(_5123__bF_buf0), .Y(_7829_) );
AOI21X1 AOI21X1_1318 ( .gnd(gnd), .vdd(vdd), .A(_5122__bF_buf1), .B(_7825_), .C(_7829_), .Y(_7830_) );
NAND2X1 NAND2X1_1013 ( .gnd(gnd), .vdd(vdd), .A(_7611_), .B(_7612_), .Y(_7831_) );
OAI21X1 OAI21X1_2171 ( .gnd(gnd), .vdd(vdd), .A(_7610_), .B(_7562__bF_buf4), .C(_7831_), .Y(_7832_) );
XNOR2X1 XNOR2X1_352 ( .gnd(gnd), .vdd(vdd), .A(_7776__bF_buf3), .B(micro_hash_ucr_2_Wx_55_), .Y(_7833_) );
OAI21X1 OAI21X1_2172 ( .gnd(gnd), .vdd(vdd), .A(_7832_), .B(_7833_), .C(micro_hash_ucr_2_pipe20_bF_buf1), .Y(_7834_) );
AOI21X1 AOI21X1_1319 ( .gnd(gnd), .vdd(vdd), .A(_7832_), .B(_7833_), .C(_7834_), .Y(_7835_) );
OAI21X1 OAI21X1_2173 ( .gnd(gnd), .vdd(vdd), .A(_7830_), .B(_7835_), .C(_5121__bF_buf4), .Y(_7836_) );
OAI21X1 OAI21X1_2174 ( .gnd(gnd), .vdd(vdd), .A(_5121__bF_buf3), .B(_7793_), .C(_7836_), .Y(_7837_) );
OAI21X1 OAI21X1_2175 ( .gnd(gnd), .vdd(vdd), .A(_4887_), .B(_7562__bF_buf3), .C(_7625_), .Y(_7838_) );
XNOR2X1 XNOR2X1_353 ( .gnd(gnd), .vdd(vdd), .A(_7776__bF_buf2), .B(micro_hash_ucr_2_Wx_71_), .Y(_7839_) );
OAI21X1 OAI21X1_2176 ( .gnd(gnd), .vdd(vdd), .A(_7838_), .B(_7839_), .C(micro_hash_ucr_2_pipe24_bF_buf3), .Y(_7840_) );
AOI21X1 AOI21X1_1320 ( .gnd(gnd), .vdd(vdd), .A(_7838_), .B(_7839_), .C(_7840_), .Y(_7841_) );
AOI21X1 AOI21X1_1321 ( .gnd(gnd), .vdd(vdd), .A(_5116__bF_buf2), .B(_7837_), .C(_7841_), .Y(_7842_) );
OAI21X1 OAI21X1_2177 ( .gnd(gnd), .vdd(vdd), .A(_5044_), .B(_7562__bF_buf2), .C(_7633_), .Y(_7843_) );
XNOR2X1 XNOR2X1_354 ( .gnd(gnd), .vdd(vdd), .A(_7776__bF_buf1), .B(_5047_), .Y(_7844_) );
NOR2X1 NOR2X1_1311 ( .gnd(gnd), .vdd(vdd), .A(_7844_), .B(_7843_), .Y(_7845_) );
AND2X2 AND2X2_498 ( .gnd(gnd), .vdd(vdd), .A(_7843_), .B(_7844_), .Y(_7846_) );
OAI21X1 OAI21X1_2178 ( .gnd(gnd), .vdd(vdd), .A(_7846_), .B(_7845_), .C(micro_hash_ucr_2_pipe26_bF_buf0), .Y(_7847_) );
OAI21X1 OAI21X1_2179 ( .gnd(gnd), .vdd(vdd), .A(_7842_), .B(micro_hash_ucr_2_pipe26_bF_buf3), .C(_7847_), .Y(_7848_) );
AND2X2 AND2X2_499 ( .gnd(gnd), .vdd(vdd), .A(_7848_), .B(_5115__bF_buf2), .Y(_7849_) );
NAND2X1 NAND2X1_1014 ( .gnd(gnd), .vdd(vdd), .A(_7637_), .B(_7639_), .Y(_7850_) );
OAI21X1 OAI21X1_2180 ( .gnd(gnd), .vdd(vdd), .A(_4953_), .B(_7562__bF_buf1), .C(_7850_), .Y(_7851_) );
XNOR2X1 XNOR2X1_355 ( .gnd(gnd), .vdd(vdd), .A(_7776__bF_buf0), .B(micro_hash_ucr_2_Wx_87_), .Y(_7852_) );
OAI21X1 OAI21X1_2181 ( .gnd(gnd), .vdd(vdd), .A(_7851_), .B(_7852_), .C(micro_hash_ucr_2_pipe28_bF_buf0), .Y(_7853_) );
AOI21X1 AOI21X1_1322 ( .gnd(gnd), .vdd(vdd), .A(_7851_), .B(_7852_), .C(_7853_), .Y(_7854_) );
OAI21X1 OAI21X1_2182 ( .gnd(gnd), .vdd(vdd), .A(_7849_), .B(_7854_), .C(_5110__bF_buf0), .Y(_7855_) );
OAI21X1 OAI21X1_2183 ( .gnd(gnd), .vdd(vdd), .A(_5110__bF_buf3), .B(_7789_), .C(_7855_), .Y(_7856_) );
OAI21X1 OAI21X1_2184 ( .gnd(gnd), .vdd(vdd), .A(_4862_), .B(_7562__bF_buf0), .C(_7653_), .Y(_7857_) );
XNOR2X1 XNOR2X1_356 ( .gnd(gnd), .vdd(vdd), .A(_7776__bF_buf4), .B(_4866_), .Y(_7858_) );
XNOR2X1 XNOR2X1_357 ( .gnd(gnd), .vdd(vdd), .A(_7857_), .B(_7858_), .Y(_7859_) );
MUX2X1 MUX2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_7856_), .B(_7859_), .S(_5111__bF_buf2), .Y(_7860_) );
NOR2X1 NOR2X1_1312 ( .gnd(gnd), .vdd(vdd), .A(_7657_), .B(_7658_), .Y(_7861_) );
AOI21X1 AOI21X1_1323 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_110_), .B(_7561__bF_buf1), .C(_7861_), .Y(_7862_) );
XNOR2X1 XNOR2X1_358 ( .gnd(gnd), .vdd(vdd), .A(_7776__bF_buf3), .B(_4890_), .Y(_7863_) );
AOI21X1 AOI21X1_1324 ( .gnd(gnd), .vdd(vdd), .A(_7863_), .B(_7862_), .C(_5109__bF_buf3), .Y(_7864_) );
OAI21X1 OAI21X1_2185 ( .gnd(gnd), .vdd(vdd), .A(_7862_), .B(_7863_), .C(_7864_), .Y(_7865_) );
OAI21X1 OAI21X1_2186 ( .gnd(gnd), .vdd(vdd), .A(_7860_), .B(micro_hash_ucr_2_pipe34_bF_buf0), .C(_7865_), .Y(_7866_) );
OAI21X1 OAI21X1_2187 ( .gnd(gnd), .vdd(vdd), .A(_4931_), .B(_7562__bF_buf4), .C(_7664_), .Y(_7867_) );
XNOR2X1 XNOR2X1_359 ( .gnd(gnd), .vdd(vdd), .A(_7776__bF_buf2), .B(micro_hash_ucr_2_Wx_119_), .Y(_7868_) );
AND2X2 AND2X2_500 ( .gnd(gnd), .vdd(vdd), .A(_7867_), .B(_7868_), .Y(_7869_) );
OAI21X1 OAI21X1_2188 ( .gnd(gnd), .vdd(vdd), .A(_7867_), .B(_7868_), .C(micro_hash_ucr_2_pipe36_bF_buf0), .Y(_7870_) );
OAI21X1 OAI21X1_2189 ( .gnd(gnd), .vdd(vdd), .A(_7869_), .B(_7870_), .C(_5105__bF_buf2), .Y(_7871_) );
AOI21X1 AOI21X1_1325 ( .gnd(gnd), .vdd(vdd), .A(_5104__bF_buf2), .B(_7866_), .C(_7871_), .Y(_7872_) );
OAI21X1 OAI21X1_2190 ( .gnd(gnd), .vdd(vdd), .A(_4909_), .B(_7562__bF_buf3), .C(_7672_), .Y(_7873_) );
XOR2X1 XOR2X1_151 ( .gnd(gnd), .vdd(vdd), .A(_7776__bF_buf1), .B(micro_hash_ucr_2_Wx_127_), .Y(_7874_) );
XNOR2X1 XNOR2X1_360 ( .gnd(gnd), .vdd(vdd), .A(_7873_), .B(_7874_), .Y(_7875_) );
OAI21X1 OAI21X1_2191 ( .gnd(gnd), .vdd(vdd), .A(_7875_), .B(_5105__bF_buf1), .C(_5103__bF_buf0), .Y(_7876_) );
NOR2X1 NOR2X1_1313 ( .gnd(gnd), .vdd(vdd), .A(_7876_), .B(_7872_), .Y(_7877_) );
OAI21X1 OAI21X1_2192 ( .gnd(gnd), .vdd(vdd), .A(_4805_), .B(_7562__bF_buf2), .C(_7679_), .Y(_7878_) );
XNOR2X1 XNOR2X1_361 ( .gnd(gnd), .vdd(vdd), .A(_7776__bF_buf0), .B(micro_hash_ucr_2_Wx_135_), .Y(_7879_) );
OAI21X1 OAI21X1_2193 ( .gnd(gnd), .vdd(vdd), .A(_7878_), .B(_7879_), .C(micro_hash_ucr_2_pipe40_bF_buf3), .Y(_7880_) );
AOI21X1 AOI21X1_1326 ( .gnd(gnd), .vdd(vdd), .A(_7878_), .B(_7879_), .C(_7880_), .Y(_7881_) );
OAI21X1 OAI21X1_2194 ( .gnd(gnd), .vdd(vdd), .A(_7877_), .B(_7881_), .C(_5098__bF_buf3), .Y(_7882_) );
OAI21X1 OAI21X1_2195 ( .gnd(gnd), .vdd(vdd), .A(_5098__bF_buf2), .B(_7786_), .C(_7882_), .Y(_7883_) );
OAI21X1 OAI21X1_2196 ( .gnd(gnd), .vdd(vdd), .A(_4833_), .B(_7562__bF_buf1), .C(_7690_), .Y(_7884_) );
XNOR2X1 XNOR2X1_362 ( .gnd(gnd), .vdd(vdd), .A(_7776__bF_buf4), .B(_4837_), .Y(_7885_) );
XNOR2X1 XNOR2X1_363 ( .gnd(gnd), .vdd(vdd), .A(_7884_), .B(_7885_), .Y(_7886_) );
MUX2X1 MUX2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_7883_), .B(_7886_), .S(_5099__bF_buf3), .Y(_7887_) );
NOR2X1 NOR2X1_1314 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe46_bF_buf0), .B(_7887_), .Y(_7888_) );
OAI21X1 OAI21X1_2197 ( .gnd(gnd), .vdd(vdd), .A(_4719_), .B(_7562__bF_buf0), .C(_7698_), .Y(_7889_) );
XNOR2X1 XNOR2X1_364 ( .gnd(gnd), .vdd(vdd), .A(_7776__bF_buf3), .B(micro_hash_ucr_2_Wx_159_), .Y(_7890_) );
OAI21X1 OAI21X1_2198 ( .gnd(gnd), .vdd(vdd), .A(_7889_), .B(_7890_), .C(micro_hash_ucr_2_pipe46_bF_buf4), .Y(_7891_) );
AOI21X1 AOI21X1_1327 ( .gnd(gnd), .vdd(vdd), .A(_7889_), .B(_7890_), .C(_7891_), .Y(_7892_) );
OAI21X1 OAI21X1_2199 ( .gnd(gnd), .vdd(vdd), .A(_7888_), .B(_7892_), .C(_5092__bF_buf4), .Y(_7893_) );
OAI21X1 OAI21X1_2200 ( .gnd(gnd), .vdd(vdd), .A(_5092__bF_buf3), .B(_7782_), .C(_7893_), .Y(_7894_) );
OAI21X1 OAI21X1_2201 ( .gnd(gnd), .vdd(vdd), .A(_4747_), .B(_7562__bF_buf4), .C(_7710_), .Y(_7895_) );
XNOR2X1 XNOR2X1_365 ( .gnd(gnd), .vdd(vdd), .A(_7776__bF_buf2), .B(_4751_), .Y(_7896_) );
XNOR2X1 XNOR2X1_366 ( .gnd(gnd), .vdd(vdd), .A(_7895_), .B(_7896_), .Y(_7897_) );
MUX2X1 MUX2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_7894_), .B(_7897_), .S(_5093__bF_buf1), .Y(_7898_) );
AOI21X1 AOI21X1_1328 ( .gnd(gnd), .vdd(vdd), .A(_7565_), .B(_7568_), .C(_7563_), .Y(_7899_) );
XNOR2X1 XNOR2X1_367 ( .gnd(gnd), .vdd(vdd), .A(_7776__bF_buf1), .B(_4809_), .Y(_7900_) );
AOI21X1 AOI21X1_1329 ( .gnd(gnd), .vdd(vdd), .A(_7900_), .B(_7899_), .C(_5091__bF_buf3), .Y(_7901_) );
OAI21X1 OAI21X1_2202 ( .gnd(gnd), .vdd(vdd), .A(_7899_), .B(_7900_), .C(_7901_), .Y(_7902_) );
OAI21X1 OAI21X1_2203 ( .gnd(gnd), .vdd(vdd), .A(_7898_), .B(micro_hash_ucr_2_pipe52_bF_buf3), .C(_7902_), .Y(_7903_) );
OAI21X1 OAI21X1_2204 ( .gnd(gnd), .vdd(vdd), .A(_4863_), .B(_7562__bF_buf3), .C(_7718_), .Y(_7904_) );
XNOR2X1 XNOR2X1_368 ( .gnd(gnd), .vdd(vdd), .A(_7776__bF_buf0), .B(micro_hash_ucr_2_Wx_191_), .Y(_7905_) );
OAI21X1 OAI21X1_2205 ( .gnd(gnd), .vdd(vdd), .A(_7904_), .B(_7905_), .C(micro_hash_ucr_2_pipe54_bF_buf0), .Y(_7906_) );
AOI21X1 AOI21X1_1330 ( .gnd(gnd), .vdd(vdd), .A(_7904_), .B(_7905_), .C(_7906_), .Y(_7907_) );
AOI21X1 AOI21X1_1331 ( .gnd(gnd), .vdd(vdd), .A(_5086__bF_buf2), .B(_7903_), .C(_7907_), .Y(_7908_) );
AOI21X1 AOI21X1_1332 ( .gnd(gnd), .vdd(vdd), .A(_7725_), .B(_7727_), .C(_7723_), .Y(_7909_) );
XNOR2X1 XNOR2X1_369 ( .gnd(gnd), .vdd(vdd), .A(_7776__bF_buf4), .B(micro_hash_ucr_2_Wx_199_), .Y(_7910_) );
AND2X2 AND2X2_501 ( .gnd(gnd), .vdd(vdd), .A(_7909_), .B(_7910_), .Y(_7911_) );
OAI21X1 OAI21X1_2206 ( .gnd(gnd), .vdd(vdd), .A(_7909_), .B(_7910_), .C(micro_hash_ucr_2_pipe56_bF_buf0), .Y(_7912_) );
OAI21X1 OAI21X1_2207 ( .gnd(gnd), .vdd(vdd), .A(_7911_), .B(_7912_), .C(_5085__bF_buf2), .Y(_7913_) );
AOI21X1 AOI21X1_1333 ( .gnd(gnd), .vdd(vdd), .A(_5087__bF_buf2), .B(_7908_), .C(_7913_), .Y(_7914_) );
NAND2X1 NAND2X1_1015 ( .gnd(gnd), .vdd(vdd), .A(_7730_), .B(_7731_), .Y(_7915_) );
OAI21X1 OAI21X1_2208 ( .gnd(gnd), .vdd(vdd), .A(_4720_), .B(_7562__bF_buf2), .C(_7915_), .Y(_7916_) );
XNOR2X1 XNOR2X1_370 ( .gnd(gnd), .vdd(vdd), .A(_7776__bF_buf3), .B(micro_hash_ucr_2_Wx_207_), .Y(_7917_) );
OAI21X1 OAI21X1_2209 ( .gnd(gnd), .vdd(vdd), .A(_7916_), .B(_7917_), .C(micro_hash_ucr_2_pipe58_bF_buf0), .Y(_7918_) );
AOI21X1 AOI21X1_1334 ( .gnd(gnd), .vdd(vdd), .A(_7916_), .B(_7917_), .C(_7918_), .Y(_7919_) );
OAI21X1 OAI21X1_2210 ( .gnd(gnd), .vdd(vdd), .A(_7914_), .B(_7919_), .C(_5080__bF_buf1), .Y(_7920_) );
OAI21X1 OAI21X1_2211 ( .gnd(gnd), .vdd(vdd), .A(_5080__bF_buf0), .B(_7778_), .C(_7920_), .Y(_7921_) );
OAI21X1 OAI21X1_2212 ( .gnd(gnd), .vdd(vdd), .A(_4748_), .B(_7562__bF_buf1), .C(_7742_), .Y(_7922_) );
XNOR2X1 XNOR2X1_371 ( .gnd(gnd), .vdd(vdd), .A(_7776__bF_buf2), .B(micro_hash_ucr_2_Wx_223_), .Y(_7923_) );
OAI21X1 OAI21X1_2213 ( .gnd(gnd), .vdd(vdd), .A(_7922_), .B(_7923_), .C(micro_hash_ucr_2_pipe62_bF_buf2), .Y(_7924_) );
AOI21X1 AOI21X1_1335 ( .gnd(gnd), .vdd(vdd), .A(_7922_), .B(_7923_), .C(_7924_), .Y(_7925_) );
AOI21X1 AOI21X1_1336 ( .gnd(gnd), .vdd(vdd), .A(_5081__bF_buf0), .B(_7921_), .C(_7925_), .Y(_7926_) );
NOR2X1 NOR2X1_1315 ( .gnd(gnd), .vdd(vdd), .A(_7746_), .B(_7562__bF_buf0), .Y(_7927_) );
AOI21X1 AOI21X1_1337 ( .gnd(gnd), .vdd(vdd), .A(_7747_), .B(_7748_), .C(_7927_), .Y(_7928_) );
XOR2X1 XOR2X1_152 ( .gnd(gnd), .vdd(vdd), .A(_7776__bF_buf1), .B(micro_hash_ucr_2_Wx_231_), .Y(_7929_) );
AOI21X1 AOI21X1_1338 ( .gnd(gnd), .vdd(vdd), .A(_7929_), .B(_7928_), .C(_5079__bF_buf3), .Y(_7930_) );
OAI21X1 OAI21X1_2214 ( .gnd(gnd), .vdd(vdd), .A(_7928_), .B(_7929_), .C(_7930_), .Y(_7931_) );
OAI21X1 OAI21X1_2215 ( .gnd(gnd), .vdd(vdd), .A(_7926_), .B(micro_hash_ucr_2_pipe64_bF_buf3), .C(_7931_), .Y(_7932_) );
OAI21X1 OAI21X1_2216 ( .gnd(gnd), .vdd(vdd), .A(_7752_), .B(_7562__bF_buf4), .C(_7756_), .Y(_7933_) );
XNOR2X1 XNOR2X1_372 ( .gnd(gnd), .vdd(vdd), .A(_7776__bF_buf0), .B(micro_hash_ucr_2_Wx_239_), .Y(_7934_) );
OAI21X1 OAI21X1_2217 ( .gnd(gnd), .vdd(vdd), .A(_7933_), .B(_7934_), .C(micro_hash_ucr_2_pipe66_bF_buf2), .Y(_7935_) );
AOI21X1 AOI21X1_1339 ( .gnd(gnd), .vdd(vdd), .A(_7933_), .B(_7934_), .C(_7935_), .Y(_7936_) );
AOI21X1 AOI21X1_1340 ( .gnd(gnd), .vdd(vdd), .A(_5074__bF_buf0), .B(_7932_), .C(_7936_), .Y(_7937_) );
NAND2X1 NAND2X1_1016 ( .gnd(gnd), .vdd(vdd), .A(_7761_), .B(_7763_), .Y(_7938_) );
OAI21X1 OAI21X1_2218 ( .gnd(gnd), .vdd(vdd), .A(_7760_), .B(_7562__bF_buf3), .C(_7938_), .Y(_7939_) );
XOR2X1 XOR2X1_153 ( .gnd(gnd), .vdd(vdd), .A(_7776__bF_buf4), .B(micro_hash_ucr_2_Wx_247_), .Y(_7940_) );
XNOR2X1 XNOR2X1_373 ( .gnd(gnd), .vdd(vdd), .A(_7939_), .B(_7940_), .Y(_7941_) );
OAI21X1 OAI21X1_2219 ( .gnd(gnd), .vdd(vdd), .A(_7941_), .B(_5075__bF_buf2), .C(_5073__bF_buf3), .Y(_7942_) );
AOI21X1 AOI21X1_1341 ( .gnd(gnd), .vdd(vdd), .A(_5075__bF_buf1), .B(_7937_), .C(_7942_), .Y(_7943_) );
NAND2X1 NAND2X1_1017 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_254_), .B(_7561__bF_buf0), .Y(_7944_) );
OAI21X1 OAI21X1_2220 ( .gnd(gnd), .vdd(vdd), .A(_7767_), .B(_7766_), .C(_7944_), .Y(_7945_) );
XNOR2X1 XNOR2X1_374 ( .gnd(gnd), .vdd(vdd), .A(_7776__bF_buf3), .B(micro_hash_ucr_2_Wx_255_), .Y(_7946_) );
AND2X2 AND2X2_502 ( .gnd(gnd), .vdd(vdd), .A(_7945_), .B(_7946_), .Y(_7947_) );
OAI21X1 OAI21X1_2221 ( .gnd(gnd), .vdd(vdd), .A(_7945_), .B(_7946_), .C(micro_hash_ucr_2_pipe69), .Y(_7948_) );
OAI21X1 OAI21X1_2222 ( .gnd(gnd), .vdd(vdd), .A(_7947_), .B(_7948_), .C(_4496__bF_buf6), .Y(_7949_) );
NOR2X1 NOR2X1_1316 ( .gnd(gnd), .vdd(vdd), .A(_7949_), .B(_7943_), .Y(_4493__7_) );
AND2X2 AND2X2_503 ( .gnd(gnd), .vdd(vdd), .A(_5384_), .B(_5494_), .Y(_7950_) );
INVX2 INVX2_253 ( .gnd(gnd), .vdd(vdd), .A(_5151_), .Y(_7951_) );
OAI21X1 OAI21X1_2223 ( .gnd(gnd), .vdd(vdd), .A(_8687_), .B(_6045_), .C(_7951_), .Y(_7952_) );
NOR2X1 NOR2X1_1317 ( .gnd(gnd), .vdd(vdd), .A(_7952_), .B(_7950_), .Y(_7953_) );
AND2X2 AND2X2_504 ( .gnd(gnd), .vdd(vdd), .A(_5272_), .B(_5133_), .Y(_7954_) );
AND2X2 AND2X2_505 ( .gnd(gnd), .vdd(vdd), .A(_7954_), .B(_5493_), .Y(_7955_) );
OAI21X1 OAI21X1_2224 ( .gnd(gnd), .vdd(vdd), .A(_7955_), .B(micro_hash_ucr_2_b_0_bF_buf3_), .C(_5125__bF_buf0), .Y(_7956_) );
OAI21X1 OAI21X1_2225 ( .gnd(gnd), .vdd(vdd), .A(_7953_), .B(_7956_), .C(_5127__bF_buf1), .Y(_7957_) );
AOI21X1 AOI21X1_1342 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe16_bF_buf3), .B(_8690_), .C(micro_hash_ucr_2_pipe17_bF_buf2), .Y(_7958_) );
AOI21X1 AOI21X1_1343 ( .gnd(gnd), .vdd(vdd), .A(_7958_), .B(_7957_), .C(micro_hash_ucr_2_pipe18_bF_buf3), .Y(_7959_) );
OAI21X1 OAI21X1_2226 ( .gnd(gnd), .vdd(vdd), .A(_5122__bF_buf0), .B(micro_hash_ucr_2_b_0_bF_buf2_), .C(_5124__bF_buf2), .Y(_7960_) );
OAI21X1 OAI21X1_2227 ( .gnd(gnd), .vdd(vdd), .A(_7959_), .B(_7960_), .C(_5123__bF_buf4), .Y(_7961_) );
AOI21X1 AOI21X1_1344 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe20_bF_buf0), .B(_8690_), .C(micro_hash_ucr_2_pipe21_bF_buf3), .Y(_7962_) );
AOI21X1 AOI21X1_1345 ( .gnd(gnd), .vdd(vdd), .A(_7962_), .B(_7961_), .C(micro_hash_ucr_2_pipe22_bF_buf1), .Y(_7963_) );
OAI21X1 OAI21X1_2228 ( .gnd(gnd), .vdd(vdd), .A(_5121__bF_buf2), .B(micro_hash_ucr_2_b_0_bF_buf1_), .C(_5120__bF_buf3), .Y(_7964_) );
OAI21X1 OAI21X1_2229 ( .gnd(gnd), .vdd(vdd), .A(_7963_), .B(_7964_), .C(_5116__bF_buf1), .Y(_7965_) );
AOI21X1 AOI21X1_1346 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe24_bF_buf2), .B(_8690_), .C(micro_hash_ucr_2_pipe25), .Y(_7966_) );
AOI21X1 AOI21X1_1347 ( .gnd(gnd), .vdd(vdd), .A(_7966_), .B(_7965_), .C(micro_hash_ucr_2_pipe26_bF_buf2), .Y(_7967_) );
OAI21X1 OAI21X1_2230 ( .gnd(gnd), .vdd(vdd), .A(_5117__bF_buf2), .B(micro_hash_ucr_2_b_0_bF_buf0_), .C(_5113_), .Y(_7968_) );
OAI21X1 OAI21X1_2231 ( .gnd(gnd), .vdd(vdd), .A(_7967_), .B(_7968_), .C(_5115__bF_buf1), .Y(_7969_) );
AOI21X1 AOI21X1_1348 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe28_bF_buf3), .B(_8690_), .C(micro_hash_ucr_2_pipe29_bF_buf1), .Y(_7970_) );
AOI21X1 AOI21X1_1349 ( .gnd(gnd), .vdd(vdd), .A(_7970_), .B(_7969_), .C(micro_hash_ucr_2_pipe30_bF_buf2), .Y(_7971_) );
OAI21X1 OAI21X1_2232 ( .gnd(gnd), .vdd(vdd), .A(_5110__bF_buf2), .B(micro_hash_ucr_2_b_0_bF_buf3_), .C(_5112__bF_buf3), .Y(_7972_) );
OAI21X1 OAI21X1_2233 ( .gnd(gnd), .vdd(vdd), .A(_7971_), .B(_7972_), .C(_5111__bF_buf1), .Y(_7973_) );
AOI21X1 AOI21X1_1350 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe32_bF_buf1), .B(_8690_), .C(micro_hash_ucr_2_pipe33_bF_buf0), .Y(_7974_) );
AOI21X1 AOI21X1_1351 ( .gnd(gnd), .vdd(vdd), .A(_7974_), .B(_7973_), .C(micro_hash_ucr_2_pipe34_bF_buf3), .Y(_7975_) );
OAI21X1 OAI21X1_2234 ( .gnd(gnd), .vdd(vdd), .A(_5109__bF_buf2), .B(micro_hash_ucr_2_b_0_bF_buf2_), .C(_5108__bF_buf2), .Y(_7976_) );
OAI21X1 OAI21X1_2235 ( .gnd(gnd), .vdd(vdd), .A(_7975_), .B(_7976_), .C(_5104__bF_buf1), .Y(_7977_) );
AOI21X1 AOI21X1_1352 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe36_bF_buf3), .B(_8690_), .C(micro_hash_ucr_2_pipe37), .Y(_7978_) );
AOI21X1 AOI21X1_1353 ( .gnd(gnd), .vdd(vdd), .A(_7978_), .B(_7977_), .C(micro_hash_ucr_2_pipe38_bF_buf0), .Y(_7979_) );
OAI21X1 OAI21X1_2236 ( .gnd(gnd), .vdd(vdd), .A(_5105__bF_buf0), .B(micro_hash_ucr_2_b_0_bF_buf1_), .C(_5101_), .Y(_7980_) );
OAI21X1 OAI21X1_2237 ( .gnd(gnd), .vdd(vdd), .A(_7979_), .B(_7980_), .C(_5103__bF_buf3), .Y(_7981_) );
AOI21X1 AOI21X1_1354 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe40_bF_buf2), .B(_8690_), .C(micro_hash_ucr_2_pipe41_bF_buf1), .Y(_7982_) );
AOI21X1 AOI21X1_1355 ( .gnd(gnd), .vdd(vdd), .A(_7982_), .B(_7981_), .C(micro_hash_ucr_2_pipe42_bF_buf3), .Y(_7983_) );
OAI21X1 OAI21X1_2238 ( .gnd(gnd), .vdd(vdd), .A(_5098__bF_buf1), .B(micro_hash_ucr_2_b_0_bF_buf0_), .C(_5100__bF_buf0), .Y(_7984_) );
OAI21X1 OAI21X1_2239 ( .gnd(gnd), .vdd(vdd), .A(_7983_), .B(_7984_), .C(_5099__bF_buf2), .Y(_7985_) );
AOI21X1 AOI21X1_1356 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe44_bF_buf0), .B(_8690_), .C(micro_hash_ucr_2_pipe45_bF_buf0), .Y(_7986_) );
AOI21X1 AOI21X1_1357 ( .gnd(gnd), .vdd(vdd), .A(_7986_), .B(_7985_), .C(micro_hash_ucr_2_pipe46_bF_buf3), .Y(_7987_) );
OAI21X1 OAI21X1_2240 ( .gnd(gnd), .vdd(vdd), .A(_5097__bF_buf2), .B(micro_hash_ucr_2_b_0_bF_buf3_), .C(_5096__bF_buf3), .Y(_7988_) );
OAI21X1 OAI21X1_2241 ( .gnd(gnd), .vdd(vdd), .A(_7987_), .B(_7988_), .C(_5092__bF_buf2), .Y(_7989_) );
AOI21X1 AOI21X1_1358 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe48_bF_buf2), .B(_8690_), .C(micro_hash_ucr_2_pipe49_bF_buf0), .Y(_7990_) );
AOI21X1 AOI21X1_1359 ( .gnd(gnd), .vdd(vdd), .A(_7990_), .B(_7989_), .C(micro_hash_ucr_2_pipe50_bF_buf1), .Y(_7991_) );
OAI21X1 OAI21X1_2242 ( .gnd(gnd), .vdd(vdd), .A(_5093__bF_buf0), .B(micro_hash_ucr_2_b_0_bF_buf2_), .C(_5089__bF_buf3), .Y(_7992_) );
OAI21X1 OAI21X1_2243 ( .gnd(gnd), .vdd(vdd), .A(_7991_), .B(_7992_), .C(_5091__bF_buf2), .Y(_7993_) );
AOI21X1 AOI21X1_1360 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe52_bF_buf2), .B(_8690_), .C(micro_hash_ucr_2_pipe53_bF_buf1), .Y(_7994_) );
AOI21X1 AOI21X1_1361 ( .gnd(gnd), .vdd(vdd), .A(_7994_), .B(_7993_), .C(micro_hash_ucr_2_pipe54_bF_buf4), .Y(_7995_) );
OAI21X1 OAI21X1_2244 ( .gnd(gnd), .vdd(vdd), .A(_5086__bF_buf1), .B(micro_hash_ucr_2_b_0_bF_buf1_), .C(_5088_), .Y(_7996_) );
OAI21X1 OAI21X1_2245 ( .gnd(gnd), .vdd(vdd), .A(_7995_), .B(_7996_), .C(_5087__bF_buf1), .Y(_7997_) );
AOI21X1 AOI21X1_1362 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe56_bF_buf3), .B(_8690_), .C(micro_hash_ucr_2_pipe57_bF_buf1), .Y(_7998_) );
AOI21X1 AOI21X1_1363 ( .gnd(gnd), .vdd(vdd), .A(_7998_), .B(_7997_), .C(micro_hash_ucr_2_pipe58_bF_buf4), .Y(_7999_) );
OAI21X1 OAI21X1_2246 ( .gnd(gnd), .vdd(vdd), .A(_5085__bF_buf1), .B(micro_hash_ucr_2_b_0_bF_buf0_), .C(_5084__bF_buf3), .Y(_8000_) );
OAI21X1 OAI21X1_2247 ( .gnd(gnd), .vdd(vdd), .A(_7999_), .B(_8000_), .C(_5080__bF_buf3), .Y(_8001_) );
AOI21X1 AOI21X1_1364 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe60_bF_buf1), .B(_8690_), .C(micro_hash_ucr_2_pipe61_bF_buf0), .Y(_8002_) );
AOI21X1 AOI21X1_1365 ( .gnd(gnd), .vdd(vdd), .A(_8002_), .B(_8001_), .C(micro_hash_ucr_2_pipe62_bF_buf1), .Y(_8003_) );
OAI21X1 OAI21X1_2248 ( .gnd(gnd), .vdd(vdd), .A(_5081__bF_buf3), .B(micro_hash_ucr_2_b_0_bF_buf3_), .C(_5077__bF_buf2), .Y(_8004_) );
OAI21X1 OAI21X1_2249 ( .gnd(gnd), .vdd(vdd), .A(_8003_), .B(_8004_), .C(_5079__bF_buf2), .Y(_8005_) );
AOI21X1 AOI21X1_1366 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe64_bF_buf2), .B(_8690_), .C(micro_hash_ucr_2_pipe65_bF_buf2), .Y(_8006_) );
AOI21X1 AOI21X1_1367 ( .gnd(gnd), .vdd(vdd), .A(_8006_), .B(_8005_), .C(micro_hash_ucr_2_pipe66_bF_buf1), .Y(_8007_) );
OAI21X1 OAI21X1_2250 ( .gnd(gnd), .vdd(vdd), .A(_5074__bF_buf3), .B(micro_hash_ucr_2_b_0_bF_buf2_), .C(_5076__bF_buf1), .Y(_8008_) );
OAI21X1 OAI21X1_2251 ( .gnd(gnd), .vdd(vdd), .A(_8007_), .B(_8008_), .C(_5075__bF_buf0), .Y(_8009_) );
OAI21X1 OAI21X1_2252 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_0_bF_buf1_), .B(_5075__bF_buf4), .C(_8009_), .Y(_8010_) );
NOR2X1 NOR2X1_1318 ( .gnd(gnd), .vdd(vdd), .A(_6147_), .B(_8010_), .Y(_4492__0_) );
OAI21X1 OAI21X1_2253 ( .gnd(gnd), .vdd(vdd), .A(_8694_), .B(_6045_), .C(_7951_), .Y(_8011_) );
NOR2X1 NOR2X1_1319 ( .gnd(gnd), .vdd(vdd), .A(_8011_), .B(_7950_), .Y(_8012_) );
OAI21X1 OAI21X1_2254 ( .gnd(gnd), .vdd(vdd), .A(_7955_), .B(micro_hash_ucr_2_b_1_bF_buf3_), .C(_5125__bF_buf3), .Y(_8013_) );
OAI21X1 OAI21X1_2255 ( .gnd(gnd), .vdd(vdd), .A(_8012_), .B(_8013_), .C(_5127__bF_buf0), .Y(_8014_) );
AOI21X1 AOI21X1_1368 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe16_bF_buf2), .B(_8696_), .C(micro_hash_ucr_2_pipe17_bF_buf1), .Y(_8015_) );
AOI21X1 AOI21X1_1369 ( .gnd(gnd), .vdd(vdd), .A(_8015_), .B(_8014_), .C(micro_hash_ucr_2_pipe18_bF_buf2), .Y(_8016_) );
OAI21X1 OAI21X1_2256 ( .gnd(gnd), .vdd(vdd), .A(_5122__bF_buf4), .B(micro_hash_ucr_2_b_1_bF_buf2_), .C(_5124__bF_buf1), .Y(_8017_) );
OAI21X1 OAI21X1_2257 ( .gnd(gnd), .vdd(vdd), .A(_8016_), .B(_8017_), .C(_5123__bF_buf3), .Y(_8018_) );
AOI21X1 AOI21X1_1370 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe20_bF_buf3), .B(_8696_), .C(micro_hash_ucr_2_pipe21_bF_buf2), .Y(_8019_) );
AOI21X1 AOI21X1_1371 ( .gnd(gnd), .vdd(vdd), .A(_8019_), .B(_8018_), .C(micro_hash_ucr_2_pipe22_bF_buf0), .Y(_8020_) );
OAI21X1 OAI21X1_2258 ( .gnd(gnd), .vdd(vdd), .A(_5121__bF_buf1), .B(micro_hash_ucr_2_b_1_bF_buf1_), .C(_5120__bF_buf2), .Y(_8021_) );
OAI21X1 OAI21X1_2259 ( .gnd(gnd), .vdd(vdd), .A(_8020_), .B(_8021_), .C(_5116__bF_buf0), .Y(_8022_) );
AOI21X1 AOI21X1_1372 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe24_bF_buf1), .B(_8696_), .C(micro_hash_ucr_2_pipe25), .Y(_8023_) );
AOI21X1 AOI21X1_1373 ( .gnd(gnd), .vdd(vdd), .A(_8023_), .B(_8022_), .C(micro_hash_ucr_2_pipe26_bF_buf1), .Y(_8024_) );
OAI21X1 OAI21X1_2260 ( .gnd(gnd), .vdd(vdd), .A(_5117__bF_buf1), .B(micro_hash_ucr_2_b_1_bF_buf0_), .C(_5113_), .Y(_8025_) );
OAI21X1 OAI21X1_2261 ( .gnd(gnd), .vdd(vdd), .A(_8024_), .B(_8025_), .C(_5115__bF_buf0), .Y(_8026_) );
AOI21X1 AOI21X1_1374 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe28_bF_buf2), .B(_8696_), .C(micro_hash_ucr_2_pipe29_bF_buf0), .Y(_8027_) );
AOI21X1 AOI21X1_1375 ( .gnd(gnd), .vdd(vdd), .A(_8027_), .B(_8026_), .C(micro_hash_ucr_2_pipe30_bF_buf1), .Y(_8028_) );
OAI21X1 OAI21X1_2262 ( .gnd(gnd), .vdd(vdd), .A(_5110__bF_buf1), .B(micro_hash_ucr_2_b_1_bF_buf3_), .C(_5112__bF_buf2), .Y(_8029_) );
OAI21X1 OAI21X1_2263 ( .gnd(gnd), .vdd(vdd), .A(_8028_), .B(_8029_), .C(_5111__bF_buf0), .Y(_8030_) );
AOI21X1 AOI21X1_1376 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe32_bF_buf0), .B(_8696_), .C(micro_hash_ucr_2_pipe33_bF_buf3), .Y(_8031_) );
AOI21X1 AOI21X1_1377 ( .gnd(gnd), .vdd(vdd), .A(_8031_), .B(_8030_), .C(micro_hash_ucr_2_pipe34_bF_buf2), .Y(_8032_) );
OAI21X1 OAI21X1_2264 ( .gnd(gnd), .vdd(vdd), .A(_5109__bF_buf1), .B(micro_hash_ucr_2_b_1_bF_buf2_), .C(_5108__bF_buf1), .Y(_8033_) );
OAI21X1 OAI21X1_2265 ( .gnd(gnd), .vdd(vdd), .A(_8032_), .B(_8033_), .C(_5104__bF_buf0), .Y(_8034_) );
AOI21X1 AOI21X1_1378 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe36_bF_buf2), .B(_8696_), .C(micro_hash_ucr_2_pipe37), .Y(_8035_) );
AOI21X1 AOI21X1_1379 ( .gnd(gnd), .vdd(vdd), .A(_8035_), .B(_8034_), .C(micro_hash_ucr_2_pipe38_bF_buf3), .Y(_8036_) );
OAI21X1 OAI21X1_2266 ( .gnd(gnd), .vdd(vdd), .A(_5105__bF_buf4), .B(micro_hash_ucr_2_b_1_bF_buf1_), .C(_5101_), .Y(_8037_) );
OAI21X1 OAI21X1_2267 ( .gnd(gnd), .vdd(vdd), .A(_8036_), .B(_8037_), .C(_5103__bF_buf2), .Y(_8038_) );
AOI21X1 AOI21X1_1380 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe40_bF_buf1), .B(_8696_), .C(micro_hash_ucr_2_pipe41_bF_buf0), .Y(_8039_) );
AOI21X1 AOI21X1_1381 ( .gnd(gnd), .vdd(vdd), .A(_8039_), .B(_8038_), .C(micro_hash_ucr_2_pipe42_bF_buf2), .Y(_8040_) );
OAI21X1 OAI21X1_2268 ( .gnd(gnd), .vdd(vdd), .A(_5098__bF_buf0), .B(micro_hash_ucr_2_b_1_bF_buf0_), .C(_5100__bF_buf3), .Y(_8041_) );
OAI21X1 OAI21X1_2269 ( .gnd(gnd), .vdd(vdd), .A(_8040_), .B(_8041_), .C(_5099__bF_buf1), .Y(_8042_) );
AOI21X1 AOI21X1_1382 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe44_bF_buf3), .B(_8696_), .C(micro_hash_ucr_2_pipe45_bF_buf3), .Y(_8043_) );
AOI21X1 AOI21X1_1383 ( .gnd(gnd), .vdd(vdd), .A(_8043_), .B(_8042_), .C(micro_hash_ucr_2_pipe46_bF_buf2), .Y(_8044_) );
OAI21X1 OAI21X1_2270 ( .gnd(gnd), .vdd(vdd), .A(_5097__bF_buf1), .B(micro_hash_ucr_2_b_1_bF_buf3_), .C(_5096__bF_buf2), .Y(_8045_) );
OAI21X1 OAI21X1_2271 ( .gnd(gnd), .vdd(vdd), .A(_8044_), .B(_8045_), .C(_5092__bF_buf1), .Y(_8046_) );
AOI21X1 AOI21X1_1384 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe48_bF_buf1), .B(_8696_), .C(micro_hash_ucr_2_pipe49_bF_buf3), .Y(_8047_) );
AOI21X1 AOI21X1_1385 ( .gnd(gnd), .vdd(vdd), .A(_8047_), .B(_8046_), .C(micro_hash_ucr_2_pipe50_bF_buf0), .Y(_8048_) );
OAI21X1 OAI21X1_2272 ( .gnd(gnd), .vdd(vdd), .A(_5093__bF_buf4), .B(micro_hash_ucr_2_b_1_bF_buf2_), .C(_5089__bF_buf2), .Y(_8049_) );
OAI21X1 OAI21X1_2273 ( .gnd(gnd), .vdd(vdd), .A(_8048_), .B(_8049_), .C(_5091__bF_buf1), .Y(_8050_) );
AOI21X1 AOI21X1_1386 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe52_bF_buf1), .B(_8696_), .C(micro_hash_ucr_2_pipe53_bF_buf0), .Y(_8051_) );
AOI21X1 AOI21X1_1387 ( .gnd(gnd), .vdd(vdd), .A(_8051_), .B(_8050_), .C(micro_hash_ucr_2_pipe54_bF_buf3), .Y(_8052_) );
OAI21X1 OAI21X1_2274 ( .gnd(gnd), .vdd(vdd), .A(_5086__bF_buf0), .B(micro_hash_ucr_2_b_1_bF_buf1_), .C(_5088_), .Y(_8053_) );
OAI21X1 OAI21X1_2275 ( .gnd(gnd), .vdd(vdd), .A(_8052_), .B(_8053_), .C(_5087__bF_buf0), .Y(_8054_) );
AOI21X1 AOI21X1_1388 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe56_bF_buf2), .B(_8696_), .C(micro_hash_ucr_2_pipe57_bF_buf0), .Y(_8055_) );
AOI21X1 AOI21X1_1389 ( .gnd(gnd), .vdd(vdd), .A(_8055_), .B(_8054_), .C(micro_hash_ucr_2_pipe58_bF_buf3), .Y(_8056_) );
OAI21X1 OAI21X1_2276 ( .gnd(gnd), .vdd(vdd), .A(_5085__bF_buf0), .B(micro_hash_ucr_2_b_1_bF_buf0_), .C(_5084__bF_buf2), .Y(_8057_) );
OAI21X1 OAI21X1_2277 ( .gnd(gnd), .vdd(vdd), .A(_8056_), .B(_8057_), .C(_5080__bF_buf2), .Y(_8058_) );
AOI21X1 AOI21X1_1390 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe60_bF_buf0), .B(_8696_), .C(micro_hash_ucr_2_pipe61_bF_buf3), .Y(_8059_) );
AOI21X1 AOI21X1_1391 ( .gnd(gnd), .vdd(vdd), .A(_8059_), .B(_8058_), .C(micro_hash_ucr_2_pipe62_bF_buf0), .Y(_8060_) );
OAI21X1 OAI21X1_2278 ( .gnd(gnd), .vdd(vdd), .A(_5081__bF_buf2), .B(micro_hash_ucr_2_b_1_bF_buf3_), .C(_5077__bF_buf1), .Y(_8061_) );
OAI21X1 OAI21X1_2279 ( .gnd(gnd), .vdd(vdd), .A(_8060_), .B(_8061_), .C(_5079__bF_buf1), .Y(_8062_) );
AOI21X1 AOI21X1_1392 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe64_bF_buf1), .B(_8696_), .C(micro_hash_ucr_2_pipe65_bF_buf1), .Y(_8063_) );
AOI21X1 AOI21X1_1393 ( .gnd(gnd), .vdd(vdd), .A(_8063_), .B(_8062_), .C(micro_hash_ucr_2_pipe66_bF_buf0), .Y(_8064_) );
OAI21X1 OAI21X1_2280 ( .gnd(gnd), .vdd(vdd), .A(_5074__bF_buf2), .B(micro_hash_ucr_2_b_1_bF_buf2_), .C(_5076__bF_buf0), .Y(_8065_) );
OAI21X1 OAI21X1_2281 ( .gnd(gnd), .vdd(vdd), .A(_8064_), .B(_8065_), .C(_5075__bF_buf3), .Y(_8066_) );
OAI21X1 OAI21X1_2282 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_1_bF_buf1_), .B(_5075__bF_buf2), .C(_8066_), .Y(_8067_) );
NOR2X1 NOR2X1_1320 ( .gnd(gnd), .vdd(vdd), .A(_6147_), .B(_8067_), .Y(_4492__1_) );
OAI21X1 OAI21X1_2283 ( .gnd(gnd), .vdd(vdd), .A(_4573_), .B(_6045_), .C(_7951_), .Y(_8068_) );
NOR2X1 NOR2X1_1321 ( .gnd(gnd), .vdd(vdd), .A(_8068_), .B(_7950_), .Y(_8069_) );
OAI21X1 OAI21X1_2284 ( .gnd(gnd), .vdd(vdd), .A(_7955_), .B(micro_hash_ucr_2_b_2_bF_buf2_), .C(_5125__bF_buf2), .Y(_8070_) );
OAI21X1 OAI21X1_2285 ( .gnd(gnd), .vdd(vdd), .A(_8069_), .B(_8070_), .C(_5127__bF_buf3), .Y(_8071_) );
AOI21X1 AOI21X1_1394 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe16_bF_buf1), .B(_4583_), .C(micro_hash_ucr_2_pipe17_bF_buf0), .Y(_8072_) );
AOI21X1 AOI21X1_1395 ( .gnd(gnd), .vdd(vdd), .A(_8072_), .B(_8071_), .C(micro_hash_ucr_2_pipe18_bF_buf1), .Y(_8073_) );
OAI21X1 OAI21X1_2286 ( .gnd(gnd), .vdd(vdd), .A(_5122__bF_buf3), .B(micro_hash_ucr_2_b_2_bF_buf1_), .C(_5124__bF_buf0), .Y(_8074_) );
OAI21X1 OAI21X1_2287 ( .gnd(gnd), .vdd(vdd), .A(_8073_), .B(_8074_), .C(_5123__bF_buf2), .Y(_8075_) );
AOI21X1 AOI21X1_1396 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe20_bF_buf2), .B(_4583_), .C(micro_hash_ucr_2_pipe21_bF_buf1), .Y(_8076_) );
AOI21X1 AOI21X1_1397 ( .gnd(gnd), .vdd(vdd), .A(_8076_), .B(_8075_), .C(micro_hash_ucr_2_pipe22_bF_buf4), .Y(_8077_) );
OAI21X1 OAI21X1_2288 ( .gnd(gnd), .vdd(vdd), .A(_5121__bF_buf0), .B(micro_hash_ucr_2_b_2_bF_buf0_), .C(_5120__bF_buf1), .Y(_8078_) );
OAI21X1 OAI21X1_2289 ( .gnd(gnd), .vdd(vdd), .A(_8077_), .B(_8078_), .C(_5116__bF_buf4), .Y(_8079_) );
AOI21X1 AOI21X1_1398 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe24_bF_buf0), .B(_4583_), .C(micro_hash_ucr_2_pipe25), .Y(_8080_) );
AOI21X1 AOI21X1_1399 ( .gnd(gnd), .vdd(vdd), .A(_8080_), .B(_8079_), .C(micro_hash_ucr_2_pipe26_bF_buf0), .Y(_8081_) );
OAI21X1 OAI21X1_2290 ( .gnd(gnd), .vdd(vdd), .A(_5117__bF_buf0), .B(micro_hash_ucr_2_b_2_bF_buf3_), .C(_5113_), .Y(_8082_) );
OAI21X1 OAI21X1_2291 ( .gnd(gnd), .vdd(vdd), .A(_8081_), .B(_8082_), .C(_5115__bF_buf4), .Y(_8083_) );
AOI21X1 AOI21X1_1400 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe28_bF_buf1), .B(_4583_), .C(micro_hash_ucr_2_pipe29_bF_buf3), .Y(_8084_) );
AOI21X1 AOI21X1_1401 ( .gnd(gnd), .vdd(vdd), .A(_8084_), .B(_8083_), .C(micro_hash_ucr_2_pipe30_bF_buf0), .Y(_8085_) );
OAI21X1 OAI21X1_2292 ( .gnd(gnd), .vdd(vdd), .A(_5110__bF_buf0), .B(micro_hash_ucr_2_b_2_bF_buf2_), .C(_5112__bF_buf1), .Y(_8086_) );
OAI21X1 OAI21X1_2293 ( .gnd(gnd), .vdd(vdd), .A(_8085_), .B(_8086_), .C(_5111__bF_buf4), .Y(_8087_) );
AOI21X1 AOI21X1_1402 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe32_bF_buf3), .B(_4583_), .C(micro_hash_ucr_2_pipe33_bF_buf2), .Y(_8088_) );
AOI21X1 AOI21X1_1403 ( .gnd(gnd), .vdd(vdd), .A(_8088_), .B(_8087_), .C(micro_hash_ucr_2_pipe34_bF_buf1), .Y(_8089_) );
OAI21X1 OAI21X1_2294 ( .gnd(gnd), .vdd(vdd), .A(_5109__bF_buf0), .B(micro_hash_ucr_2_b_2_bF_buf1_), .C(_5108__bF_buf0), .Y(_8090_) );
OAI21X1 OAI21X1_2295 ( .gnd(gnd), .vdd(vdd), .A(_8089_), .B(_8090_), .C(_5104__bF_buf4), .Y(_8091_) );
AOI21X1 AOI21X1_1404 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe36_bF_buf1), .B(_4583_), .C(micro_hash_ucr_2_pipe37), .Y(_8092_) );
AOI21X1 AOI21X1_1405 ( .gnd(gnd), .vdd(vdd), .A(_8092_), .B(_8091_), .C(micro_hash_ucr_2_pipe38_bF_buf2), .Y(_8093_) );
OAI21X1 OAI21X1_2296 ( .gnd(gnd), .vdd(vdd), .A(_5105__bF_buf3), .B(micro_hash_ucr_2_b_2_bF_buf0_), .C(_5101_), .Y(_8094_) );
OAI21X1 OAI21X1_2297 ( .gnd(gnd), .vdd(vdd), .A(_8093_), .B(_8094_), .C(_5103__bF_buf1), .Y(_8095_) );
AOI21X1 AOI21X1_1406 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe40_bF_buf0), .B(_4583_), .C(micro_hash_ucr_2_pipe41_bF_buf3), .Y(_8096_) );
AOI21X1 AOI21X1_1407 ( .gnd(gnd), .vdd(vdd), .A(_8096_), .B(_8095_), .C(micro_hash_ucr_2_pipe42_bF_buf1), .Y(_8097_) );
OAI21X1 OAI21X1_2298 ( .gnd(gnd), .vdd(vdd), .A(_5098__bF_buf4), .B(micro_hash_ucr_2_b_2_bF_buf3_), .C(_5100__bF_buf2), .Y(_8098_) );
OAI21X1 OAI21X1_2299 ( .gnd(gnd), .vdd(vdd), .A(_8097_), .B(_8098_), .C(_5099__bF_buf0), .Y(_8099_) );
AOI21X1 AOI21X1_1408 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe44_bF_buf2), .B(_4583_), .C(micro_hash_ucr_2_pipe45_bF_buf2), .Y(_8100_) );
AOI21X1 AOI21X1_1409 ( .gnd(gnd), .vdd(vdd), .A(_8100_), .B(_8099_), .C(micro_hash_ucr_2_pipe46_bF_buf1), .Y(_8101_) );
OAI21X1 OAI21X1_2300 ( .gnd(gnd), .vdd(vdd), .A(_5097__bF_buf0), .B(micro_hash_ucr_2_b_2_bF_buf2_), .C(_5096__bF_buf1), .Y(_8102_) );
OAI21X1 OAI21X1_2301 ( .gnd(gnd), .vdd(vdd), .A(_8101_), .B(_8102_), .C(_5092__bF_buf0), .Y(_8103_) );
AOI21X1 AOI21X1_1410 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe48_bF_buf0), .B(_4583_), .C(micro_hash_ucr_2_pipe49_bF_buf2), .Y(_8104_) );
AOI21X1 AOI21X1_1411 ( .gnd(gnd), .vdd(vdd), .A(_8104_), .B(_8103_), .C(micro_hash_ucr_2_pipe50_bF_buf3), .Y(_8105_) );
OAI21X1 OAI21X1_2302 ( .gnd(gnd), .vdd(vdd), .A(_5093__bF_buf3), .B(micro_hash_ucr_2_b_2_bF_buf1_), .C(_5089__bF_buf1), .Y(_8106_) );
OAI21X1 OAI21X1_2303 ( .gnd(gnd), .vdd(vdd), .A(_8105_), .B(_8106_), .C(_5091__bF_buf0), .Y(_8107_) );
AOI21X1 AOI21X1_1412 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe52_bF_buf0), .B(_4583_), .C(micro_hash_ucr_2_pipe53_bF_buf3), .Y(_8108_) );
AOI21X1 AOI21X1_1413 ( .gnd(gnd), .vdd(vdd), .A(_8108_), .B(_8107_), .C(micro_hash_ucr_2_pipe54_bF_buf2), .Y(_8109_) );
OAI21X1 OAI21X1_2304 ( .gnd(gnd), .vdd(vdd), .A(_5086__bF_buf3), .B(micro_hash_ucr_2_b_2_bF_buf0_), .C(_5088_), .Y(_8110_) );
OAI21X1 OAI21X1_2305 ( .gnd(gnd), .vdd(vdd), .A(_8109_), .B(_8110_), .C(_5087__bF_buf4), .Y(_8111_) );
AOI21X1 AOI21X1_1414 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe56_bF_buf1), .B(_4583_), .C(micro_hash_ucr_2_pipe57_bF_buf3), .Y(_8112_) );
AOI21X1 AOI21X1_1415 ( .gnd(gnd), .vdd(vdd), .A(_8112_), .B(_8111_), .C(micro_hash_ucr_2_pipe58_bF_buf2), .Y(_8113_) );
OAI21X1 OAI21X1_2306 ( .gnd(gnd), .vdd(vdd), .A(_5085__bF_buf3), .B(micro_hash_ucr_2_b_2_bF_buf3_), .C(_5084__bF_buf1), .Y(_8114_) );
OAI21X1 OAI21X1_2307 ( .gnd(gnd), .vdd(vdd), .A(_8113_), .B(_8114_), .C(_5080__bF_buf1), .Y(_8115_) );
AOI21X1 AOI21X1_1416 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe60_bF_buf4), .B(_4583_), .C(micro_hash_ucr_2_pipe61_bF_buf2), .Y(_8116_) );
AOI21X1 AOI21X1_1417 ( .gnd(gnd), .vdd(vdd), .A(_8116_), .B(_8115_), .C(micro_hash_ucr_2_pipe62_bF_buf4), .Y(_8117_) );
OAI21X1 OAI21X1_2308 ( .gnd(gnd), .vdd(vdd), .A(_5081__bF_buf1), .B(micro_hash_ucr_2_b_2_bF_buf2_), .C(_5077__bF_buf0), .Y(_8118_) );
OAI21X1 OAI21X1_2309 ( .gnd(gnd), .vdd(vdd), .A(_8117_), .B(_8118_), .C(_5079__bF_buf0), .Y(_8119_) );
AOI21X1 AOI21X1_1418 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe64_bF_buf0), .B(_4583_), .C(micro_hash_ucr_2_pipe65_bF_buf0), .Y(_8120_) );
AOI21X1 AOI21X1_1419 ( .gnd(gnd), .vdd(vdd), .A(_8120_), .B(_8119_), .C(micro_hash_ucr_2_pipe66_bF_buf4), .Y(_8121_) );
OAI21X1 OAI21X1_2310 ( .gnd(gnd), .vdd(vdd), .A(_5074__bF_buf1), .B(micro_hash_ucr_2_b_2_bF_buf1_), .C(_5076__bF_buf3), .Y(_8122_) );
OAI21X1 OAI21X1_2311 ( .gnd(gnd), .vdd(vdd), .A(_8121_), .B(_8122_), .C(_5075__bF_buf1), .Y(_8123_) );
OAI21X1 OAI21X1_2312 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_2_bF_buf0_), .B(_5075__bF_buf0), .C(_8123_), .Y(_8124_) );
NOR2X1 NOR2X1_1322 ( .gnd(gnd), .vdd(vdd), .A(_6147_), .B(_8124_), .Y(_4492__2_) );
OAI21X1 OAI21X1_2313 ( .gnd(gnd), .vdd(vdd), .A(_4587_), .B(_6045_), .C(_7951_), .Y(_8125_) );
NOR2X1 NOR2X1_1323 ( .gnd(gnd), .vdd(vdd), .A(_8125_), .B(_7950_), .Y(_8126_) );
OAI21X1 OAI21X1_2314 ( .gnd(gnd), .vdd(vdd), .A(_7955_), .B(micro_hash_ucr_2_b_3_bF_buf2_), .C(_5125__bF_buf1), .Y(_8127_) );
OAI21X1 OAI21X1_2315 ( .gnd(gnd), .vdd(vdd), .A(_8126_), .B(_8127_), .C(_5127__bF_buf2), .Y(_8128_) );
AOI21X1 AOI21X1_1420 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe16_bF_buf0), .B(_4588_), .C(micro_hash_ucr_2_pipe17_bF_buf3), .Y(_8129_) );
AOI21X1 AOI21X1_1421 ( .gnd(gnd), .vdd(vdd), .A(_8129_), .B(_8128_), .C(micro_hash_ucr_2_pipe18_bF_buf0), .Y(_8130_) );
OAI21X1 OAI21X1_2316 ( .gnd(gnd), .vdd(vdd), .A(_5122__bF_buf2), .B(micro_hash_ucr_2_b_3_bF_buf1_), .C(_5124__bF_buf3), .Y(_8131_) );
OAI21X1 OAI21X1_2317 ( .gnd(gnd), .vdd(vdd), .A(_8130_), .B(_8131_), .C(_5123__bF_buf1), .Y(_8132_) );
AOI21X1 AOI21X1_1422 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe20_bF_buf1), .B(_4588_), .C(micro_hash_ucr_2_pipe21_bF_buf0), .Y(_8133_) );
AOI21X1 AOI21X1_1423 ( .gnd(gnd), .vdd(vdd), .A(_8133_), .B(_8132_), .C(micro_hash_ucr_2_pipe22_bF_buf3), .Y(_8134_) );
OAI21X1 OAI21X1_2318 ( .gnd(gnd), .vdd(vdd), .A(_5121__bF_buf4), .B(micro_hash_ucr_2_b_3_bF_buf0_), .C(_5120__bF_buf0), .Y(_8135_) );
OAI21X1 OAI21X1_2319 ( .gnd(gnd), .vdd(vdd), .A(_8134_), .B(_8135_), .C(_5116__bF_buf3), .Y(_8136_) );
AOI21X1 AOI21X1_1424 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe24_bF_buf3), .B(_4588_), .C(micro_hash_ucr_2_pipe25), .Y(_8137_) );
AOI21X1 AOI21X1_1425 ( .gnd(gnd), .vdd(vdd), .A(_8137_), .B(_8136_), .C(micro_hash_ucr_2_pipe26_bF_buf3), .Y(_8138_) );
OAI21X1 OAI21X1_2320 ( .gnd(gnd), .vdd(vdd), .A(_5117__bF_buf4), .B(micro_hash_ucr_2_b_3_bF_buf3_), .C(_5113_), .Y(_8139_) );
OAI21X1 OAI21X1_2321 ( .gnd(gnd), .vdd(vdd), .A(_8138_), .B(_8139_), .C(_5115__bF_buf3), .Y(_8140_) );
AOI21X1 AOI21X1_1426 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe28_bF_buf0), .B(_4588_), .C(micro_hash_ucr_2_pipe29_bF_buf2), .Y(_8141_) );
AOI21X1 AOI21X1_1427 ( .gnd(gnd), .vdd(vdd), .A(_8141_), .B(_8140_), .C(micro_hash_ucr_2_pipe30_bF_buf4), .Y(_8142_) );
OAI21X1 OAI21X1_2322 ( .gnd(gnd), .vdd(vdd), .A(_5110__bF_buf3), .B(micro_hash_ucr_2_b_3_bF_buf2_), .C(_5112__bF_buf0), .Y(_8143_) );
OAI21X1 OAI21X1_2323 ( .gnd(gnd), .vdd(vdd), .A(_8142_), .B(_8143_), .C(_5111__bF_buf3), .Y(_8144_) );
AOI21X1 AOI21X1_1428 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe32_bF_buf2), .B(_4588_), .C(micro_hash_ucr_2_pipe33_bF_buf1), .Y(_8145_) );
AOI21X1 AOI21X1_1429 ( .gnd(gnd), .vdd(vdd), .A(_8145_), .B(_8144_), .C(micro_hash_ucr_2_pipe34_bF_buf0), .Y(_8146_) );
OAI21X1 OAI21X1_2324 ( .gnd(gnd), .vdd(vdd), .A(_5109__bF_buf4), .B(micro_hash_ucr_2_b_3_bF_buf1_), .C(_5108__bF_buf3), .Y(_8147_) );
OAI21X1 OAI21X1_2325 ( .gnd(gnd), .vdd(vdd), .A(_8146_), .B(_8147_), .C(_5104__bF_buf3), .Y(_8148_) );
AOI21X1 AOI21X1_1430 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe36_bF_buf0), .B(_4588_), .C(micro_hash_ucr_2_pipe37), .Y(_8149_) );
AOI21X1 AOI21X1_1431 ( .gnd(gnd), .vdd(vdd), .A(_8149_), .B(_8148_), .C(micro_hash_ucr_2_pipe38_bF_buf1), .Y(_8150_) );
OAI21X1 OAI21X1_2326 ( .gnd(gnd), .vdd(vdd), .A(_5105__bF_buf2), .B(micro_hash_ucr_2_b_3_bF_buf0_), .C(_5101_), .Y(_8151_) );
OAI21X1 OAI21X1_2327 ( .gnd(gnd), .vdd(vdd), .A(_8150_), .B(_8151_), .C(_5103__bF_buf0), .Y(_8152_) );
AOI21X1 AOI21X1_1432 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe40_bF_buf4), .B(_4588_), .C(micro_hash_ucr_2_pipe41_bF_buf2), .Y(_8153_) );
AOI21X1 AOI21X1_1433 ( .gnd(gnd), .vdd(vdd), .A(_8153_), .B(_8152_), .C(micro_hash_ucr_2_pipe42_bF_buf0), .Y(_8154_) );
OAI21X1 OAI21X1_2328 ( .gnd(gnd), .vdd(vdd), .A(_5098__bF_buf3), .B(micro_hash_ucr_2_b_3_bF_buf3_), .C(_5100__bF_buf1), .Y(_8155_) );
OAI21X1 OAI21X1_2329 ( .gnd(gnd), .vdd(vdd), .A(_8154_), .B(_8155_), .C(_5099__bF_buf4), .Y(_8156_) );
AOI21X1 AOI21X1_1434 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe44_bF_buf1), .B(_4588_), .C(micro_hash_ucr_2_pipe45_bF_buf1), .Y(_8157_) );
AOI21X1 AOI21X1_1435 ( .gnd(gnd), .vdd(vdd), .A(_8157_), .B(_8156_), .C(micro_hash_ucr_2_pipe46_bF_buf0), .Y(_8158_) );
OAI21X1 OAI21X1_2330 ( .gnd(gnd), .vdd(vdd), .A(_5097__bF_buf3), .B(micro_hash_ucr_2_b_3_bF_buf2_), .C(_5096__bF_buf0), .Y(_8159_) );
OAI21X1 OAI21X1_2331 ( .gnd(gnd), .vdd(vdd), .A(_8158_), .B(_8159_), .C(_5092__bF_buf4), .Y(_8160_) );
AOI21X1 AOI21X1_1436 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe48_bF_buf4), .B(_4588_), .C(micro_hash_ucr_2_pipe49_bF_buf1), .Y(_8161_) );
AOI21X1 AOI21X1_1437 ( .gnd(gnd), .vdd(vdd), .A(_8161_), .B(_8160_), .C(micro_hash_ucr_2_pipe50_bF_buf2), .Y(_8162_) );
OAI21X1 OAI21X1_2332 ( .gnd(gnd), .vdd(vdd), .A(_5093__bF_buf2), .B(micro_hash_ucr_2_b_3_bF_buf1_), .C(_5089__bF_buf0), .Y(_8163_) );
OAI21X1 OAI21X1_2333 ( .gnd(gnd), .vdd(vdd), .A(_8162_), .B(_8163_), .C(_5091__bF_buf4), .Y(_8164_) );
AOI21X1 AOI21X1_1438 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe52_bF_buf3), .B(_4588_), .C(micro_hash_ucr_2_pipe53_bF_buf2), .Y(_8165_) );
AOI21X1 AOI21X1_1439 ( .gnd(gnd), .vdd(vdd), .A(_8165_), .B(_8164_), .C(micro_hash_ucr_2_pipe54_bF_buf1), .Y(_8166_) );
OAI21X1 OAI21X1_2334 ( .gnd(gnd), .vdd(vdd), .A(_5086__bF_buf2), .B(micro_hash_ucr_2_b_3_bF_buf0_), .C(_5088_), .Y(_8167_) );
OAI21X1 OAI21X1_2335 ( .gnd(gnd), .vdd(vdd), .A(_8166_), .B(_8167_), .C(_5087__bF_buf3), .Y(_8168_) );
AOI21X1 AOI21X1_1440 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe56_bF_buf0), .B(_4588_), .C(micro_hash_ucr_2_pipe57_bF_buf2), .Y(_8169_) );
AOI21X1 AOI21X1_1441 ( .gnd(gnd), .vdd(vdd), .A(_8169_), .B(_8168_), .C(micro_hash_ucr_2_pipe58_bF_buf1), .Y(_8170_) );
OAI21X1 OAI21X1_2336 ( .gnd(gnd), .vdd(vdd), .A(_5085__bF_buf2), .B(micro_hash_ucr_2_b_3_bF_buf3_), .C(_5084__bF_buf0), .Y(_8171_) );
OAI21X1 OAI21X1_2337 ( .gnd(gnd), .vdd(vdd), .A(_8170_), .B(_8171_), .C(_5080__bF_buf0), .Y(_8172_) );
AOI21X1 AOI21X1_1442 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe60_bF_buf3), .B(_4588_), .C(micro_hash_ucr_2_pipe61_bF_buf1), .Y(_8173_) );
AOI21X1 AOI21X1_1443 ( .gnd(gnd), .vdd(vdd), .A(_8173_), .B(_8172_), .C(micro_hash_ucr_2_pipe62_bF_buf3), .Y(_8174_) );
OAI21X1 OAI21X1_2338 ( .gnd(gnd), .vdd(vdd), .A(_5081__bF_buf0), .B(micro_hash_ucr_2_b_3_bF_buf2_), .C(_5077__bF_buf3), .Y(_8175_) );
OAI21X1 OAI21X1_2339 ( .gnd(gnd), .vdd(vdd), .A(_8174_), .B(_8175_), .C(_5079__bF_buf4), .Y(_8176_) );
AOI21X1 AOI21X1_1444 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe64_bF_buf4), .B(_4588_), .C(micro_hash_ucr_2_pipe65_bF_buf3), .Y(_8177_) );
AOI21X1 AOI21X1_1445 ( .gnd(gnd), .vdd(vdd), .A(_8177_), .B(_8176_), .C(micro_hash_ucr_2_pipe66_bF_buf3), .Y(_8178_) );
OAI21X1 OAI21X1_2340 ( .gnd(gnd), .vdd(vdd), .A(_5074__bF_buf0), .B(micro_hash_ucr_2_b_3_bF_buf1_), .C(_5076__bF_buf2), .Y(_8179_) );
OAI21X1 OAI21X1_2341 ( .gnd(gnd), .vdd(vdd), .A(_8178_), .B(_8179_), .C(_5075__bF_buf4), .Y(_8180_) );
OAI21X1 OAI21X1_2342 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_3_bF_buf0_), .B(_5075__bF_buf3), .C(_8180_), .Y(_8181_) );
NOR2X1 NOR2X1_1324 ( .gnd(gnd), .vdd(vdd), .A(_6147_), .B(_8181_), .Y(_4492__3_) );
NAND2X1 NAND2X1_1018 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_0_bF_buf3_), .B(_4563_), .Y(_8182_) );
NAND2X1 NAND2X1_1019 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_4_bF_buf2_), .B(micro_hash_ucr_2_pipe66_bF_buf2), .Y(_8183_) );
NAND2X1 NAND2X1_1020 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe65_bF_buf2), .B(_8632__bF_buf0), .Y(_8184_) );
NAND2X1 NAND2X1_1021 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_4_bF_buf1_), .B(micro_hash_ucr_2_pipe64_bF_buf3), .Y(_8185_) );
NAND2X1 NAND2X1_1022 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe63), .B(_8632__bF_buf3), .Y(_8186_) );
NAND2X1 NAND2X1_1023 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe52_bF_buf2), .B(_5593_), .Y(_8187_) );
NAND2X1 NAND2X1_1024 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_0_bF_buf2_), .B(micro_hash_ucr_2_pipe51), .Y(_8188_) );
NAND2X1 NAND2X1_1025 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe50_bF_buf1), .B(_5593_), .Y(_8189_) );
NAND2X1 NAND2X1_1026 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_0_bF_buf1_), .B(micro_hash_ucr_2_pipe49_bF_buf0), .Y(_8190_) );
NAND2X1 NAND2X1_1027 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe48_bF_buf3), .B(_5593_), .Y(_8191_) );
NAND2X1 NAND2X1_1028 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_0_bF_buf0_), .B(micro_hash_ucr_2_pipe47), .Y(_8192_) );
NOR2X1 NOR2X1_1325 ( .gnd(gnd), .vdd(vdd), .A(_5593_), .B(_5097__bF_buf2), .Y(_8193_) );
NAND2X1 NAND2X1_1029 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_0_bF_buf3_), .B(micro_hash_ucr_2_pipe45_bF_buf0), .Y(_8194_) );
NAND2X1 NAND2X1_1030 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe29_bF_buf1), .B(_8632__bF_buf2), .Y(_8195_) );
NOR2X1 NOR2X1_1326 ( .gnd(gnd), .vdd(vdd), .A(_8632__bF_buf1), .B(_5120__bF_buf3), .Y(_8196_) );
NAND2X1 NAND2X1_1031 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_4_bF_buf0_), .B(micro_hash_ucr_2_pipe22_bF_buf2), .Y(_8197_) );
NOR2X1 NOR2X1_1327 ( .gnd(gnd), .vdd(vdd), .A(_8632__bF_buf0), .B(_5119_), .Y(_8198_) );
NAND2X1 NAND2X1_1032 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_4_bF_buf3_), .B(micro_hash_ucr_2_pipe20_bF_buf0), .Y(_8199_) );
NOR2X1 NOR2X1_1328 ( .gnd(gnd), .vdd(vdd), .A(_8632__bF_buf3), .B(_5124__bF_buf2), .Y(_8200_) );
NAND2X1 NAND2X1_1033 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_4_bF_buf2_), .B(micro_hash_ucr_2_pipe18_bF_buf4), .Y(_8201_) );
NOR2X1 NOR2X1_1329 ( .gnd(gnd), .vdd(vdd), .A(_8632__bF_buf2), .B(_5126_), .Y(_8202_) );
NAND2X1 NAND2X1_1034 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_4_bF_buf1_), .B(micro_hash_ucr_2_pipe16_bF_buf4), .Y(_8203_) );
NAND2X1 NAND2X1_1035 ( .gnd(gnd), .vdd(vdd), .A(_8632__bF_buf1), .B(_5270_), .Y(_8204_) );
NAND2X1 NAND2X1_1036 ( .gnd(gnd), .vdd(vdd), .A(_4599_), .B(_5128_), .Y(_8205_) );
NAND2X1 NAND2X1_1037 ( .gnd(gnd), .vdd(vdd), .A(_5132_), .B(_5133_), .Y(_8206_) );
NOR2X1 NOR2X1_1330 ( .gnd(gnd), .vdd(vdd), .A(_8205_), .B(_8206_), .Y(_8207_) );
NOR2X1 NOR2X1_1331 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe14_bF_buf2), .B(micro_hash_ucr_2_pipe13), .Y(_8208_) );
NAND3X1 NAND3X1_324 ( .gnd(gnd), .vdd(vdd), .A(_5168_), .B(_8208_), .C(_8207_), .Y(_8209_) );
OAI22X1 OAI22X1_105 ( .gnd(gnd), .vdd(vdd), .A(_5158_), .B(_8209_), .C(_5278_), .D(micro_hash_ucr_2_b_4_bF_buf0_), .Y(_8210_) );
AOI21X1 AOI21X1_1446 ( .gnd(gnd), .vdd(vdd), .A(_5125__bF_buf0), .B(_8210_), .C(micro_hash_ucr_2_pipe16_bF_buf3), .Y(_8211_) );
NAND2X1 NAND2X1_1038 ( .gnd(gnd), .vdd(vdd), .A(_8204_), .B(_8211_), .Y(_8212_) );
AOI21X1 AOI21X1_1447 ( .gnd(gnd), .vdd(vdd), .A(_8203_), .B(_8212_), .C(micro_hash_ucr_2_pipe17_bF_buf2), .Y(_8213_) );
OAI21X1 OAI21X1_2343 ( .gnd(gnd), .vdd(vdd), .A(_8213_), .B(_8202_), .C(_5122__bF_buf1), .Y(_8214_) );
AOI21X1 AOI21X1_1448 ( .gnd(gnd), .vdd(vdd), .A(_8201_), .B(_8214_), .C(micro_hash_ucr_2_pipe19), .Y(_8215_) );
OAI21X1 OAI21X1_2344 ( .gnd(gnd), .vdd(vdd), .A(_8215_), .B(_8200_), .C(_5123__bF_buf0), .Y(_8216_) );
AOI21X1 AOI21X1_1449 ( .gnd(gnd), .vdd(vdd), .A(_8199_), .B(_8216_), .C(micro_hash_ucr_2_pipe21_bF_buf3), .Y(_8217_) );
OAI21X1 OAI21X1_2345 ( .gnd(gnd), .vdd(vdd), .A(_8217_), .B(_8198_), .C(_5121__bF_buf3), .Y(_8218_) );
AOI21X1 AOI21X1_1450 ( .gnd(gnd), .vdd(vdd), .A(_8197_), .B(_8218_), .C(micro_hash_ucr_2_pipe23), .Y(_8219_) );
OAI21X1 OAI21X1_2346 ( .gnd(gnd), .vdd(vdd), .A(_8219_), .B(_8196_), .C(_5116__bF_buf2), .Y(_8220_) );
OAI21X1 OAI21X1_2347 ( .gnd(gnd), .vdd(vdd), .A(_5593_), .B(_5116__bF_buf1), .C(_8220_), .Y(_8221_) );
NAND2X1 NAND2X1_1039 ( .gnd(gnd), .vdd(vdd), .A(_5118__bF_buf0), .B(_8221_), .Y(_8222_) );
OAI21X1 OAI21X1_2348 ( .gnd(gnd), .vdd(vdd), .A(_8632__bF_buf0), .B(_5118__bF_buf3), .C(_8222_), .Y(_8223_) );
AOI21X1 AOI21X1_1451 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe26_bF_buf2), .B(_5593_), .C(micro_hash_ucr_2_pipe27), .Y(_8224_) );
OAI21X1 OAI21X1_2349 ( .gnd(gnd), .vdd(vdd), .A(_8223_), .B(micro_hash_ucr_2_pipe26_bF_buf1), .C(_8224_), .Y(_8225_) );
AOI21X1 AOI21X1_1452 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_0_bF_buf2_), .B(micro_hash_ucr_2_pipe27), .C(micro_hash_ucr_2_pipe28_bF_buf3), .Y(_8226_) );
AND2X2 AND2X2_506 ( .gnd(gnd), .vdd(vdd), .A(_8225_), .B(_8226_), .Y(_8227_) );
NOR2X1 NOR2X1_1332 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_4_bF_buf3_), .B(_5115__bF_buf2), .Y(_8228_) );
OAI21X1 OAI21X1_2350 ( .gnd(gnd), .vdd(vdd), .A(_8227_), .B(_8228_), .C(_5114_), .Y(_8229_) );
NAND3X1 NAND3X1_325 ( .gnd(gnd), .vdd(vdd), .A(_5110__bF_buf2), .B(_8195_), .C(_8229_), .Y(_8230_) );
AOI21X1 AOI21X1_1453 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_4_bF_buf2_), .B(micro_hash_ucr_2_pipe30_bF_buf3), .C(micro_hash_ucr_2_pipe31), .Y(_8231_) );
OAI21X1 OAI21X1_2351 ( .gnd(gnd), .vdd(vdd), .A(_5112__bF_buf3), .B(micro_hash_ucr_2_c_0_bF_buf1_), .C(_5111__bF_buf2), .Y(_8232_) );
AOI21X1 AOI21X1_1454 ( .gnd(gnd), .vdd(vdd), .A(_8231_), .B(_8230_), .C(_8232_), .Y(_8233_) );
NOR2X1 NOR2X1_1333 ( .gnd(gnd), .vdd(vdd), .A(_5593_), .B(_5111__bF_buf1), .Y(_8234_) );
OAI21X1 OAI21X1_2352 ( .gnd(gnd), .vdd(vdd), .A(_8233_), .B(_8234_), .C(_5107_), .Y(_8235_) );
AOI21X1 AOI21X1_1455 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_0_bF_buf0_), .B(micro_hash_ucr_2_pipe33_bF_buf0), .C(micro_hash_ucr_2_pipe34_bF_buf3), .Y(_8236_) );
OAI21X1 OAI21X1_2353 ( .gnd(gnd), .vdd(vdd), .A(_5109__bF_buf3), .B(micro_hash_ucr_2_b_4_bF_buf1_), .C(_5108__bF_buf2), .Y(_8237_) );
AOI21X1 AOI21X1_1456 ( .gnd(gnd), .vdd(vdd), .A(_8236_), .B(_8235_), .C(_8237_), .Y(_8238_) );
OAI21X1 OAI21X1_2354 ( .gnd(gnd), .vdd(vdd), .A(_8632__bF_buf3), .B(_5108__bF_buf1), .C(_5104__bF_buf2), .Y(_8239_) );
OAI22X1 OAI22X1_106 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_4_bF_buf0_), .B(_5104__bF_buf1), .C(_8238_), .D(_8239_), .Y(_8240_) );
OAI21X1 OAI21X1_2355 ( .gnd(gnd), .vdd(vdd), .A(_5106_), .B(micro_hash_ucr_2_c_0_bF_buf3_), .C(_5105__bF_buf1), .Y(_8241_) );
AOI21X1 AOI21X1_1457 ( .gnd(gnd), .vdd(vdd), .A(_5106_), .B(_8240_), .C(_8241_), .Y(_8242_) );
NOR2X1 NOR2X1_1334 ( .gnd(gnd), .vdd(vdd), .A(_5593_), .B(_5105__bF_buf0), .Y(_8243_) );
OAI21X1 OAI21X1_2356 ( .gnd(gnd), .vdd(vdd), .A(_8242_), .B(_8243_), .C(_5101_), .Y(_8244_) );
AOI21X1 AOI21X1_1458 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_0_bF_buf2_), .B(micro_hash_ucr_2_pipe39), .C(micro_hash_ucr_2_pipe40_bF_buf3), .Y(_8245_) );
OAI21X1 OAI21X1_2357 ( .gnd(gnd), .vdd(vdd), .A(_5103__bF_buf3), .B(micro_hash_ucr_2_b_4_bF_buf3_), .C(_5102_), .Y(_8246_) );
AOI21X1 AOI21X1_1459 ( .gnd(gnd), .vdd(vdd), .A(_8245_), .B(_8244_), .C(_8246_), .Y(_8247_) );
OAI21X1 OAI21X1_2358 ( .gnd(gnd), .vdd(vdd), .A(_8632__bF_buf2), .B(_5102_), .C(_5098__bF_buf2), .Y(_8248_) );
OAI22X1 OAI22X1_107 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_4_bF_buf2_), .B(_5098__bF_buf1), .C(_8247_), .D(_8248_), .Y(_8249_) );
OAI21X1 OAI21X1_2359 ( .gnd(gnd), .vdd(vdd), .A(_5100__bF_buf0), .B(micro_hash_ucr_2_c_0_bF_buf1_), .C(_5099__bF_buf3), .Y(_8250_) );
AOI21X1 AOI21X1_1460 ( .gnd(gnd), .vdd(vdd), .A(_5100__bF_buf3), .B(_8249_), .C(_8250_), .Y(_8251_) );
NOR2X1 NOR2X1_1335 ( .gnd(gnd), .vdd(vdd), .A(_5593_), .B(_5099__bF_buf2), .Y(_8252_) );
OAI21X1 OAI21X1_2360 ( .gnd(gnd), .vdd(vdd), .A(_8251_), .B(_8252_), .C(_5095_), .Y(_8253_) );
AOI21X1 AOI21X1_1461 ( .gnd(gnd), .vdd(vdd), .A(_8194_), .B(_8253_), .C(micro_hash_ucr_2_pipe46_bF_buf4), .Y(_8254_) );
OAI21X1 OAI21X1_2361 ( .gnd(gnd), .vdd(vdd), .A(_8254_), .B(_8193_), .C(_5096__bF_buf3), .Y(_8255_) );
NAND3X1 NAND3X1_326 ( .gnd(gnd), .vdd(vdd), .A(_5092__bF_buf3), .B(_8192_), .C(_8255_), .Y(_8256_) );
NAND3X1 NAND3X1_327 ( .gnd(gnd), .vdd(vdd), .A(_5094_), .B(_8191_), .C(_8256_), .Y(_8257_) );
NAND3X1 NAND3X1_328 ( .gnd(gnd), .vdd(vdd), .A(_5093__bF_buf1), .B(_8190_), .C(_8257_), .Y(_8258_) );
NAND3X1 NAND3X1_329 ( .gnd(gnd), .vdd(vdd), .A(_5089__bF_buf3), .B(_8189_), .C(_8258_), .Y(_8259_) );
NAND3X1 NAND3X1_330 ( .gnd(gnd), .vdd(vdd), .A(_5091__bF_buf3), .B(_8188_), .C(_8259_), .Y(_8260_) );
NAND3X1 NAND3X1_331 ( .gnd(gnd), .vdd(vdd), .A(_5090_), .B(_8187_), .C(_8260_), .Y(_8261_) );
AOI21X1 AOI21X1_1462 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_0_bF_buf0_), .B(micro_hash_ucr_2_pipe53_bF_buf1), .C(micro_hash_ucr_2_pipe54_bF_buf0), .Y(_8262_) );
OAI21X1 OAI21X1_2362 ( .gnd(gnd), .vdd(vdd), .A(_5086__bF_buf1), .B(micro_hash_ucr_2_b_4_bF_buf1_), .C(_5088_), .Y(_8263_) );
AOI21X1 AOI21X1_1463 ( .gnd(gnd), .vdd(vdd), .A(_8262_), .B(_8261_), .C(_8263_), .Y(_8264_) );
OAI21X1 OAI21X1_2363 ( .gnd(gnd), .vdd(vdd), .A(_8632__bF_buf1), .B(_5088_), .C(_5087__bF_buf2), .Y(_8265_) );
NAND2X1 NAND2X1_1040 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe56_bF_buf3), .B(_5593_), .Y(_8266_) );
OAI21X1 OAI21X1_2364 ( .gnd(gnd), .vdd(vdd), .A(_8264_), .B(_8265_), .C(_8266_), .Y(_8267_) );
NAND2X1 NAND2X1_1041 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_0_bF_buf3_), .B(micro_hash_ucr_2_pipe57_bF_buf1), .Y(_8268_) );
OAI21X1 OAI21X1_2365 ( .gnd(gnd), .vdd(vdd), .A(_8267_), .B(micro_hash_ucr_2_pipe57_bF_buf0), .C(_8268_), .Y(_8269_) );
AOI21X1 AOI21X1_1464 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe58_bF_buf0), .B(_5593_), .C(micro_hash_ucr_2_pipe59), .Y(_8270_) );
OAI21X1 OAI21X1_2366 ( .gnd(gnd), .vdd(vdd), .A(_8269_), .B(micro_hash_ucr_2_pipe58_bF_buf4), .C(_8270_), .Y(_8271_) );
AOI21X1 AOI21X1_1465 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_0_bF_buf2_), .B(micro_hash_ucr_2_pipe59), .C(micro_hash_ucr_2_pipe60_bF_buf2), .Y(_8272_) );
AOI22X1 AOI22X1_60 ( .gnd(gnd), .vdd(vdd), .A(_5593_), .B(micro_hash_ucr_2_pipe60_bF_buf1), .C(_8271_), .D(_8272_), .Y(_8273_) );
AOI21X1 AOI21X1_1466 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe61_bF_buf0), .B(_8632__bF_buf0), .C(micro_hash_ucr_2_pipe62_bF_buf2), .Y(_8274_) );
OAI21X1 OAI21X1_2367 ( .gnd(gnd), .vdd(vdd), .A(_8273_), .B(micro_hash_ucr_2_pipe61_bF_buf3), .C(_8274_), .Y(_8275_) );
NAND2X1 NAND2X1_1042 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_4_bF_buf0_), .B(micro_hash_ucr_2_pipe62_bF_buf1), .Y(_8276_) );
NAND3X1 NAND3X1_332 ( .gnd(gnd), .vdd(vdd), .A(_5077__bF_buf2), .B(_8276_), .C(_8275_), .Y(_8277_) );
NAND3X1 NAND3X1_333 ( .gnd(gnd), .vdd(vdd), .A(_5079__bF_buf3), .B(_8186_), .C(_8277_), .Y(_8278_) );
NAND3X1 NAND3X1_334 ( .gnd(gnd), .vdd(vdd), .A(_5078_), .B(_8185_), .C(_8278_), .Y(_8279_) );
NAND3X1 NAND3X1_335 ( .gnd(gnd), .vdd(vdd), .A(_5074__bF_buf3), .B(_8184_), .C(_8279_), .Y(_8280_) );
NAND2X1 NAND2X1_1043 ( .gnd(gnd), .vdd(vdd), .A(_8183_), .B(_8280_), .Y(_8281_) );
OAI21X1 OAI21X1_2368 ( .gnd(gnd), .vdd(vdd), .A(_8632__bF_buf3), .B(_5076__bF_buf1), .C(_5075__bF_buf2), .Y(_8282_) );
AOI21X1 AOI21X1_1467 ( .gnd(gnd), .vdd(vdd), .A(_5076__bF_buf0), .B(_8281_), .C(_8282_), .Y(_8283_) );
OAI21X1 OAI21X1_2369 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_4_bF_buf3_), .B(_5075__bF_buf1), .C(_6146_), .Y(_8284_) );
OAI21X1 OAI21X1_2370 ( .gnd(gnd), .vdd(vdd), .A(_8283_), .B(_8284_), .C(_8182_), .Y(_4492__4_) );
NAND2X1 NAND2X1_1044 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_1_bF_buf3_), .B(_4563_), .Y(_8285_) );
NAND2X1 NAND2X1_1045 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe64_bF_buf2), .B(_4608__bF_buf2), .Y(_8286_) );
NAND2X1 NAND2X1_1046 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_1_bF_buf2_), .B(micro_hash_ucr_2_pipe63), .Y(_8287_) );
NAND2X1 NAND2X1_1047 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe62_bF_buf0), .B(_4608__bF_buf1), .Y(_8288_) );
NAND2X1 NAND2X1_1048 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_1_bF_buf1_), .B(micro_hash_ucr_2_pipe61_bF_buf2), .Y(_8289_) );
NAND2X1 NAND2X1_1049 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe60_bF_buf0), .B(_4608__bF_buf0), .Y(_8290_) );
NAND2X1 NAND2X1_1050 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_1_bF_buf0_), .B(micro_hash_ucr_2_pipe59), .Y(_8291_) );
NAND2X1 NAND2X1_1051 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe58_bF_buf3), .B(_4608__bF_buf3), .Y(_8292_) );
NAND2X1 NAND2X1_1052 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_1_bF_buf3_), .B(micro_hash_ucr_2_pipe57_bF_buf3), .Y(_8293_) );
NAND2X1 NAND2X1_1053 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe56_bF_buf2), .B(_4608__bF_buf2), .Y(_8294_) );
NAND2X1 NAND2X1_1054 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_1_bF_buf2_), .B(micro_hash_ucr_2_pipe55), .Y(_8295_) );
NAND2X1 NAND2X1_1055 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe54_bF_buf4), .B(_4608__bF_buf1), .Y(_8296_) );
NAND2X1 NAND2X1_1056 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_1_bF_buf1_), .B(micro_hash_ucr_2_pipe53_bF_buf0), .Y(_8297_) );
NAND2X1 NAND2X1_1057 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe52_bF_buf1), .B(_4608__bF_buf0), .Y(_8298_) );
NAND2X1 NAND2X1_1058 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_1_bF_buf0_), .B(micro_hash_ucr_2_pipe51), .Y(_8299_) );
NAND2X1 NAND2X1_1059 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_1_bF_buf3_), .B(micro_hash_ucr_2_pipe43), .Y(_8300_) );
NAND2X1 NAND2X1_1060 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_5_bF_buf1_), .B(micro_hash_ucr_2_pipe36_bF_buf3), .Y(_8301_) );
NAND2X1 NAND2X1_1061 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe35), .B(_5255_), .Y(_8302_) );
NAND2X1 NAND2X1_1062 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_5_bF_buf0_), .B(micro_hash_ucr_2_pipe34_bF_buf2), .Y(_8303_) );
NAND2X1 NAND2X1_1063 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe33_bF_buf3), .B(_5255_), .Y(_8304_) );
NAND2X1 NAND2X1_1064 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_5_bF_buf3_), .B(micro_hash_ucr_2_pipe32_bF_buf1), .Y(_8305_) );
NAND2X1 NAND2X1_1065 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe31), .B(_5255_), .Y(_8306_) );
NAND2X1 NAND2X1_1066 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_1_bF_buf2_), .B(micro_hash_ucr_2_pipe27), .Y(_8307_) );
NAND2X1 NAND2X1_1067 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_5_bF_buf2_), .B(micro_hash_ucr_2_pipe16_bF_buf2), .Y(_8308_) );
NAND2X1 NAND2X1_1068 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_5_bF_buf1_), .B(micro_hash_ucr_2_pipe14_bF_buf1), .Y(_8309_) );
NAND2X1 NAND2X1_1069 ( .gnd(gnd), .vdd(vdd), .A(_5131_), .B(_5383_), .Y(_8310_) );
NOR2X1 NOR2X1_1336 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe10), .B(micro_hash_ucr_2_pipe7), .Y(_8311_) );
NAND3X1 NAND3X1_336 ( .gnd(gnd), .vdd(vdd), .A(_4607_), .B(_5132_), .C(_8311_), .Y(_8312_) );
OAI22X1 OAI22X1_108 ( .gnd(gnd), .vdd(vdd), .A(_8310_), .B(_8312_), .C(_5172_), .D(micro_hash_ucr_2_c_1_bF_buf1_), .Y(_8313_) );
NAND2X1 NAND2X1_1070 ( .gnd(gnd), .vdd(vdd), .A(_5128_), .B(_8313_), .Y(_8314_) );
AOI21X1 AOI21X1_1468 ( .gnd(gnd), .vdd(vdd), .A(_4608__bF_buf3), .B(_5160_), .C(micro_hash_ucr_2_pipe13), .Y(_8315_) );
AOI22X1 AOI22X1_61 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_1_bF_buf0_), .B(micro_hash_ucr_2_pipe13), .C(_8315_), .D(_8314_), .Y(_8316_) );
OAI21X1 OAI21X1_2371 ( .gnd(gnd), .vdd(vdd), .A(_8316_), .B(micro_hash_ucr_2_pipe14_bF_buf0), .C(_8309_), .Y(_8317_) );
NAND2X1 NAND2X1_1071 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe15), .B(_5255_), .Y(_8318_) );
OAI21X1 OAI21X1_2372 ( .gnd(gnd), .vdd(vdd), .A(_8317_), .B(micro_hash_ucr_2_pipe15), .C(_8318_), .Y(_8319_) );
OAI21X1 OAI21X1_2373 ( .gnd(gnd), .vdd(vdd), .A(_8319_), .B(micro_hash_ucr_2_pipe16_bF_buf1), .C(_8308_), .Y(_8320_) );
NAND2X1 NAND2X1_1072 ( .gnd(gnd), .vdd(vdd), .A(_5126_), .B(_8320_), .Y(_8321_) );
OAI21X1 OAI21X1_2374 ( .gnd(gnd), .vdd(vdd), .A(_5255_), .B(_5126_), .C(_8321_), .Y(_8322_) );
AOI21X1 AOI21X1_1469 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe18_bF_buf3), .B(_4608__bF_buf2), .C(micro_hash_ucr_2_pipe19), .Y(_8323_) );
OAI21X1 OAI21X1_2375 ( .gnd(gnd), .vdd(vdd), .A(_8322_), .B(micro_hash_ucr_2_pipe18_bF_buf2), .C(_8323_), .Y(_8324_) );
OAI21X1 OAI21X1_2376 ( .gnd(gnd), .vdd(vdd), .A(_5255_), .B(_5124__bF_buf1), .C(_8324_), .Y(_8325_) );
NAND2X1 NAND2X1_1073 ( .gnd(gnd), .vdd(vdd), .A(_5123__bF_buf4), .B(_8325_), .Y(_8326_) );
OAI21X1 OAI21X1_2377 ( .gnd(gnd), .vdd(vdd), .A(_4608__bF_buf1), .B(_5123__bF_buf3), .C(_8326_), .Y(_8327_) );
NAND2X1 NAND2X1_1074 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe21_bF_buf2), .B(_5255_), .Y(_8328_) );
OAI21X1 OAI21X1_2378 ( .gnd(gnd), .vdd(vdd), .A(_8327_), .B(micro_hash_ucr_2_pipe21_bF_buf1), .C(_8328_), .Y(_8329_) );
OAI21X1 OAI21X1_2379 ( .gnd(gnd), .vdd(vdd), .A(_5121__bF_buf2), .B(micro_hash_ucr_2_b_5_bF_buf0_), .C(_5120__bF_buf2), .Y(_8330_) );
AOI21X1 AOI21X1_1470 ( .gnd(gnd), .vdd(vdd), .A(_5121__bF_buf1), .B(_8329_), .C(_8330_), .Y(_8331_) );
OAI21X1 OAI21X1_2380 ( .gnd(gnd), .vdd(vdd), .A(_5255_), .B(_5120__bF_buf1), .C(_5116__bF_buf0), .Y(_8332_) );
OAI22X1 OAI22X1_109 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_5_bF_buf3_), .B(_5116__bF_buf4), .C(_8331_), .D(_8332_), .Y(_8333_) );
OAI21X1 OAI21X1_2381 ( .gnd(gnd), .vdd(vdd), .A(_5118__bF_buf2), .B(micro_hash_ucr_2_c_1_bF_buf3_), .C(_5117__bF_buf3), .Y(_8334_) );
AOI21X1 AOI21X1_1471 ( .gnd(gnd), .vdd(vdd), .A(_5118__bF_buf1), .B(_8333_), .C(_8334_), .Y(_8335_) );
NOR2X1 NOR2X1_1337 ( .gnd(gnd), .vdd(vdd), .A(_4608__bF_buf0), .B(_5117__bF_buf2), .Y(_8336_) );
OAI21X1 OAI21X1_2382 ( .gnd(gnd), .vdd(vdd), .A(_8335_), .B(_8336_), .C(_5113_), .Y(_8337_) );
AOI21X1 AOI21X1_1472 ( .gnd(gnd), .vdd(vdd), .A(_8307_), .B(_8337_), .C(micro_hash_ucr_2_pipe28_bF_buf2), .Y(_8338_) );
OAI21X1 OAI21X1_2383 ( .gnd(gnd), .vdd(vdd), .A(_4608__bF_buf3), .B(_5115__bF_buf1), .C(_5114_), .Y(_8339_) );
AOI21X1 AOI21X1_1473 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe29_bF_buf0), .B(_5255_), .C(micro_hash_ucr_2_pipe30_bF_buf2), .Y(_8340_) );
OAI21X1 OAI21X1_2384 ( .gnd(gnd), .vdd(vdd), .A(_8338_), .B(_8339_), .C(_8340_), .Y(_8341_) );
NAND2X1 NAND2X1_1075 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_5_bF_buf2_), .B(micro_hash_ucr_2_pipe30_bF_buf1), .Y(_8342_) );
NAND3X1 NAND3X1_337 ( .gnd(gnd), .vdd(vdd), .A(_5112__bF_buf2), .B(_8342_), .C(_8341_), .Y(_8343_) );
NAND3X1 NAND3X1_338 ( .gnd(gnd), .vdd(vdd), .A(_5111__bF_buf0), .B(_8306_), .C(_8343_), .Y(_8344_) );
NAND3X1 NAND3X1_339 ( .gnd(gnd), .vdd(vdd), .A(_5107_), .B(_8305_), .C(_8344_), .Y(_8345_) );
NAND3X1 NAND3X1_340 ( .gnd(gnd), .vdd(vdd), .A(_5109__bF_buf2), .B(_8304_), .C(_8345_), .Y(_8346_) );
NAND3X1 NAND3X1_341 ( .gnd(gnd), .vdd(vdd), .A(_5108__bF_buf0), .B(_8303_), .C(_8346_), .Y(_8347_) );
NAND3X1 NAND3X1_342 ( .gnd(gnd), .vdd(vdd), .A(_5104__bF_buf0), .B(_8302_), .C(_8347_), .Y(_8348_) );
AOI21X1 AOI21X1_1474 ( .gnd(gnd), .vdd(vdd), .A(_8301_), .B(_8348_), .C(micro_hash_ucr_2_pipe37), .Y(_8349_) );
OAI21X1 OAI21X1_2385 ( .gnd(gnd), .vdd(vdd), .A(_5255_), .B(_5106_), .C(_5105__bF_buf4), .Y(_8350_) );
AOI21X1 AOI21X1_1475 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe38_bF_buf0), .B(_4608__bF_buf2), .C(micro_hash_ucr_2_pipe39), .Y(_8351_) );
OAI21X1 OAI21X1_2386 ( .gnd(gnd), .vdd(vdd), .A(_8349_), .B(_8350_), .C(_8351_), .Y(_8352_) );
AOI21X1 AOI21X1_1476 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_1_bF_buf2_), .B(micro_hash_ucr_2_pipe39), .C(micro_hash_ucr_2_pipe40_bF_buf2), .Y(_8353_) );
AOI22X1 AOI22X1_62 ( .gnd(gnd), .vdd(vdd), .A(_4608__bF_buf1), .B(micro_hash_ucr_2_pipe40_bF_buf1), .C(_8352_), .D(_8353_), .Y(_8354_) );
OAI21X1 OAI21X1_2387 ( .gnd(gnd), .vdd(vdd), .A(_5255_), .B(_5102_), .C(_5098__bF_buf0), .Y(_8355_) );
AOI21X1 AOI21X1_1477 ( .gnd(gnd), .vdd(vdd), .A(_5102_), .B(_8354_), .C(_8355_), .Y(_8356_) );
OAI21X1 OAI21X1_2388 ( .gnd(gnd), .vdd(vdd), .A(_5098__bF_buf4), .B(micro_hash_ucr_2_b_5_bF_buf1_), .C(_5100__bF_buf2), .Y(_8357_) );
OAI21X1 OAI21X1_2389 ( .gnd(gnd), .vdd(vdd), .A(_8356_), .B(_8357_), .C(_8300_), .Y(_8358_) );
OAI21X1 OAI21X1_2390 ( .gnd(gnd), .vdd(vdd), .A(_4608__bF_buf0), .B(_5099__bF_buf1), .C(_5095_), .Y(_8359_) );
AOI21X1 AOI21X1_1478 ( .gnd(gnd), .vdd(vdd), .A(_5099__bF_buf0), .B(_8358_), .C(_8359_), .Y(_8360_) );
OAI21X1 OAI21X1_2391 ( .gnd(gnd), .vdd(vdd), .A(_5095_), .B(micro_hash_ucr_2_c_1_bF_buf1_), .C(_5097__bF_buf1), .Y(_8361_) );
NAND2X1 NAND2X1_1076 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_5_bF_buf0_), .B(micro_hash_ucr_2_pipe46_bF_buf3), .Y(_8362_) );
OAI21X1 OAI21X1_2392 ( .gnd(gnd), .vdd(vdd), .A(_8360_), .B(_8361_), .C(_8362_), .Y(_8363_) );
OAI21X1 OAI21X1_2393 ( .gnd(gnd), .vdd(vdd), .A(_5255_), .B(_5096__bF_buf2), .C(_5092__bF_buf2), .Y(_8364_) );
AOI21X1 AOI21X1_1479 ( .gnd(gnd), .vdd(vdd), .A(_5096__bF_buf1), .B(_8363_), .C(_8364_), .Y(_8365_) );
OAI21X1 OAI21X1_2394 ( .gnd(gnd), .vdd(vdd), .A(_5092__bF_buf1), .B(micro_hash_ucr_2_b_5_bF_buf3_), .C(_5094_), .Y(_8366_) );
AOI21X1 AOI21X1_1480 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_1_bF_buf0_), .B(micro_hash_ucr_2_pipe49_bF_buf3), .C(micro_hash_ucr_2_pipe50_bF_buf0), .Y(_8367_) );
OAI21X1 OAI21X1_2395 ( .gnd(gnd), .vdd(vdd), .A(_8365_), .B(_8366_), .C(_8367_), .Y(_8368_) );
NAND2X1 NAND2X1_1077 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe50_bF_buf3), .B(_4608__bF_buf3), .Y(_8369_) );
NAND3X1 NAND3X1_343 ( .gnd(gnd), .vdd(vdd), .A(_5089__bF_buf2), .B(_8369_), .C(_8368_), .Y(_8370_) );
NAND3X1 NAND3X1_344 ( .gnd(gnd), .vdd(vdd), .A(_5091__bF_buf2), .B(_8299_), .C(_8370_), .Y(_8371_) );
NAND3X1 NAND3X1_345 ( .gnd(gnd), .vdd(vdd), .A(_5090_), .B(_8298_), .C(_8371_), .Y(_8372_) );
NAND3X1 NAND3X1_346 ( .gnd(gnd), .vdd(vdd), .A(_5086__bF_buf0), .B(_8297_), .C(_8372_), .Y(_8373_) );
NAND3X1 NAND3X1_347 ( .gnd(gnd), .vdd(vdd), .A(_5088_), .B(_8296_), .C(_8373_), .Y(_8374_) );
NAND3X1 NAND3X1_348 ( .gnd(gnd), .vdd(vdd), .A(_5087__bF_buf1), .B(_8295_), .C(_8374_), .Y(_8375_) );
NAND3X1 NAND3X1_349 ( .gnd(gnd), .vdd(vdd), .A(_5083_), .B(_8294_), .C(_8375_), .Y(_8376_) );
NAND3X1 NAND3X1_350 ( .gnd(gnd), .vdd(vdd), .A(_5085__bF_buf1), .B(_8293_), .C(_8376_), .Y(_8377_) );
NAND3X1 NAND3X1_351 ( .gnd(gnd), .vdd(vdd), .A(_5084__bF_buf3), .B(_8292_), .C(_8377_), .Y(_8378_) );
NAND3X1 NAND3X1_352 ( .gnd(gnd), .vdd(vdd), .A(_5080__bF_buf3), .B(_8291_), .C(_8378_), .Y(_8379_) );
NAND3X1 NAND3X1_353 ( .gnd(gnd), .vdd(vdd), .A(_5082_), .B(_8290_), .C(_8379_), .Y(_8380_) );
NAND3X1 NAND3X1_354 ( .gnd(gnd), .vdd(vdd), .A(_5081__bF_buf3), .B(_8289_), .C(_8380_), .Y(_8381_) );
NAND3X1 NAND3X1_355 ( .gnd(gnd), .vdd(vdd), .A(_5077__bF_buf1), .B(_8288_), .C(_8381_), .Y(_8382_) );
NAND3X1 NAND3X1_356 ( .gnd(gnd), .vdd(vdd), .A(_5079__bF_buf2), .B(_8287_), .C(_8382_), .Y(_8383_) );
NAND3X1 NAND3X1_357 ( .gnd(gnd), .vdd(vdd), .A(_5078_), .B(_8286_), .C(_8383_), .Y(_8384_) );
AOI21X1 AOI21X1_1481 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_1_bF_buf3_), .B(micro_hash_ucr_2_pipe65_bF_buf1), .C(micro_hash_ucr_2_pipe66_bF_buf1), .Y(_8385_) );
NAND2X1 NAND2X1_1078 ( .gnd(gnd), .vdd(vdd), .A(_8385_), .B(_8384_), .Y(_8386_) );
AOI21X1 AOI21X1_1482 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe66_bF_buf0), .B(_4608__bF_buf2), .C(micro_hash_ucr_2_pipe67), .Y(_8387_) );
OAI21X1 OAI21X1_2396 ( .gnd(gnd), .vdd(vdd), .A(_5255_), .B(_5076__bF_buf3), .C(_5075__bF_buf0), .Y(_8388_) );
AOI21X1 AOI21X1_1483 ( .gnd(gnd), .vdd(vdd), .A(_8387_), .B(_8386_), .C(_8388_), .Y(_8389_) );
OAI21X1 OAI21X1_2397 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_5_bF_buf2_), .B(_5075__bF_buf4), .C(_6146_), .Y(_8390_) );
OAI21X1 OAI21X1_2398 ( .gnd(gnd), .vdd(vdd), .A(_8389_), .B(_8390_), .C(_8285_), .Y(_4492__5_) );
NAND2X1 NAND2X1_1079 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe64_bF_buf1), .B(_4622__bF_buf1), .Y(_8391_) );
NAND2X1 NAND2X1_1080 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_2_bF_buf3_), .B(micro_hash_ucr_2_pipe63), .Y(_8392_) );
NAND2X1 NAND2X1_1081 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe62_bF_buf4), .B(_4622__bF_buf0), .Y(_8393_) );
NAND2X1 NAND2X1_1082 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_2_bF_buf2_), .B(micro_hash_ucr_2_pipe61_bF_buf1), .Y(_8394_) );
NAND2X1 NAND2X1_1083 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe60_bF_buf4), .B(_4622__bF_buf3), .Y(_8395_) );
NAND2X1 NAND2X1_1084 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_2_bF_buf1_), .B(micro_hash_ucr_2_pipe59), .Y(_8396_) );
NAND2X1 NAND2X1_1085 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe58_bF_buf2), .B(_4622__bF_buf2), .Y(_8397_) );
NAND2X1 NAND2X1_1086 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_2_bF_buf0_), .B(micro_hash_ucr_2_pipe57_bF_buf2), .Y(_8398_) );
NAND2X1 NAND2X1_1087 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe56_bF_buf1), .B(_4622__bF_buf1), .Y(_8399_) );
NAND2X1 NAND2X1_1088 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_2_bF_buf3_), .B(micro_hash_ucr_2_pipe55), .Y(_8400_) );
NAND2X1 NAND2X1_1089 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe54_bF_buf3), .B(_4622__bF_buf0), .Y(_8401_) );
NAND2X1 NAND2X1_1090 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_2_bF_buf2_), .B(micro_hash_ucr_2_pipe53_bF_buf3), .Y(_8402_) );
NAND2X1 NAND2X1_1091 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe52_bF_buf0), .B(_4622__bF_buf3), .Y(_8403_) );
NAND2X1 NAND2X1_1092 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_2_bF_buf1_), .B(micro_hash_ucr_2_pipe51), .Y(_8404_) );
NAND2X1 NAND2X1_1093 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_6_), .B(micro_hash_ucr_2_pipe46_bF_buf2), .Y(_8405_) );
NAND2X1 NAND2X1_1094 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_6_), .B(micro_hash_ucr_2_pipe44_bF_buf0), .Y(_8406_) );
NAND2X1 NAND2X1_1095 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_6_), .B(micro_hash_ucr_2_pipe38_bF_buf3), .Y(_8407_) );
NAND2X1 NAND2X1_1096 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe37), .B(_5372_), .Y(_8408_) );
NAND2X1 NAND2X1_1097 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_2_bF_buf0_), .B(micro_hash_ucr_2_pipe33_bF_buf2), .Y(_8409_) );
NAND2X1 NAND2X1_1098 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe29_bF_buf3), .B(_5372_), .Y(_8410_) );
NAND2X1 NAND2X1_1099 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_6_), .B(micro_hash_ucr_2_pipe28_bF_buf1), .Y(_8411_) );
NAND2X1 NAND2X1_1100 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe27), .B(_5372_), .Y(_8412_) );
NAND2X1 NAND2X1_1101 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_6_), .B(micro_hash_ucr_2_pipe26_bF_buf0), .Y(_8413_) );
NAND2X1 NAND2X1_1102 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe25), .B(_5372_), .Y(_8414_) );
NAND2X1 NAND2X1_1103 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_2_bF_buf3_), .B(micro_hash_ucr_2_pipe21_bF_buf0), .Y(_8415_) );
NAND2X1 NAND2X1_1104 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe20_bF_buf3), .B(_4622__bF_buf2), .Y(_8416_) );
NAND2X1 NAND2X1_1105 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_2_bF_buf2_), .B(micro_hash_ucr_2_pipe19), .Y(_8417_) );
NAND2X1 NAND2X1_1106 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe18_bF_buf1), .B(_4622__bF_buf1), .Y(_8418_) );
NAND2X1 NAND2X1_1107 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_2_bF_buf1_), .B(micro_hash_ucr_2_pipe17_bF_buf1), .Y(_8419_) );
NAND2X1 NAND2X1_1108 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe16_bF_buf0), .B(_4622__bF_buf0), .Y(_8420_) );
NAND2X1 NAND2X1_1109 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_2_bF_buf0_), .B(micro_hash_ucr_2_pipe15), .Y(_8421_) );
NAND2X1 NAND2X1_1110 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_2_bF_buf3_), .B(_5268_), .Y(_8422_) );
NAND3X1 NAND3X1_358 ( .gnd(gnd), .vdd(vdd), .A(H_2_14_), .B(_5132_), .C(_8311_), .Y(_8423_) );
OR2X2 OR2X2_64 ( .gnd(gnd), .vdd(vdd), .A(_8310_), .B(_8423_), .Y(_8424_) );
AOI21X1 AOI21X1_1484 ( .gnd(gnd), .vdd(vdd), .A(_8422_), .B(_8424_), .C(micro_hash_ucr_2_pipe12_bF_buf2), .Y(_8425_) );
OAI21X1 OAI21X1_2399 ( .gnd(gnd), .vdd(vdd), .A(_5385_), .B(_4622__bF_buf3), .C(_8208_), .Y(_8426_) );
NOR2X1 NOR2X1_1338 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe14_bF_buf4), .B(_5130_), .Y(_8427_) );
OAI21X1 OAI21X1_2400 ( .gnd(gnd), .vdd(vdd), .A(_5129_), .B(micro_hash_ucr_2_b_6_), .C(_5125__bF_buf3), .Y(_8428_) );
AOI21X1 AOI21X1_1485 ( .gnd(gnd), .vdd(vdd), .A(_5372_), .B(_8427_), .C(_8428_), .Y(_8429_) );
OAI21X1 OAI21X1_2401 ( .gnd(gnd), .vdd(vdd), .A(_8426_), .B(_8425_), .C(_8429_), .Y(_8430_) );
NAND3X1 NAND3X1_359 ( .gnd(gnd), .vdd(vdd), .A(_5127__bF_buf1), .B(_8421_), .C(_8430_), .Y(_8431_) );
NAND3X1 NAND3X1_360 ( .gnd(gnd), .vdd(vdd), .A(_5126_), .B(_8420_), .C(_8431_), .Y(_8432_) );
NAND3X1 NAND3X1_361 ( .gnd(gnd), .vdd(vdd), .A(_5122__bF_buf0), .B(_8419_), .C(_8432_), .Y(_8433_) );
NAND3X1 NAND3X1_362 ( .gnd(gnd), .vdd(vdd), .A(_5124__bF_buf0), .B(_8418_), .C(_8433_), .Y(_8434_) );
NAND3X1 NAND3X1_363 ( .gnd(gnd), .vdd(vdd), .A(_5123__bF_buf2), .B(_8417_), .C(_8434_), .Y(_8435_) );
NAND3X1 NAND3X1_364 ( .gnd(gnd), .vdd(vdd), .A(_5119_), .B(_8416_), .C(_8435_), .Y(_8436_) );
AOI21X1 AOI21X1_1486 ( .gnd(gnd), .vdd(vdd), .A(_8415_), .B(_8436_), .C(micro_hash_ucr_2_pipe22_bF_buf1), .Y(_8437_) );
OAI21X1 OAI21X1_2402 ( .gnd(gnd), .vdd(vdd), .A(_4622__bF_buf2), .B(_5121__bF_buf0), .C(_5120__bF_buf0), .Y(_8438_) );
AOI21X1 AOI21X1_1487 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe23), .B(_5372_), .C(micro_hash_ucr_2_pipe24_bF_buf2), .Y(_8439_) );
OAI21X1 OAI21X1_2403 ( .gnd(gnd), .vdd(vdd), .A(_8437_), .B(_8438_), .C(_8439_), .Y(_8440_) );
NAND2X1 NAND2X1_1111 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_6_), .B(micro_hash_ucr_2_pipe24_bF_buf1), .Y(_8441_) );
NAND3X1 NAND3X1_365 ( .gnd(gnd), .vdd(vdd), .A(_5118__bF_buf0), .B(_8441_), .C(_8440_), .Y(_8442_) );
NAND3X1 NAND3X1_366 ( .gnd(gnd), .vdd(vdd), .A(_5117__bF_buf1), .B(_8414_), .C(_8442_), .Y(_8443_) );
NAND3X1 NAND3X1_367 ( .gnd(gnd), .vdd(vdd), .A(_5113_), .B(_8413_), .C(_8443_), .Y(_8444_) );
NAND3X1 NAND3X1_368 ( .gnd(gnd), .vdd(vdd), .A(_5115__bF_buf0), .B(_8412_), .C(_8444_), .Y(_8445_) );
NAND3X1 NAND3X1_369 ( .gnd(gnd), .vdd(vdd), .A(_5114_), .B(_8411_), .C(_8445_), .Y(_8446_) );
NAND3X1 NAND3X1_370 ( .gnd(gnd), .vdd(vdd), .A(_5110__bF_buf1), .B(_8410_), .C(_8446_), .Y(_8447_) );
AOI21X1 AOI21X1_1488 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_6_), .B(micro_hash_ucr_2_pipe30_bF_buf0), .C(micro_hash_ucr_2_pipe31), .Y(_8448_) );
OAI21X1 OAI21X1_2404 ( .gnd(gnd), .vdd(vdd), .A(_5112__bF_buf1), .B(micro_hash_ucr_2_c_2_bF_buf2_), .C(_5111__bF_buf4), .Y(_8449_) );
AOI21X1 AOI21X1_1489 ( .gnd(gnd), .vdd(vdd), .A(_8448_), .B(_8447_), .C(_8449_), .Y(_8450_) );
NOR2X1 NOR2X1_1339 ( .gnd(gnd), .vdd(vdd), .A(_4622__bF_buf1), .B(_5111__bF_buf3), .Y(_8451_) );
OAI21X1 OAI21X1_2405 ( .gnd(gnd), .vdd(vdd), .A(_8450_), .B(_8451_), .C(_5107_), .Y(_8452_) );
AOI21X1 AOI21X1_1490 ( .gnd(gnd), .vdd(vdd), .A(_8409_), .B(_8452_), .C(micro_hash_ucr_2_pipe34_bF_buf1), .Y(_8453_) );
OAI21X1 OAI21X1_2406 ( .gnd(gnd), .vdd(vdd), .A(_4622__bF_buf0), .B(_5109__bF_buf1), .C(_5108__bF_buf3), .Y(_8454_) );
AOI21X1 AOI21X1_1491 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe35), .B(_5372_), .C(micro_hash_ucr_2_pipe36_bF_buf2), .Y(_8455_) );
OAI21X1 OAI21X1_2407 ( .gnd(gnd), .vdd(vdd), .A(_8453_), .B(_8454_), .C(_8455_), .Y(_8456_) );
NAND2X1 NAND2X1_1112 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_6_), .B(micro_hash_ucr_2_pipe36_bF_buf1), .Y(_8457_) );
NAND3X1 NAND3X1_371 ( .gnd(gnd), .vdd(vdd), .A(_5106_), .B(_8457_), .C(_8456_), .Y(_8458_) );
NAND3X1 NAND3X1_372 ( .gnd(gnd), .vdd(vdd), .A(_5105__bF_buf3), .B(_8408_), .C(_8458_), .Y(_8459_) );
AOI21X1 AOI21X1_1492 ( .gnd(gnd), .vdd(vdd), .A(_8407_), .B(_8459_), .C(micro_hash_ucr_2_pipe39), .Y(_8460_) );
OAI21X1 OAI21X1_2408 ( .gnd(gnd), .vdd(vdd), .A(_5372_), .B(_5101_), .C(_5103__bF_buf2), .Y(_8461_) );
AOI21X1 AOI21X1_1493 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe40_bF_buf0), .B(_4622__bF_buf3), .C(micro_hash_ucr_2_pipe41_bF_buf1), .Y(_8462_) );
OAI21X1 OAI21X1_2409 ( .gnd(gnd), .vdd(vdd), .A(_8460_), .B(_8461_), .C(_8462_), .Y(_8463_) );
AOI21X1 AOI21X1_1494 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_2_bF_buf1_), .B(micro_hash_ucr_2_pipe41_bF_buf0), .C(micro_hash_ucr_2_pipe42_bF_buf3), .Y(_8464_) );
AOI22X1 AOI22X1_63 ( .gnd(gnd), .vdd(vdd), .A(_4622__bF_buf2), .B(micro_hash_ucr_2_pipe42_bF_buf2), .C(_8463_), .D(_8464_), .Y(_8465_) );
NAND2X1 NAND2X1_1113 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe43), .B(_5372_), .Y(_8466_) );
OAI21X1 OAI21X1_2410 ( .gnd(gnd), .vdd(vdd), .A(_8465_), .B(micro_hash_ucr_2_pipe43), .C(_8466_), .Y(_8467_) );
OAI21X1 OAI21X1_2411 ( .gnd(gnd), .vdd(vdd), .A(_8467_), .B(micro_hash_ucr_2_pipe44_bF_buf3), .C(_8406_), .Y(_8468_) );
NAND2X1 NAND2X1_1114 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe45_bF_buf3), .B(_5372_), .Y(_8469_) );
OAI21X1 OAI21X1_2412 ( .gnd(gnd), .vdd(vdd), .A(_8468_), .B(micro_hash_ucr_2_pipe45_bF_buf2), .C(_8469_), .Y(_8470_) );
OAI21X1 OAI21X1_2413 ( .gnd(gnd), .vdd(vdd), .A(_8470_), .B(micro_hash_ucr_2_pipe46_bF_buf1), .C(_8405_), .Y(_8471_) );
NAND2X1 NAND2X1_1115 ( .gnd(gnd), .vdd(vdd), .A(_5096__bF_buf0), .B(_8471_), .Y(_8472_) );
OAI21X1 OAI21X1_2414 ( .gnd(gnd), .vdd(vdd), .A(_5372_), .B(_5096__bF_buf3), .C(_8472_), .Y(_8473_) );
AOI21X1 AOI21X1_1495 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe48_bF_buf2), .B(_4622__bF_buf1), .C(micro_hash_ucr_2_pipe49_bF_buf2), .Y(_8474_) );
OAI21X1 OAI21X1_2415 ( .gnd(gnd), .vdd(vdd), .A(_8473_), .B(micro_hash_ucr_2_pipe48_bF_buf1), .C(_8474_), .Y(_8475_) );
AOI21X1 AOI21X1_1496 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_2_bF_buf0_), .B(micro_hash_ucr_2_pipe49_bF_buf1), .C(micro_hash_ucr_2_pipe50_bF_buf2), .Y(_8476_) );
NAND2X1 NAND2X1_1116 ( .gnd(gnd), .vdd(vdd), .A(_8476_), .B(_8475_), .Y(_8477_) );
NAND2X1 NAND2X1_1117 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe50_bF_buf1), .B(_4622__bF_buf0), .Y(_8478_) );
NAND3X1 NAND3X1_373 ( .gnd(gnd), .vdd(vdd), .A(_5089__bF_buf1), .B(_8478_), .C(_8477_), .Y(_8479_) );
NAND3X1 NAND3X1_374 ( .gnd(gnd), .vdd(vdd), .A(_5091__bF_buf1), .B(_8404_), .C(_8479_), .Y(_8480_) );
NAND3X1 NAND3X1_375 ( .gnd(gnd), .vdd(vdd), .A(_5090_), .B(_8403_), .C(_8480_), .Y(_8481_) );
NAND3X1 NAND3X1_376 ( .gnd(gnd), .vdd(vdd), .A(_5086__bF_buf3), .B(_8402_), .C(_8481_), .Y(_8482_) );
NAND3X1 NAND3X1_377 ( .gnd(gnd), .vdd(vdd), .A(_5088_), .B(_8401_), .C(_8482_), .Y(_8483_) );
NAND3X1 NAND3X1_378 ( .gnd(gnd), .vdd(vdd), .A(_5087__bF_buf0), .B(_8400_), .C(_8483_), .Y(_8484_) );
NAND3X1 NAND3X1_379 ( .gnd(gnd), .vdd(vdd), .A(_5083_), .B(_8399_), .C(_8484_), .Y(_8485_) );
NAND3X1 NAND3X1_380 ( .gnd(gnd), .vdd(vdd), .A(_5085__bF_buf0), .B(_8398_), .C(_8485_), .Y(_8486_) );
NAND3X1 NAND3X1_381 ( .gnd(gnd), .vdd(vdd), .A(_5084__bF_buf2), .B(_8397_), .C(_8486_), .Y(_8487_) );
NAND3X1 NAND3X1_382 ( .gnd(gnd), .vdd(vdd), .A(_5080__bF_buf2), .B(_8396_), .C(_8487_), .Y(_8488_) );
NAND3X1 NAND3X1_383 ( .gnd(gnd), .vdd(vdd), .A(_5082_), .B(_8395_), .C(_8488_), .Y(_8489_) );
NAND3X1 NAND3X1_384 ( .gnd(gnd), .vdd(vdd), .A(_5081__bF_buf2), .B(_8394_), .C(_8489_), .Y(_8490_) );
NAND3X1 NAND3X1_385 ( .gnd(gnd), .vdd(vdd), .A(_5077__bF_buf0), .B(_8393_), .C(_8490_), .Y(_8491_) );
NAND3X1 NAND3X1_386 ( .gnd(gnd), .vdd(vdd), .A(_5079__bF_buf1), .B(_8392_), .C(_8491_), .Y(_8492_) );
NAND3X1 NAND3X1_387 ( .gnd(gnd), .vdd(vdd), .A(_5078_), .B(_8391_), .C(_8492_), .Y(_8493_) );
AOI21X1 AOI21X1_1497 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_2_bF_buf3_), .B(micro_hash_ucr_2_pipe65_bF_buf0), .C(micro_hash_ucr_2_pipe66_bF_buf4), .Y(_8494_) );
NAND2X1 NAND2X1_1118 ( .gnd(gnd), .vdd(vdd), .A(_8494_), .B(_8493_), .Y(_8495_) );
AOI21X1 AOI21X1_1498 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe66_bF_buf3), .B(_4622__bF_buf3), .C(micro_hash_ucr_2_pipe67), .Y(_8496_) );
OAI21X1 OAI21X1_2416 ( .gnd(gnd), .vdd(vdd), .A(_5372_), .B(_5076__bF_buf2), .C(_5075__bF_buf3), .Y(_8497_) );
AOI21X1 AOI21X1_1499 ( .gnd(gnd), .vdd(vdd), .A(_8496_), .B(_8495_), .C(_8497_), .Y(_8498_) );
OAI21X1 OAI21X1_2417 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_6_), .B(_5075__bF_buf2), .C(_6146_), .Y(_8499_) );
OAI22X1 OAI22X1_110 ( .gnd(gnd), .vdd(vdd), .A(_5372_), .B(_7300_), .C(_8498_), .D(_8499_), .Y(_4492__6_) );
NAND2X1 NAND2X1_1119 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_3_bF_buf0_), .B(_4563_), .Y(_8500_) );
NAND2X1 NAND2X1_1120 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_7_bF_buf2_), .B(micro_hash_ucr_2_pipe66_bF_buf2), .Y(_8501_) );
NAND2X1 NAND2X1_1121 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe65_bF_buf3), .B(_8654_), .Y(_8502_) );
NAND2X1 NAND2X1_1122 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_7_bF_buf1_), .B(micro_hash_ucr_2_pipe64_bF_buf0), .Y(_8503_) );
NAND2X1 NAND2X1_1123 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe63), .B(_8654_), .Y(_8504_) );
NAND2X1 NAND2X1_1124 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_7_bF_buf0_), .B(micro_hash_ucr_2_pipe62_bF_buf3), .Y(_8505_) );
NAND2X1 NAND2X1_1125 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe61_bF_buf0), .B(_8654_), .Y(_8506_) );
NAND2X1 NAND2X1_1126 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_3_bF_buf3_), .B(micro_hash_ucr_2_pipe57_bF_buf1), .Y(_8507_) );
NAND2X1 NAND2X1_1127 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe56_bF_buf0), .B(_6135__bF_buf2), .Y(_8508_) );
NAND2X1 NAND2X1_1128 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_3_bF_buf2_), .B(micro_hash_ucr_2_pipe55), .Y(_8509_) );
NAND2X1 NAND2X1_1129 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe54_bF_buf2), .B(_6135__bF_buf1), .Y(_8510_) );
NAND2X1 NAND2X1_1130 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_3_bF_buf1_), .B(micro_hash_ucr_2_pipe53_bF_buf2), .Y(_8511_) );
NAND2X1 NAND2X1_1131 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe43), .B(_8654_), .Y(_8512_) );
NAND2X1 NAND2X1_1132 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_7_bF_buf3_), .B(micro_hash_ucr_2_pipe42_bF_buf1), .Y(_8513_) );
NAND2X1 NAND2X1_1133 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe41_bF_buf3), .B(_8654_), .Y(_8514_) );
NAND2X1 NAND2X1_1134 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_3_bF_buf0_), .B(micro_hash_ucr_2_pipe39), .Y(_8515_) );
NAND2X1 NAND2X1_1135 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe34_bF_buf0), .B(_6135__bF_buf0), .Y(_8516_) );
NAND2X1 NAND2X1_1136 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_3_bF_buf3_), .B(micro_hash_ucr_2_pipe33_bF_buf1), .Y(_8517_) );
NAND2X1 NAND2X1_1137 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe29_bF_buf2), .B(_8654_), .Y(_8518_) );
NAND2X1 NAND2X1_1138 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_7_bF_buf2_), .B(micro_hash_ucr_2_pipe28_bF_buf0), .Y(_8519_) );
NAND2X1 NAND2X1_1139 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe27), .B(_8654_), .Y(_8520_) );
NAND2X1 NAND2X1_1140 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_3_bF_buf2_), .B(micro_hash_ucr_2_pipe23), .Y(_8521_) );
NAND2X1 NAND2X1_1141 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe22_bF_buf0), .B(_6135__bF_buf3), .Y(_8522_) );
NAND2X1 NAND2X1_1142 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_3_bF_buf1_), .B(micro_hash_ucr_2_pipe21_bF_buf3), .Y(_8523_) );
NAND2X1 NAND2X1_1143 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe20_bF_buf2), .B(_6135__bF_buf2), .Y(_8524_) );
NAND2X1 NAND2X1_1144 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_3_bF_buf0_), .B(micro_hash_ucr_2_pipe19), .Y(_8525_) );
NAND2X1 NAND2X1_1145 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe18_bF_buf0), .B(_6135__bF_buf1), .Y(_8526_) );
NAND2X1 NAND2X1_1146 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_3_bF_buf3_), .B(micro_hash_ucr_2_pipe17_bF_buf0), .Y(_8527_) );
NAND2X1 NAND2X1_1147 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe16_bF_buf4), .B(_6135__bF_buf0), .Y(_8528_) );
NAND2X1 NAND2X1_1148 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_3_bF_buf2_), .B(micro_hash_ucr_2_pipe15), .Y(_8529_) );
NAND2X1 NAND2X1_1149 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe14_bF_buf3), .B(_6135__bF_buf3), .Y(_8530_) );
NAND2X1 NAND2X1_1150 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_3_bF_buf1_), .B(micro_hash_ucr_2_pipe13), .Y(_8531_) );
NOR2X1 NOR2X1_1340 ( .gnd(gnd), .vdd(vdd), .A(H_2_15_), .B(micro_hash_ucr_2_pipe11), .Y(_8532_) );
NAND2X1 NAND2X1_1151 ( .gnd(gnd), .vdd(vdd), .A(_8311_), .B(_8532_), .Y(_8533_) );
NOR2X1 NOR2X1_1341 ( .gnd(gnd), .vdd(vdd), .A(_8533_), .B(_8310_), .Y(_8534_) );
AOI21X1 AOI21X1_1500 ( .gnd(gnd), .vdd(vdd), .A(_8654_), .B(_5268_), .C(_8534_), .Y(_8535_) );
AOI21X1 AOI21X1_1501 ( .gnd(gnd), .vdd(vdd), .A(_6135__bF_buf2), .B(_5160_), .C(micro_hash_ucr_2_pipe13), .Y(_8536_) );
OAI21X1 OAI21X1_2418 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe12_bF_buf1), .B(_8535_), .C(_8536_), .Y(_8537_) );
NAND3X1 NAND3X1_388 ( .gnd(gnd), .vdd(vdd), .A(_5129_), .B(_8531_), .C(_8537_), .Y(_8538_) );
NAND3X1 NAND3X1_389 ( .gnd(gnd), .vdd(vdd), .A(_5125__bF_buf2), .B(_8530_), .C(_8538_), .Y(_8539_) );
NAND3X1 NAND3X1_390 ( .gnd(gnd), .vdd(vdd), .A(_5127__bF_buf0), .B(_8529_), .C(_8539_), .Y(_8540_) );
NAND3X1 NAND3X1_391 ( .gnd(gnd), .vdd(vdd), .A(_5126_), .B(_8528_), .C(_8540_), .Y(_8541_) );
NAND3X1 NAND3X1_392 ( .gnd(gnd), .vdd(vdd), .A(_5122__bF_buf4), .B(_8527_), .C(_8541_), .Y(_8542_) );
NAND3X1 NAND3X1_393 ( .gnd(gnd), .vdd(vdd), .A(_5124__bF_buf3), .B(_8526_), .C(_8542_), .Y(_8543_) );
NAND3X1 NAND3X1_394 ( .gnd(gnd), .vdd(vdd), .A(_5123__bF_buf1), .B(_8525_), .C(_8543_), .Y(_8544_) );
NAND3X1 NAND3X1_395 ( .gnd(gnd), .vdd(vdd), .A(_5119_), .B(_8524_), .C(_8544_), .Y(_8545_) );
NAND3X1 NAND3X1_396 ( .gnd(gnd), .vdd(vdd), .A(_5121__bF_buf4), .B(_8523_), .C(_8545_), .Y(_8546_) );
NAND3X1 NAND3X1_397 ( .gnd(gnd), .vdd(vdd), .A(_5120__bF_buf3), .B(_8522_), .C(_8546_), .Y(_8547_) );
AOI21X1 AOI21X1_1502 ( .gnd(gnd), .vdd(vdd), .A(_8521_), .B(_8547_), .C(micro_hash_ucr_2_pipe24_bF_buf0), .Y(_8548_) );
OAI21X1 OAI21X1_2419 ( .gnd(gnd), .vdd(vdd), .A(_6135__bF_buf1), .B(_5116__bF_buf3), .C(_5118__bF_buf3), .Y(_8549_) );
AOI21X1 AOI21X1_1503 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe25), .B(_8654_), .C(micro_hash_ucr_2_pipe26_bF_buf3), .Y(_8550_) );
OAI21X1 OAI21X1_2420 ( .gnd(gnd), .vdd(vdd), .A(_8548_), .B(_8549_), .C(_8550_), .Y(_8551_) );
NAND2X1 NAND2X1_1152 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_7_bF_buf1_), .B(micro_hash_ucr_2_pipe26_bF_buf2), .Y(_8552_) );
NAND3X1 NAND3X1_398 ( .gnd(gnd), .vdd(vdd), .A(_5113_), .B(_8552_), .C(_8551_), .Y(_8553_) );
NAND3X1 NAND3X1_399 ( .gnd(gnd), .vdd(vdd), .A(_5115__bF_buf4), .B(_8520_), .C(_8553_), .Y(_8554_) );
NAND3X1 NAND3X1_400 ( .gnd(gnd), .vdd(vdd), .A(_5114_), .B(_8519_), .C(_8554_), .Y(_8555_) );
NAND3X1 NAND3X1_401 ( .gnd(gnd), .vdd(vdd), .A(_5110__bF_buf0), .B(_8518_), .C(_8555_), .Y(_8556_) );
AOI21X1 AOI21X1_1504 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_7_bF_buf0_), .B(micro_hash_ucr_2_pipe30_bF_buf4), .C(micro_hash_ucr_2_pipe31), .Y(_8557_) );
OAI21X1 OAI21X1_2421 ( .gnd(gnd), .vdd(vdd), .A(_5112__bF_buf0), .B(micro_hash_ucr_2_c_3_bF_buf0_), .C(_5111__bF_buf2), .Y(_8558_) );
AOI21X1 AOI21X1_1505 ( .gnd(gnd), .vdd(vdd), .A(_8557_), .B(_8556_), .C(_8558_), .Y(_8559_) );
NOR2X1 NOR2X1_1342 ( .gnd(gnd), .vdd(vdd), .A(_6135__bF_buf0), .B(_5111__bF_buf1), .Y(_8560_) );
OAI21X1 OAI21X1_2422 ( .gnd(gnd), .vdd(vdd), .A(_8559_), .B(_8560_), .C(_5107_), .Y(_8561_) );
NAND3X1 NAND3X1_402 ( .gnd(gnd), .vdd(vdd), .A(_5109__bF_buf0), .B(_8517_), .C(_8561_), .Y(_8562_) );
NAND3X1 NAND3X1_403 ( .gnd(gnd), .vdd(vdd), .A(_5108__bF_buf2), .B(_8516_), .C(_8562_), .Y(_8563_) );
AOI21X1 AOI21X1_1506 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_3_bF_buf3_), .B(micro_hash_ucr_2_pipe35), .C(micro_hash_ucr_2_pipe36_bF_buf0), .Y(_8564_) );
OAI21X1 OAI21X1_2423 ( .gnd(gnd), .vdd(vdd), .A(_5104__bF_buf4), .B(micro_hash_ucr_2_b_7_bF_buf3_), .C(_5106_), .Y(_8565_) );
AOI21X1 AOI21X1_1507 ( .gnd(gnd), .vdd(vdd), .A(_8564_), .B(_8563_), .C(_8565_), .Y(_8566_) );
OAI21X1 OAI21X1_2424 ( .gnd(gnd), .vdd(vdd), .A(_8654_), .B(_5106_), .C(_5105__bF_buf2), .Y(_8567_) );
NAND2X1 NAND2X1_1153 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe38_bF_buf2), .B(_6135__bF_buf3), .Y(_8568_) );
OAI21X1 OAI21X1_2425 ( .gnd(gnd), .vdd(vdd), .A(_8566_), .B(_8567_), .C(_8568_), .Y(_8569_) );
OAI21X1 OAI21X1_2426 ( .gnd(gnd), .vdd(vdd), .A(_8569_), .B(micro_hash_ucr_2_pipe39), .C(_8515_), .Y(_8570_) );
NAND2X1 NAND2X1_1154 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe40_bF_buf4), .B(_6135__bF_buf2), .Y(_8571_) );
OAI21X1 OAI21X1_2427 ( .gnd(gnd), .vdd(vdd), .A(_8570_), .B(micro_hash_ucr_2_pipe40_bF_buf3), .C(_8571_), .Y(_8572_) );
NAND2X1 NAND2X1_1155 ( .gnd(gnd), .vdd(vdd), .A(_5102_), .B(_8572_), .Y(_8573_) );
NAND3X1 NAND3X1_404 ( .gnd(gnd), .vdd(vdd), .A(_5098__bF_buf3), .B(_8514_), .C(_8573_), .Y(_8574_) );
NAND3X1 NAND3X1_405 ( .gnd(gnd), .vdd(vdd), .A(_5100__bF_buf1), .B(_8513_), .C(_8574_), .Y(_8575_) );
NAND3X1 NAND3X1_406 ( .gnd(gnd), .vdd(vdd), .A(_5099__bF_buf4), .B(_8512_), .C(_8575_), .Y(_8576_) );
AOI21X1 AOI21X1_1508 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_7_bF_buf2_), .B(micro_hash_ucr_2_pipe44_bF_buf2), .C(micro_hash_ucr_2_pipe45_bF_buf1), .Y(_8577_) );
OAI21X1 OAI21X1_2428 ( .gnd(gnd), .vdd(vdd), .A(_5095_), .B(micro_hash_ucr_2_c_3_bF_buf2_), .C(_5097__bF_buf0), .Y(_8578_) );
AOI21X1 AOI21X1_1509 ( .gnd(gnd), .vdd(vdd), .A(_8577_), .B(_8576_), .C(_8578_), .Y(_8579_) );
NOR2X1 NOR2X1_1343 ( .gnd(gnd), .vdd(vdd), .A(_6135__bF_buf1), .B(_5097__bF_buf3), .Y(_8580_) );
OAI21X1 OAI21X1_2429 ( .gnd(gnd), .vdd(vdd), .A(_8579_), .B(_8580_), .C(_5096__bF_buf2), .Y(_8581_) );
AOI21X1 AOI21X1_1510 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_c_3_bF_buf1_), .B(micro_hash_ucr_2_pipe47), .C(micro_hash_ucr_2_pipe48_bF_buf0), .Y(_8582_) );
OAI21X1 OAI21X1_2430 ( .gnd(gnd), .vdd(vdd), .A(_5092__bF_buf0), .B(micro_hash_ucr_2_b_7_bF_buf1_), .C(_5094_), .Y(_8583_) );
AOI21X1 AOI21X1_1511 ( .gnd(gnd), .vdd(vdd), .A(_8582_), .B(_8581_), .C(_8583_), .Y(_8584_) );
OAI21X1 OAI21X1_2431 ( .gnd(gnd), .vdd(vdd), .A(_8654_), .B(_5094_), .C(_5093__bF_buf0), .Y(_8585_) );
OAI22X1 OAI22X1_111 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_7_bF_buf0_), .B(_5093__bF_buf4), .C(_8584_), .D(_8585_), .Y(_8586_) );
OAI21X1 OAI21X1_2432 ( .gnd(gnd), .vdd(vdd), .A(_5089__bF_buf0), .B(micro_hash_ucr_2_c_3_bF_buf0_), .C(_5091__bF_buf0), .Y(_8587_) );
AOI21X1 AOI21X1_1512 ( .gnd(gnd), .vdd(vdd), .A(_5089__bF_buf3), .B(_8586_), .C(_8587_), .Y(_8588_) );
NOR2X1 NOR2X1_1344 ( .gnd(gnd), .vdd(vdd), .A(_6135__bF_buf0), .B(_5091__bF_buf4), .Y(_8589_) );
OAI21X1 OAI21X1_2433 ( .gnd(gnd), .vdd(vdd), .A(_8588_), .B(_8589_), .C(_5090_), .Y(_8590_) );
NAND3X1 NAND3X1_407 ( .gnd(gnd), .vdd(vdd), .A(_5086__bF_buf2), .B(_8511_), .C(_8590_), .Y(_8591_) );
NAND3X1 NAND3X1_408 ( .gnd(gnd), .vdd(vdd), .A(_5088_), .B(_8510_), .C(_8591_), .Y(_8592_) );
NAND3X1 NAND3X1_409 ( .gnd(gnd), .vdd(vdd), .A(_5087__bF_buf4), .B(_8509_), .C(_8592_), .Y(_8593_) );
NAND3X1 NAND3X1_410 ( .gnd(gnd), .vdd(vdd), .A(_5083_), .B(_8508_), .C(_8593_), .Y(_8594_) );
AOI21X1 AOI21X1_1513 ( .gnd(gnd), .vdd(vdd), .A(_8507_), .B(_8594_), .C(micro_hash_ucr_2_pipe58_bF_buf1), .Y(_8595_) );
OAI21X1 OAI21X1_2434 ( .gnd(gnd), .vdd(vdd), .A(_6135__bF_buf3), .B(_5085__bF_buf3), .C(_5084__bF_buf1), .Y(_8596_) );
AOI21X1 AOI21X1_1514 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe59), .B(_8654_), .C(micro_hash_ucr_2_pipe60_bF_buf3), .Y(_8597_) );
OAI21X1 OAI21X1_2435 ( .gnd(gnd), .vdd(vdd), .A(_8595_), .B(_8596_), .C(_8597_), .Y(_8598_) );
NAND2X1 NAND2X1_1156 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_7_bF_buf3_), .B(micro_hash_ucr_2_pipe60_bF_buf2), .Y(_8599_) );
NAND3X1 NAND3X1_411 ( .gnd(gnd), .vdd(vdd), .A(_5082_), .B(_8599_), .C(_8598_), .Y(_8600_) );
NAND3X1 NAND3X1_412 ( .gnd(gnd), .vdd(vdd), .A(_5081__bF_buf1), .B(_8506_), .C(_8600_), .Y(_8601_) );
NAND3X1 NAND3X1_413 ( .gnd(gnd), .vdd(vdd), .A(_5077__bF_buf3), .B(_8505_), .C(_8601_), .Y(_8602_) );
NAND3X1 NAND3X1_414 ( .gnd(gnd), .vdd(vdd), .A(_5079__bF_buf0), .B(_8504_), .C(_8602_), .Y(_8603_) );
NAND3X1 NAND3X1_415 ( .gnd(gnd), .vdd(vdd), .A(_5078_), .B(_8503_), .C(_8603_), .Y(_8604_) );
NAND3X1 NAND3X1_416 ( .gnd(gnd), .vdd(vdd), .A(_5074__bF_buf2), .B(_8502_), .C(_8604_), .Y(_8605_) );
NAND2X1 NAND2X1_1157 ( .gnd(gnd), .vdd(vdd), .A(_8501_), .B(_8605_), .Y(_8606_) );
OAI21X1 OAI21X1_2436 ( .gnd(gnd), .vdd(vdd), .A(_8654_), .B(_5076__bF_buf1), .C(_5075__bF_buf1), .Y(_8607_) );
AOI21X1 AOI21X1_1515 ( .gnd(gnd), .vdd(vdd), .A(_5076__bF_buf0), .B(_8606_), .C(_8607_), .Y(_8608_) );
OAI21X1 OAI21X1_2437 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_b_7_bF_buf2_), .B(_5075__bF_buf0), .C(_6146_), .Y(_8609_) );
OAI21X1 OAI21X1_2438 ( .gnd(gnd), .vdd(vdd), .A(_8608_), .B(_8609_), .C(_8500_), .Y(_4492__7_) );
AOI21X1 AOI21X1_1516 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_136_), .B(_4782_), .C(micro_hash_ucr_2_Wx_224_), .Y(_8610_) );
OAI21X1 OAI21X1_2439 ( .gnd(gnd), .vdd(vdd), .A(_4782_), .B(micro_hash_ucr_2_Wx_136_), .C(_8610_), .Y(_8611_) );
AND2X2 AND2X2_507 ( .gnd(gnd), .vdd(vdd), .A(_8611_), .B(_4496__bF_buf5), .Y(_4490__248_) );
OAI21X1 OAI21X1_2440 ( .gnd(gnd), .vdd(vdd), .A(_4786_), .B(micro_hash_ucr_2_Wx_137_), .C(_6476_), .Y(_8612_) );
AOI21X1 AOI21X1_1517 ( .gnd(gnd), .vdd(vdd), .A(_4786_), .B(micro_hash_ucr_2_Wx_137_), .C(_8612_), .Y(_8613_) );
NOR2X1 NOR2X1_1345 ( .gnd(gnd), .vdd(vdd), .A(_8613_), .B(_4594__bF_buf10), .Y(_4490__249_) );
OAI21X1 OAI21X1_2441 ( .gnd(gnd), .vdd(vdd), .A(_4790_), .B(micro_hash_ucr_2_Wx_138_), .C(_6504_), .Y(_8614_) );
AOI21X1 AOI21X1_1518 ( .gnd(gnd), .vdd(vdd), .A(_4790_), .B(micro_hash_ucr_2_Wx_138_), .C(_8614_), .Y(_8615_) );
NOR2X1 NOR2X1_1346 ( .gnd(gnd), .vdd(vdd), .A(_8615_), .B(_4594__bF_buf9), .Y(_4490__250_) );
OAI21X1 OAI21X1_2442 ( .gnd(gnd), .vdd(vdd), .A(_4794_), .B(micro_hash_ucr_2_Wx_139_), .C(_7023_), .Y(_8616_) );
AOI21X1 AOI21X1_1519 ( .gnd(gnd), .vdd(vdd), .A(_4794_), .B(micro_hash_ucr_2_Wx_139_), .C(_8616_), .Y(_8617_) );
NOR2X1 NOR2X1_1347 ( .gnd(gnd), .vdd(vdd), .A(_8617_), .B(_4594__bF_buf8), .Y(_4490__251_) );
AOI21X1 AOI21X1_1520 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_140_), .B(_4798_), .C(micro_hash_ucr_2_Wx_228_), .Y(_8618_) );
OAI21X1 OAI21X1_2443 ( .gnd(gnd), .vdd(vdd), .A(_4798_), .B(micro_hash_ucr_2_Wx_140_), .C(_8618_), .Y(_8619_) );
AND2X2 AND2X2_508 ( .gnd(gnd), .vdd(vdd), .A(_8619_), .B(_4496__bF_buf4), .Y(_4490__252_) );
AOI21X1 AOI21X1_1521 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_141_), .B(_4802_), .C(micro_hash_ucr_2_Wx_229_), .Y(_8620_) );
OAI21X1 OAI21X1_2444 ( .gnd(gnd), .vdd(vdd), .A(_4802_), .B(micro_hash_ucr_2_Wx_141_), .C(_8620_), .Y(_8621_) );
AND2X2 AND2X2_509 ( .gnd(gnd), .vdd(vdd), .A(_8621_), .B(_4496__bF_buf3), .Y(_4490__253_) );
OAI21X1 OAI21X1_2445 ( .gnd(gnd), .vdd(vdd), .A(_4806_), .B(micro_hash_ucr_2_Wx_142_), .C(_7746_), .Y(_8622_) );
AOI21X1 AOI21X1_1522 ( .gnd(gnd), .vdd(vdd), .A(_4806_), .B(micro_hash_ucr_2_Wx_142_), .C(_8622_), .Y(_8623_) );
NOR2X1 NOR2X1_1348 ( .gnd(gnd), .vdd(vdd), .A(_8623_), .B(_4594__bF_buf7), .Y(_4490__254_) );
AOI21X1 AOI21X1_1523 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_Wx_143_), .B(_4809_), .C(micro_hash_ucr_2_Wx_231_), .Y(_8624_) );
OAI21X1 OAI21X1_2446 ( .gnd(gnd), .vdd(vdd), .A(_4809_), .B(micro_hash_ucr_2_Wx_143_), .C(_8624_), .Y(_8625_) );
AND2X2 AND2X2_510 ( .gnd(gnd), .vdd(vdd), .A(_8625_), .B(_4496__bF_buf2), .Y(_4490__255_) );
OAI21X1 OAI21X1_2447 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe70_bF_buf1), .B(comparador_2_valid_hash), .C(_4496__bF_buf1), .Y(_8626_) );
NOR2X1 NOR2X1_1349 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_2_pipe71), .B(_8626_), .Y(_4568_) );
DFFPOSX1 DFFPOSX1_784 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_4494__0_), .Q(H_2_0_) );
DFFPOSX1 DFFPOSX1_785 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_4494__1_), .Q(H_2_1_) );
DFFPOSX1 DFFPOSX1_786 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_4494__2_), .Q(H_2_2_) );
DFFPOSX1 DFFPOSX1_787 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_4494__3_), .Q(H_2_3_) );
DFFPOSX1 DFFPOSX1_788 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_4494__4_), .Q(H_2_4_) );
DFFPOSX1 DFFPOSX1_789 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_4494__5_), .Q(H_2_5_) );
DFFPOSX1 DFFPOSX1_790 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_4494__6_), .Q(H_2_6_) );
DFFPOSX1 DFFPOSX1_791 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf157), .D(_4494__7_), .Q(H_2_7_) );
DFFPOSX1 DFFPOSX1_792 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf156), .D(_4494__8_), .Q(H_2_8_) );
DFFPOSX1 DFFPOSX1_793 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf155), .D(_4494__9_), .Q(H_2_9_) );
DFFPOSX1 DFFPOSX1_794 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf154), .D(_4494__10_), .Q(H_2_10_) );
DFFPOSX1 DFFPOSX1_795 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf153), .D(_4494__11_), .Q(H_2_11_) );
DFFPOSX1 DFFPOSX1_796 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf152), .D(_4494__12_), .Q(H_2_12_) );
DFFPOSX1 DFFPOSX1_797 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf151), .D(_4494__13_), .Q(H_2_13_) );
DFFPOSX1 DFFPOSX1_798 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf150), .D(_4494__14_), .Q(H_2_14_) );
DFFPOSX1 DFFPOSX1_799 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf149), .D(_4494__15_), .Q(H_2_15_) );
DFFPOSX1 DFFPOSX1_800 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf148), .D(_4494__16_), .Q(H_2_16_) );
DFFPOSX1 DFFPOSX1_801 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf147), .D(_4494__17_), .Q(H_2_17_) );
DFFPOSX1 DFFPOSX1_802 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf146), .D(_4494__18_), .Q(H_2_18_) );
DFFPOSX1 DFFPOSX1_803 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf145), .D(_4494__19_), .Q(H_2_19_) );
DFFPOSX1 DFFPOSX1_804 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf144), .D(_4494__20_), .Q(H_2_20_) );
DFFPOSX1 DFFPOSX1_805 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf143), .D(_4494__21_), .Q(H_2_21_) );
DFFPOSX1 DFFPOSX1_806 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf142), .D(_4494__22_), .Q(H_2_22_) );
DFFPOSX1 DFFPOSX1_807 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf141), .D(_4494__23_), .Q(H_2_23_) );
DFFPOSX1 DFFPOSX1_808 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf140), .D(_4568_), .Q(comparador_2_valid_hash) );
DFFPOSX1 DFFPOSX1_809 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf139), .D(_4492__0_), .Q(micro_hash_ucr_2_b_0_) );
DFFPOSX1 DFFPOSX1_810 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf138), .D(_4492__1_), .Q(micro_hash_ucr_2_b_1_) );
DFFPOSX1 DFFPOSX1_811 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf137), .D(_4492__2_), .Q(micro_hash_ucr_2_b_2_) );
DFFPOSX1 DFFPOSX1_812 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf136), .D(_4492__3_), .Q(micro_hash_ucr_2_b_3_) );
DFFPOSX1 DFFPOSX1_813 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf135), .D(_4492__4_), .Q(micro_hash_ucr_2_b_4_) );
DFFPOSX1 DFFPOSX1_814 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf134), .D(_4492__5_), .Q(micro_hash_ucr_2_b_5_) );
DFFPOSX1 DFFPOSX1_815 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf133), .D(_4492__6_), .Q(micro_hash_ucr_2_b_6_) );
DFFPOSX1 DFFPOSX1_816 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf132), .D(_4492__7_), .Q(micro_hash_ucr_2_b_7_) );
DFFPOSX1 DFFPOSX1_817 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf131), .D(_4493__0_), .Q(micro_hash_ucr_2_c_0_) );
DFFPOSX1 DFFPOSX1_818 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf130), .D(_4493__1_), .Q(micro_hash_ucr_2_c_1_) );
DFFPOSX1 DFFPOSX1_819 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf129), .D(_4493__2_), .Q(micro_hash_ucr_2_c_2_) );
DFFPOSX1 DFFPOSX1_820 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf128), .D(_4493__3_), .Q(micro_hash_ucr_2_c_3_) );
DFFPOSX1 DFFPOSX1_821 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf127), .D(_4493__4_), .Q(micro_hash_ucr_2_c_4_) );
DFFPOSX1 DFFPOSX1_822 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf126), .D(_4493__5_), .Q(micro_hash_ucr_2_c_5_) );
DFFPOSX1 DFFPOSX1_823 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf125), .D(_4493__6_), .Q(micro_hash_ucr_2_c_6_) );
DFFPOSX1 DFFPOSX1_824 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf124), .D(_4493__7_), .Q(micro_hash_ucr_2_c_7_) );
DFFPOSX1 DFFPOSX1_825 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf123), .D(_4569__0_), .Q(micro_hash_ucr_2_x_0_) );
DFFPOSX1 DFFPOSX1_826 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf122), .D(_4569__1_), .Q(micro_hash_ucr_2_x_1_) );
DFFPOSX1 DFFPOSX1_827 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf121), .D(_4569__2_), .Q(micro_hash_ucr_2_x_2_) );
DFFPOSX1 DFFPOSX1_828 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf120), .D(_4569__3_), .Q(micro_hash_ucr_2_x_3_) );
DFFPOSX1 DFFPOSX1_829 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf119), .D(_4569__4_), .Q(micro_hash_ucr_2_x_4_) );
DFFPOSX1 DFFPOSX1_830 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf118), .D(_4569__5_), .Q(micro_hash_ucr_2_x_5_) );
DFFPOSX1 DFFPOSX1_831 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf117), .D(_4569__6_), .Q(micro_hash_ucr_2_x_6_) );
DFFPOSX1 DFFPOSX1_832 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf116), .D(_4569__7_), .Q(micro_hash_ucr_2_x_7_) );
DFFPOSX1 DFFPOSX1_833 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf115), .D(_4495__0_), .Q(micro_hash_ucr_2_k_0_) );
DFFPOSX1 DFFPOSX1_834 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf114), .D(_4495__1_), .Q(micro_hash_ucr_2_k_1_) );
DFFPOSX1 DFFPOSX1_835 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf113), .D(_4495__2_), .Q(micro_hash_ucr_2_k_2_) );
DFFPOSX1 DFFPOSX1_836 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf112), .D(_4495__3_), .Q(micro_hash_ucr_2_k_3_) );
DFFPOSX1 DFFPOSX1_837 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf111), .D(_4495__4_), .Q(micro_hash_ucr_2_k_4_) );
DFFPOSX1 DFFPOSX1_838 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf110), .D(_4495__5_), .Q(micro_hash_ucr_2_k_5_) );
DFFPOSX1 DFFPOSX1_839 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf109), .D(_4495__6_), .Q(micro_hash_ucr_2_k_6_) );
DFFPOSX1 DFFPOSX1_840 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf108), .D(_4495__7_), .Q(micro_hash_ucr_2_k_7_) );
DFFPOSX1 DFFPOSX1_841 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf107), .D(_4491__0_), .Q(micro_hash_ucr_2_a_0_) );
DFFPOSX1 DFFPOSX1_842 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(_4491__1_), .Q(micro_hash_ucr_2_a_1_) );
DFFPOSX1 DFFPOSX1_843 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(_4491__2_), .Q(micro_hash_ucr_2_a_2_) );
DFFPOSX1 DFFPOSX1_844 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(_4491__3_), .Q(micro_hash_ucr_2_a_3_) );
DFFPOSX1 DFFPOSX1_845 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(_4491__4_), .Q(micro_hash_ucr_2_a_4_) );
DFFPOSX1 DFFPOSX1_846 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(_4491__5_), .Q(micro_hash_ucr_2_a_5_) );
DFFPOSX1 DFFPOSX1_847 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(_4491__6_), .Q(micro_hash_ucr_2_a_6_) );
DFFPOSX1 DFFPOSX1_848 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(_4491__7_), .Q(micro_hash_ucr_2_a_7_) );
DFFPOSX1 DFFPOSX1_849 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(_4496__bF_buf0), .Q(micro_hash_ucr_2_pipe0) );
DFFPOSX1 DFFPOSX1_850 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_4490__0_), .Q(micro_hash_ucr_2_Wx_0_) );
DFFPOSX1 DFFPOSX1_851 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_4490__1_), .Q(micro_hash_ucr_2_Wx_1_) );
DFFPOSX1 DFFPOSX1_852 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_4490__2_), .Q(micro_hash_ucr_2_Wx_2_) );
DFFPOSX1 DFFPOSX1_853 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_4490__3_), .Q(micro_hash_ucr_2_Wx_3_) );
DFFPOSX1 DFFPOSX1_854 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_4490__4_), .Q(micro_hash_ucr_2_Wx_4_) );
DFFPOSX1 DFFPOSX1_855 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_4490__5_), .Q(micro_hash_ucr_2_Wx_5_) );
DFFPOSX1 DFFPOSX1_856 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_4490__6_), .Q(micro_hash_ucr_2_Wx_6_) );
DFFPOSX1 DFFPOSX1_857 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_4490__7_), .Q(micro_hash_ucr_2_Wx_7_) );
DFFPOSX1 DFFPOSX1_858 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_4490__8_), .Q(micro_hash_ucr_2_Wx_8_) );
DFFPOSX1 DFFPOSX1_859 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_4490__9_), .Q(micro_hash_ucr_2_Wx_9_) );
DFFPOSX1 DFFPOSX1_860 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_4490__10_), .Q(micro_hash_ucr_2_Wx_10_) );
DFFPOSX1 DFFPOSX1_861 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_4490__11_), .Q(micro_hash_ucr_2_Wx_11_) );
DFFPOSX1 DFFPOSX1_862 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_4490__12_), .Q(micro_hash_ucr_2_Wx_12_) );
DFFPOSX1 DFFPOSX1_863 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_4490__13_), .Q(micro_hash_ucr_2_Wx_13_) );
DFFPOSX1 DFFPOSX1_864 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_4490__14_), .Q(micro_hash_ucr_2_Wx_14_) );
DFFPOSX1 DFFPOSX1_865 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_4490__15_), .Q(micro_hash_ucr_2_Wx_15_) );
DFFPOSX1 DFFPOSX1_866 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_4490__16_), .Q(micro_hash_ucr_2_Wx_16_) );
DFFPOSX1 DFFPOSX1_867 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_4490__17_), .Q(micro_hash_ucr_2_Wx_17_) );
DFFPOSX1 DFFPOSX1_868 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_4490__18_), .Q(micro_hash_ucr_2_Wx_18_) );
DFFPOSX1 DFFPOSX1_869 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_4490__19_), .Q(micro_hash_ucr_2_Wx_19_) );
DFFPOSX1 DFFPOSX1_870 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_4490__20_), .Q(micro_hash_ucr_2_Wx_20_) );
DFFPOSX1 DFFPOSX1_871 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_4490__21_), .Q(micro_hash_ucr_2_Wx_21_) );
DFFPOSX1 DFFPOSX1_872 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_4490__22_), .Q(micro_hash_ucr_2_Wx_22_) );
DFFPOSX1 DFFPOSX1_873 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_4490__23_), .Q(micro_hash_ucr_2_Wx_23_) );
DFFPOSX1 DFFPOSX1_874 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_4490__24_), .Q(micro_hash_ucr_2_Wx_24_) );
DFFPOSX1 DFFPOSX1_875 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_4490__25_), .Q(micro_hash_ucr_2_Wx_25_) );
DFFPOSX1 DFFPOSX1_876 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_4490__26_), .Q(micro_hash_ucr_2_Wx_26_) );
DFFPOSX1 DFFPOSX1_877 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_4490__27_), .Q(micro_hash_ucr_2_Wx_27_) );
DFFPOSX1 DFFPOSX1_878 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_4490__28_), .Q(micro_hash_ucr_2_Wx_28_) );
DFFPOSX1 DFFPOSX1_879 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_4490__29_), .Q(micro_hash_ucr_2_Wx_29_) );
DFFPOSX1 DFFPOSX1_880 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_4490__30_), .Q(micro_hash_ucr_2_Wx_30_) );
DFFPOSX1 DFFPOSX1_881 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_4490__31_), .Q(micro_hash_ucr_2_Wx_31_) );
DFFPOSX1 DFFPOSX1_882 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_4490__32_), .Q(micro_hash_ucr_2_Wx_32_) );
DFFPOSX1 DFFPOSX1_883 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_4490__33_), .Q(micro_hash_ucr_2_Wx_33_) );
DFFPOSX1 DFFPOSX1_884 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_4490__34_), .Q(micro_hash_ucr_2_Wx_34_) );
DFFPOSX1 DFFPOSX1_885 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_4490__35_), .Q(micro_hash_ucr_2_Wx_35_) );
DFFPOSX1 DFFPOSX1_886 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_4490__36_), .Q(micro_hash_ucr_2_Wx_36_) );
DFFPOSX1 DFFPOSX1_887 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_4490__37_), .Q(micro_hash_ucr_2_Wx_37_) );
DFFPOSX1 DFFPOSX1_888 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_4490__38_), .Q(micro_hash_ucr_2_Wx_38_) );
DFFPOSX1 DFFPOSX1_889 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_4490__39_), .Q(micro_hash_ucr_2_Wx_39_) );
DFFPOSX1 DFFPOSX1_890 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_4490__40_), .Q(micro_hash_ucr_2_Wx_40_) );
DFFPOSX1 DFFPOSX1_891 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_4490__41_), .Q(micro_hash_ucr_2_Wx_41_) );
DFFPOSX1 DFFPOSX1_892 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_4490__42_), .Q(micro_hash_ucr_2_Wx_42_) );
DFFPOSX1 DFFPOSX1_893 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_4490__43_), .Q(micro_hash_ucr_2_Wx_43_) );
DFFPOSX1 DFFPOSX1_894 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_4490__44_), .Q(micro_hash_ucr_2_Wx_44_) );
DFFPOSX1 DFFPOSX1_895 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_4490__45_), .Q(micro_hash_ucr_2_Wx_45_) );
DFFPOSX1 DFFPOSX1_896 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_4490__46_), .Q(micro_hash_ucr_2_Wx_46_) );
DFFPOSX1 DFFPOSX1_897 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_4490__47_), .Q(micro_hash_ucr_2_Wx_47_) );
DFFPOSX1 DFFPOSX1_898 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_4490__48_), .Q(micro_hash_ucr_2_Wx_48_) );
DFFPOSX1 DFFPOSX1_899 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_4490__49_), .Q(micro_hash_ucr_2_Wx_49_) );
DFFPOSX1 DFFPOSX1_900 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_4490__50_), .Q(micro_hash_ucr_2_Wx_50_) );
DFFPOSX1 DFFPOSX1_901 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_4490__51_), .Q(micro_hash_ucr_2_Wx_51_) );
DFFPOSX1 DFFPOSX1_902 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_4490__52_), .Q(micro_hash_ucr_2_Wx_52_) );
DFFPOSX1 DFFPOSX1_903 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_4490__53_), .Q(micro_hash_ucr_2_Wx_53_) );
DFFPOSX1 DFFPOSX1_904 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_4490__54_), .Q(micro_hash_ucr_2_Wx_54_) );
DFFPOSX1 DFFPOSX1_905 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_4490__55_), .Q(micro_hash_ucr_2_Wx_55_) );
DFFPOSX1 DFFPOSX1_906 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_4490__56_), .Q(micro_hash_ucr_2_Wx_56_) );
DFFPOSX1 DFFPOSX1_907 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_4490__57_), .Q(micro_hash_ucr_2_Wx_57_) );
DFFPOSX1 DFFPOSX1_908 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_4490__58_), .Q(micro_hash_ucr_2_Wx_58_) );
DFFPOSX1 DFFPOSX1_909 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_4490__59_), .Q(micro_hash_ucr_2_Wx_59_) );
DFFPOSX1 DFFPOSX1_910 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_4490__60_), .Q(micro_hash_ucr_2_Wx_60_) );
DFFPOSX1 DFFPOSX1_911 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_4490__61_), .Q(micro_hash_ucr_2_Wx_61_) );
DFFPOSX1 DFFPOSX1_912 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_4490__62_), .Q(micro_hash_ucr_2_Wx_62_) );
DFFPOSX1 DFFPOSX1_913 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_4490__63_), .Q(micro_hash_ucr_2_Wx_63_) );
DFFPOSX1 DFFPOSX1_914 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_4490__64_), .Q(micro_hash_ucr_2_Wx_64_) );
DFFPOSX1 DFFPOSX1_915 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_4490__65_), .Q(micro_hash_ucr_2_Wx_65_) );
DFFPOSX1 DFFPOSX1_916 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_4490__66_), .Q(micro_hash_ucr_2_Wx_66_) );
DFFPOSX1 DFFPOSX1_917 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_4490__67_), .Q(micro_hash_ucr_2_Wx_67_) );
DFFPOSX1 DFFPOSX1_918 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_4490__68_), .Q(micro_hash_ucr_2_Wx_68_) );
DFFPOSX1 DFFPOSX1_919 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_4490__69_), .Q(micro_hash_ucr_2_Wx_69_) );
DFFPOSX1 DFFPOSX1_920 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_4490__70_), .Q(micro_hash_ucr_2_Wx_70_) );
DFFPOSX1 DFFPOSX1_921 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_4490__71_), .Q(micro_hash_ucr_2_Wx_71_) );
DFFPOSX1 DFFPOSX1_922 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_4490__72_), .Q(micro_hash_ucr_2_Wx_72_) );
DFFPOSX1 DFFPOSX1_923 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_4490__73_), .Q(micro_hash_ucr_2_Wx_73_) );
DFFPOSX1 DFFPOSX1_924 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_4490__74_), .Q(micro_hash_ucr_2_Wx_74_) );
DFFPOSX1 DFFPOSX1_925 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_4490__75_), .Q(micro_hash_ucr_2_Wx_75_) );
DFFPOSX1 DFFPOSX1_926 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_4490__76_), .Q(micro_hash_ucr_2_Wx_76_) );
DFFPOSX1 DFFPOSX1_927 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_4490__77_), .Q(micro_hash_ucr_2_Wx_77_) );
DFFPOSX1 DFFPOSX1_928 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_4490__78_), .Q(micro_hash_ucr_2_Wx_78_) );
DFFPOSX1 DFFPOSX1_929 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_4490__79_), .Q(micro_hash_ucr_2_Wx_79_) );
DFFPOSX1 DFFPOSX1_930 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_4490__80_), .Q(micro_hash_ucr_2_Wx_80_) );
DFFPOSX1 DFFPOSX1_931 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_4490__81_), .Q(micro_hash_ucr_2_Wx_81_) );
DFFPOSX1 DFFPOSX1_932 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_4490__82_), .Q(micro_hash_ucr_2_Wx_82_) );
DFFPOSX1 DFFPOSX1_933 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_4490__83_), .Q(micro_hash_ucr_2_Wx_83_) );
DFFPOSX1 DFFPOSX1_934 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_4490__84_), .Q(micro_hash_ucr_2_Wx_84_) );
DFFPOSX1 DFFPOSX1_935 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_4490__85_), .Q(micro_hash_ucr_2_Wx_85_) );
DFFPOSX1 DFFPOSX1_936 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_4490__86_), .Q(micro_hash_ucr_2_Wx_86_) );
DFFPOSX1 DFFPOSX1_937 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_4490__87_), .Q(micro_hash_ucr_2_Wx_87_) );
DFFPOSX1 DFFPOSX1_938 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_4490__88_), .Q(micro_hash_ucr_2_Wx_88_) );
DFFPOSX1 DFFPOSX1_939 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_4490__89_), .Q(micro_hash_ucr_2_Wx_89_) );
DFFPOSX1 DFFPOSX1_940 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_4490__90_), .Q(micro_hash_ucr_2_Wx_90_) );
DFFPOSX1 DFFPOSX1_941 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_4490__91_), .Q(micro_hash_ucr_2_Wx_91_) );
DFFPOSX1 DFFPOSX1_942 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_4490__92_), .Q(micro_hash_ucr_2_Wx_92_) );
DFFPOSX1 DFFPOSX1_943 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_4490__93_), .Q(micro_hash_ucr_2_Wx_93_) );
DFFPOSX1 DFFPOSX1_944 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_4490__94_), .Q(micro_hash_ucr_2_Wx_94_) );
DFFPOSX1 DFFPOSX1_945 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_4490__95_), .Q(micro_hash_ucr_2_Wx_95_) );
DFFPOSX1 DFFPOSX1_946 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_4490__96_), .Q(micro_hash_ucr_2_Wx_96_) );
DFFPOSX1 DFFPOSX1_947 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_4490__97_), .Q(micro_hash_ucr_2_Wx_97_) );
DFFPOSX1 DFFPOSX1_948 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_4490__98_), .Q(micro_hash_ucr_2_Wx_98_) );
DFFPOSX1 DFFPOSX1_949 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf157), .D(_4490__99_), .Q(micro_hash_ucr_2_Wx_99_) );
DFFPOSX1 DFFPOSX1_950 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf156), .D(_4490__100_), .Q(micro_hash_ucr_2_Wx_100_) );
DFFPOSX1 DFFPOSX1_951 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf155), .D(_4490__101_), .Q(micro_hash_ucr_2_Wx_101_) );
DFFPOSX1 DFFPOSX1_952 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf154), .D(_4490__102_), .Q(micro_hash_ucr_2_Wx_102_) );
DFFPOSX1 DFFPOSX1_953 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf153), .D(_4490__103_), .Q(micro_hash_ucr_2_Wx_103_) );
DFFPOSX1 DFFPOSX1_954 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf152), .D(_4490__104_), .Q(micro_hash_ucr_2_Wx_104_) );
DFFPOSX1 DFFPOSX1_955 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf151), .D(_4490__105_), .Q(micro_hash_ucr_2_Wx_105_) );
DFFPOSX1 DFFPOSX1_956 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf150), .D(_4490__106_), .Q(micro_hash_ucr_2_Wx_106_) );
DFFPOSX1 DFFPOSX1_957 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf149), .D(_4490__107_), .Q(micro_hash_ucr_2_Wx_107_) );
DFFPOSX1 DFFPOSX1_958 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf148), .D(_4490__108_), .Q(micro_hash_ucr_2_Wx_108_) );
DFFPOSX1 DFFPOSX1_959 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf147), .D(_4490__109_), .Q(micro_hash_ucr_2_Wx_109_) );
DFFPOSX1 DFFPOSX1_960 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf146), .D(_4490__110_), .Q(micro_hash_ucr_2_Wx_110_) );
DFFPOSX1 DFFPOSX1_961 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf145), .D(_4490__111_), .Q(micro_hash_ucr_2_Wx_111_) );
DFFPOSX1 DFFPOSX1_962 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf144), .D(_4490__112_), .Q(micro_hash_ucr_2_Wx_112_) );
DFFPOSX1 DFFPOSX1_963 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf143), .D(_4490__113_), .Q(micro_hash_ucr_2_Wx_113_) );
DFFPOSX1 DFFPOSX1_964 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf142), .D(_4490__114_), .Q(micro_hash_ucr_2_Wx_114_) );
DFFPOSX1 DFFPOSX1_965 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf141), .D(_4490__115_), .Q(micro_hash_ucr_2_Wx_115_) );
DFFPOSX1 DFFPOSX1_966 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf140), .D(_4490__116_), .Q(micro_hash_ucr_2_Wx_116_) );
DFFPOSX1 DFFPOSX1_967 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf139), .D(_4490__117_), .Q(micro_hash_ucr_2_Wx_117_) );
DFFPOSX1 DFFPOSX1_968 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf138), .D(_4490__118_), .Q(micro_hash_ucr_2_Wx_118_) );
DFFPOSX1 DFFPOSX1_969 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf137), .D(_4490__119_), .Q(micro_hash_ucr_2_Wx_119_) );
DFFPOSX1 DFFPOSX1_970 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf136), .D(_4490__120_), .Q(micro_hash_ucr_2_Wx_120_) );
DFFPOSX1 DFFPOSX1_971 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf135), .D(_4490__121_), .Q(micro_hash_ucr_2_Wx_121_) );
DFFPOSX1 DFFPOSX1_972 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf134), .D(_4490__122_), .Q(micro_hash_ucr_2_Wx_122_) );
DFFPOSX1 DFFPOSX1_973 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf133), .D(_4490__123_), .Q(micro_hash_ucr_2_Wx_123_) );
DFFPOSX1 DFFPOSX1_974 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf132), .D(_4490__124_), .Q(micro_hash_ucr_2_Wx_124_) );
DFFPOSX1 DFFPOSX1_975 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf131), .D(_4490__125_), .Q(micro_hash_ucr_2_Wx_125_) );
DFFPOSX1 DFFPOSX1_976 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf130), .D(_4490__126_), .Q(micro_hash_ucr_2_Wx_126_) );
DFFPOSX1 DFFPOSX1_977 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf129), .D(_4490__127_), .Q(micro_hash_ucr_2_Wx_127_) );
DFFPOSX1 DFFPOSX1_978 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf128), .D(_4490__128_), .Q(micro_hash_ucr_2_Wx_128_) );
DFFPOSX1 DFFPOSX1_979 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf127), .D(_4490__129_), .Q(micro_hash_ucr_2_Wx_129_) );
DFFPOSX1 DFFPOSX1_980 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf126), .D(_4490__130_), .Q(micro_hash_ucr_2_Wx_130_) );
DFFPOSX1 DFFPOSX1_981 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf125), .D(_4490__131_), .Q(micro_hash_ucr_2_Wx_131_) );
DFFPOSX1 DFFPOSX1_982 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf124), .D(_4490__132_), .Q(micro_hash_ucr_2_Wx_132_) );
DFFPOSX1 DFFPOSX1_983 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf123), .D(_4490__133_), .Q(micro_hash_ucr_2_Wx_133_) );
DFFPOSX1 DFFPOSX1_984 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf122), .D(_4490__134_), .Q(micro_hash_ucr_2_Wx_134_) );
DFFPOSX1 DFFPOSX1_985 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf121), .D(_4490__135_), .Q(micro_hash_ucr_2_Wx_135_) );
DFFPOSX1 DFFPOSX1_986 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf120), .D(_4490__136_), .Q(micro_hash_ucr_2_Wx_136_) );
DFFPOSX1 DFFPOSX1_987 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf119), .D(_4490__137_), .Q(micro_hash_ucr_2_Wx_137_) );
DFFPOSX1 DFFPOSX1_988 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf118), .D(_4490__138_), .Q(micro_hash_ucr_2_Wx_138_) );
DFFPOSX1 DFFPOSX1_989 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf117), .D(_4490__139_), .Q(micro_hash_ucr_2_Wx_139_) );
DFFPOSX1 DFFPOSX1_990 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf116), .D(_4490__140_), .Q(micro_hash_ucr_2_Wx_140_) );
DFFPOSX1 DFFPOSX1_991 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf115), .D(_4490__141_), .Q(micro_hash_ucr_2_Wx_141_) );
DFFPOSX1 DFFPOSX1_992 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf114), .D(_4490__142_), .Q(micro_hash_ucr_2_Wx_142_) );
DFFPOSX1 DFFPOSX1_993 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf113), .D(_4490__143_), .Q(micro_hash_ucr_2_Wx_143_) );
DFFPOSX1 DFFPOSX1_994 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf112), .D(_4490__144_), .Q(micro_hash_ucr_2_Wx_144_) );
DFFPOSX1 DFFPOSX1_995 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf111), .D(_4490__145_), .Q(micro_hash_ucr_2_Wx_145_) );
DFFPOSX1 DFFPOSX1_996 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf110), .D(_4490__146_), .Q(micro_hash_ucr_2_Wx_146_) );
DFFPOSX1 DFFPOSX1_997 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf109), .D(_4490__147_), .Q(micro_hash_ucr_2_Wx_147_) );
DFFPOSX1 DFFPOSX1_998 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf108), .D(_4490__148_), .Q(micro_hash_ucr_2_Wx_148_) );
DFFPOSX1 DFFPOSX1_999 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf107), .D(_4490__149_), .Q(micro_hash_ucr_2_Wx_149_) );
DFFPOSX1 DFFPOSX1_1000 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(_4490__150_), .Q(micro_hash_ucr_2_Wx_150_) );
DFFPOSX1 DFFPOSX1_1001 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(_4490__151_), .Q(micro_hash_ucr_2_Wx_151_) );
DFFPOSX1 DFFPOSX1_1002 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(_4490__152_), .Q(micro_hash_ucr_2_Wx_152_) );
DFFPOSX1 DFFPOSX1_1003 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(_4490__153_), .Q(micro_hash_ucr_2_Wx_153_) );
DFFPOSX1 DFFPOSX1_1004 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(_4490__154_), .Q(micro_hash_ucr_2_Wx_154_) );
DFFPOSX1 DFFPOSX1_1005 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(_4490__155_), .Q(micro_hash_ucr_2_Wx_155_) );
DFFPOSX1 DFFPOSX1_1006 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(_4490__156_), .Q(micro_hash_ucr_2_Wx_156_) );
DFFPOSX1 DFFPOSX1_1007 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(_4490__157_), .Q(micro_hash_ucr_2_Wx_157_) );
DFFPOSX1 DFFPOSX1_1008 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_4490__158_), .Q(micro_hash_ucr_2_Wx_158_) );
DFFPOSX1 DFFPOSX1_1009 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_4490__159_), .Q(micro_hash_ucr_2_Wx_159_) );
DFFPOSX1 DFFPOSX1_1010 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_4490__160_), .Q(micro_hash_ucr_2_Wx_160_) );
DFFPOSX1 DFFPOSX1_1011 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_4490__161_), .Q(micro_hash_ucr_2_Wx_161_) );
DFFPOSX1 DFFPOSX1_1012 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_4490__162_), .Q(micro_hash_ucr_2_Wx_162_) );
DFFPOSX1 DFFPOSX1_1013 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_4490__163_), .Q(micro_hash_ucr_2_Wx_163_) );
DFFPOSX1 DFFPOSX1_1014 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_4490__164_), .Q(micro_hash_ucr_2_Wx_164_) );
DFFPOSX1 DFFPOSX1_1015 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_4490__165_), .Q(micro_hash_ucr_2_Wx_165_) );
DFFPOSX1 DFFPOSX1_1016 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_4490__166_), .Q(micro_hash_ucr_2_Wx_166_) );
DFFPOSX1 DFFPOSX1_1017 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_4490__167_), .Q(micro_hash_ucr_2_Wx_167_) );
DFFPOSX1 DFFPOSX1_1018 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_4490__168_), .Q(micro_hash_ucr_2_Wx_168_) );
DFFPOSX1 DFFPOSX1_1019 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_4490__169_), .Q(micro_hash_ucr_2_Wx_169_) );
DFFPOSX1 DFFPOSX1_1020 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_4490__170_), .Q(micro_hash_ucr_2_Wx_170_) );
DFFPOSX1 DFFPOSX1_1021 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_4490__171_), .Q(micro_hash_ucr_2_Wx_171_) );
DFFPOSX1 DFFPOSX1_1022 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_4490__172_), .Q(micro_hash_ucr_2_Wx_172_) );
DFFPOSX1 DFFPOSX1_1023 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_4490__173_), .Q(micro_hash_ucr_2_Wx_173_) );
DFFPOSX1 DFFPOSX1_1024 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_4490__174_), .Q(micro_hash_ucr_2_Wx_174_) );
DFFPOSX1 DFFPOSX1_1025 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_4490__175_), .Q(micro_hash_ucr_2_Wx_175_) );
DFFPOSX1 DFFPOSX1_1026 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_4490__176_), .Q(micro_hash_ucr_2_Wx_176_) );
DFFPOSX1 DFFPOSX1_1027 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_4490__177_), .Q(micro_hash_ucr_2_Wx_177_) );
DFFPOSX1 DFFPOSX1_1028 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_4490__178_), .Q(micro_hash_ucr_2_Wx_178_) );
DFFPOSX1 DFFPOSX1_1029 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_4490__179_), .Q(micro_hash_ucr_2_Wx_179_) );
DFFPOSX1 DFFPOSX1_1030 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_4490__180_), .Q(micro_hash_ucr_2_Wx_180_) );
DFFPOSX1 DFFPOSX1_1031 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_4490__181_), .Q(micro_hash_ucr_2_Wx_181_) );
DFFPOSX1 DFFPOSX1_1032 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_4490__182_), .Q(micro_hash_ucr_2_Wx_182_) );
DFFPOSX1 DFFPOSX1_1033 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_4490__183_), .Q(micro_hash_ucr_2_Wx_183_) );
DFFPOSX1 DFFPOSX1_1034 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_4490__184_), .Q(micro_hash_ucr_2_Wx_184_) );
DFFPOSX1 DFFPOSX1_1035 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_4490__185_), .Q(micro_hash_ucr_2_Wx_185_) );
DFFPOSX1 DFFPOSX1_1036 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_4490__186_), .Q(micro_hash_ucr_2_Wx_186_) );
DFFPOSX1 DFFPOSX1_1037 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_4490__187_), .Q(micro_hash_ucr_2_Wx_187_) );
DFFPOSX1 DFFPOSX1_1038 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_4490__188_), .Q(micro_hash_ucr_2_Wx_188_) );
DFFPOSX1 DFFPOSX1_1039 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_4490__189_), .Q(micro_hash_ucr_2_Wx_189_) );
DFFPOSX1 DFFPOSX1_1040 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_4490__190_), .Q(micro_hash_ucr_2_Wx_190_) );
DFFPOSX1 DFFPOSX1_1041 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_4490__191_), .Q(micro_hash_ucr_2_Wx_191_) );
DFFPOSX1 DFFPOSX1_1042 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_4490__192_), .Q(micro_hash_ucr_2_Wx_192_) );
DFFPOSX1 DFFPOSX1_1043 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_4490__193_), .Q(micro_hash_ucr_2_Wx_193_) );
DFFPOSX1 DFFPOSX1_1044 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_4490__194_), .Q(micro_hash_ucr_2_Wx_194_) );
DFFPOSX1 DFFPOSX1_1045 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_4490__195_), .Q(micro_hash_ucr_2_Wx_195_) );
DFFPOSX1 DFFPOSX1_1046 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_4490__196_), .Q(micro_hash_ucr_2_Wx_196_) );
DFFPOSX1 DFFPOSX1_1047 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_4490__197_), .Q(micro_hash_ucr_2_Wx_197_) );
DFFPOSX1 DFFPOSX1_1048 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_4490__198_), .Q(micro_hash_ucr_2_Wx_198_) );
DFFPOSX1 DFFPOSX1_1049 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_4490__199_), .Q(micro_hash_ucr_2_Wx_199_) );
DFFPOSX1 DFFPOSX1_1050 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_4490__200_), .Q(micro_hash_ucr_2_Wx_200_) );
DFFPOSX1 DFFPOSX1_1051 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_4490__201_), .Q(micro_hash_ucr_2_Wx_201_) );
DFFPOSX1 DFFPOSX1_1052 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_4490__202_), .Q(micro_hash_ucr_2_Wx_202_) );
DFFPOSX1 DFFPOSX1_1053 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_4490__203_), .Q(micro_hash_ucr_2_Wx_203_) );
DFFPOSX1 DFFPOSX1_1054 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_4490__204_), .Q(micro_hash_ucr_2_Wx_204_) );
DFFPOSX1 DFFPOSX1_1055 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_4490__205_), .Q(micro_hash_ucr_2_Wx_205_) );
DFFPOSX1 DFFPOSX1_1056 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_4490__206_), .Q(micro_hash_ucr_2_Wx_206_) );
DFFPOSX1 DFFPOSX1_1057 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_4490__207_), .Q(micro_hash_ucr_2_Wx_207_) );
DFFPOSX1 DFFPOSX1_1058 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_4490__208_), .Q(micro_hash_ucr_2_Wx_208_) );
DFFPOSX1 DFFPOSX1_1059 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_4490__209_), .Q(micro_hash_ucr_2_Wx_209_) );
DFFPOSX1 DFFPOSX1_1060 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_4490__210_), .Q(micro_hash_ucr_2_Wx_210_) );
DFFPOSX1 DFFPOSX1_1061 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_4490__211_), .Q(micro_hash_ucr_2_Wx_211_) );
DFFPOSX1 DFFPOSX1_1062 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_4490__212_), .Q(micro_hash_ucr_2_Wx_212_) );
DFFPOSX1 DFFPOSX1_1063 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_4490__213_), .Q(micro_hash_ucr_2_Wx_213_) );
DFFPOSX1 DFFPOSX1_1064 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_4490__214_), .Q(micro_hash_ucr_2_Wx_214_) );
DFFPOSX1 DFFPOSX1_1065 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_4490__215_), .Q(micro_hash_ucr_2_Wx_215_) );
DFFPOSX1 DFFPOSX1_1066 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_4490__216_), .Q(micro_hash_ucr_2_Wx_216_) );
DFFPOSX1 DFFPOSX1_1067 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_4490__217_), .Q(micro_hash_ucr_2_Wx_217_) );
DFFPOSX1 DFFPOSX1_1068 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_4490__218_), .Q(micro_hash_ucr_2_Wx_218_) );
DFFPOSX1 DFFPOSX1_1069 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_4490__219_), .Q(micro_hash_ucr_2_Wx_219_) );
DFFPOSX1 DFFPOSX1_1070 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_4490__220_), .Q(micro_hash_ucr_2_Wx_220_) );
DFFPOSX1 DFFPOSX1_1071 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_4490__221_), .Q(micro_hash_ucr_2_Wx_221_) );
DFFPOSX1 DFFPOSX1_1072 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_4490__222_), .Q(micro_hash_ucr_2_Wx_222_) );
DFFPOSX1 DFFPOSX1_1073 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_4490__223_), .Q(micro_hash_ucr_2_Wx_223_) );
DFFPOSX1 DFFPOSX1_1074 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_4490__224_), .Q(micro_hash_ucr_2_Wx_224_) );
DFFPOSX1 DFFPOSX1_1075 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_4490__225_), .Q(micro_hash_ucr_2_Wx_225_) );
DFFPOSX1 DFFPOSX1_1076 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_4490__226_), .Q(micro_hash_ucr_2_Wx_226_) );
DFFPOSX1 DFFPOSX1_1077 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_4490__227_), .Q(micro_hash_ucr_2_Wx_227_) );
DFFPOSX1 DFFPOSX1_1078 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_4490__228_), .Q(micro_hash_ucr_2_Wx_228_) );
DFFPOSX1 DFFPOSX1_1079 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_4490__229_), .Q(micro_hash_ucr_2_Wx_229_) );
DFFPOSX1 DFFPOSX1_1080 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_4490__230_), .Q(micro_hash_ucr_2_Wx_230_) );
DFFPOSX1 DFFPOSX1_1081 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_4490__231_), .Q(micro_hash_ucr_2_Wx_231_) );
DFFPOSX1 DFFPOSX1_1082 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_4490__232_), .Q(micro_hash_ucr_2_Wx_232_) );
DFFPOSX1 DFFPOSX1_1083 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_4490__233_), .Q(micro_hash_ucr_2_Wx_233_) );
DFFPOSX1 DFFPOSX1_1084 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_4490__234_), .Q(micro_hash_ucr_2_Wx_234_) );
DFFPOSX1 DFFPOSX1_1085 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_4490__235_), .Q(micro_hash_ucr_2_Wx_235_) );
DFFPOSX1 DFFPOSX1_1086 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_4490__236_), .Q(micro_hash_ucr_2_Wx_236_) );
DFFPOSX1 DFFPOSX1_1087 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_4490__237_), .Q(micro_hash_ucr_2_Wx_237_) );
DFFPOSX1 DFFPOSX1_1088 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_4490__238_), .Q(micro_hash_ucr_2_Wx_238_) );
DFFPOSX1 DFFPOSX1_1089 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_4490__239_), .Q(micro_hash_ucr_2_Wx_239_) );
DFFPOSX1 DFFPOSX1_1090 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_4490__240_), .Q(micro_hash_ucr_2_Wx_240_) );
DFFPOSX1 DFFPOSX1_1091 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_4490__241_), .Q(micro_hash_ucr_2_Wx_241_) );
DFFPOSX1 DFFPOSX1_1092 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_4490__242_), .Q(micro_hash_ucr_2_Wx_242_) );
DFFPOSX1 DFFPOSX1_1093 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_4490__243_), .Q(micro_hash_ucr_2_Wx_243_) );
DFFPOSX1 DFFPOSX1_1094 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_4490__244_), .Q(micro_hash_ucr_2_Wx_244_) );
DFFPOSX1 DFFPOSX1_1095 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_4490__245_), .Q(micro_hash_ucr_2_Wx_245_) );
DFFPOSX1 DFFPOSX1_1096 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_4490__246_), .Q(micro_hash_ucr_2_Wx_246_) );
DFFPOSX1 DFFPOSX1_1097 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_4490__247_), .Q(micro_hash_ucr_2_Wx_247_) );
DFFPOSX1 DFFPOSX1_1098 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_4490__248_), .Q(micro_hash_ucr_2_Wx_248_) );
DFFPOSX1 DFFPOSX1_1099 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_4490__249_), .Q(micro_hash_ucr_2_Wx_249_) );
DFFPOSX1 DFFPOSX1_1100 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_4490__250_), .Q(micro_hash_ucr_2_Wx_250_) );
DFFPOSX1 DFFPOSX1_1101 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_4490__251_), .Q(micro_hash_ucr_2_Wx_251_) );
DFFPOSX1 DFFPOSX1_1102 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_4490__252_), .Q(micro_hash_ucr_2_Wx_252_) );
DFFPOSX1 DFFPOSX1_1103 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_4490__253_), .Q(micro_hash_ucr_2_Wx_253_) );
DFFPOSX1 DFFPOSX1_1104 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_4490__254_), .Q(micro_hash_ucr_2_Wx_254_) );
DFFPOSX1 DFFPOSX1_1105 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_4490__255_), .Q(micro_hash_ucr_2_Wx_255_) );
DFFPOSX1 DFFPOSX1_1106 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_4507_), .Q(micro_hash_ucr_2_pipe1) );
DFFPOSX1 DFFPOSX1_1107 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf157), .D(_4518_), .Q(micro_hash_ucr_2_pipe2) );
DFFPOSX1 DFFPOSX1_1108 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf156), .D(_4529_), .Q(micro_hash_ucr_2_pipe3) );
DFFPOSX1 DFFPOSX1_1109 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf155), .D(_4540_), .Q(micro_hash_ucr_2_pipe4) );
DFFPOSX1 DFFPOSX1_1110 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf154), .D(_4551_), .Q(micro_hash_ucr_2_pipe5) );
DFFPOSX1 DFFPOSX1_1111 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf153), .D(_4562_), .Q(micro_hash_ucr_2_pipe6) );
DFFPOSX1 DFFPOSX1_1112 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf152), .D(_4565_), .Q(micro_hash_ucr_2_pipe7) );
DFFPOSX1 DFFPOSX1_1113 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf151), .D(_4566_), .Q(micro_hash_ucr_2_pipe8) );
DFFPOSX1 DFFPOSX1_1114 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf150), .D(_4567_), .Q(micro_hash_ucr_2_pipe9) );
DFFPOSX1 DFFPOSX1_1115 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf149), .D(_4497_), .Q(micro_hash_ucr_2_pipe10) );
DFFPOSX1 DFFPOSX1_1116 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf148), .D(_4498_), .Q(micro_hash_ucr_2_pipe11) );
DFFPOSX1 DFFPOSX1_1117 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf147), .D(_4499_), .Q(micro_hash_ucr_2_pipe12) );
DFFPOSX1 DFFPOSX1_1118 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf146), .D(_4500_), .Q(micro_hash_ucr_2_pipe13) );
DFFPOSX1 DFFPOSX1_1119 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf145), .D(_4501_), .Q(micro_hash_ucr_2_pipe14) );
DFFPOSX1 DFFPOSX1_1120 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf144), .D(_4502_), .Q(micro_hash_ucr_2_pipe15) );
DFFPOSX1 DFFPOSX1_1121 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf143), .D(_4503_), .Q(micro_hash_ucr_2_pipe16) );
DFFPOSX1 DFFPOSX1_1122 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf142), .D(_4504_), .Q(micro_hash_ucr_2_pipe17) );
DFFPOSX1 DFFPOSX1_1123 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf141), .D(_4505_), .Q(micro_hash_ucr_2_pipe18) );
DFFPOSX1 DFFPOSX1_1124 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf140), .D(_4506_), .Q(micro_hash_ucr_2_pipe19) );
DFFPOSX1 DFFPOSX1_1125 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf139), .D(_4508_), .Q(micro_hash_ucr_2_pipe20) );
DFFPOSX1 DFFPOSX1_1126 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf138), .D(_4509_), .Q(micro_hash_ucr_2_pipe21) );
DFFPOSX1 DFFPOSX1_1127 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf137), .D(_4510_), .Q(micro_hash_ucr_2_pipe22) );
DFFPOSX1 DFFPOSX1_1128 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf136), .D(_4511_), .Q(micro_hash_ucr_2_pipe23) );
DFFPOSX1 DFFPOSX1_1129 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf135), .D(_4512_), .Q(micro_hash_ucr_2_pipe24) );
DFFPOSX1 DFFPOSX1_1130 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf134), .D(_4513_), .Q(micro_hash_ucr_2_pipe25) );
DFFPOSX1 DFFPOSX1_1131 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf133), .D(_4514_), .Q(micro_hash_ucr_2_pipe26) );
DFFPOSX1 DFFPOSX1_1132 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf132), .D(_4515_), .Q(micro_hash_ucr_2_pipe27) );
DFFPOSX1 DFFPOSX1_1133 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf131), .D(_4516_), .Q(micro_hash_ucr_2_pipe28) );
DFFPOSX1 DFFPOSX1_1134 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf130), .D(_4517_), .Q(micro_hash_ucr_2_pipe29) );
DFFPOSX1 DFFPOSX1_1135 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf129), .D(_4519_), .Q(micro_hash_ucr_2_pipe30) );
DFFPOSX1 DFFPOSX1_1136 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf128), .D(_4520_), .Q(micro_hash_ucr_2_pipe31) );
DFFPOSX1 DFFPOSX1_1137 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf127), .D(_4521_), .Q(micro_hash_ucr_2_pipe32) );
DFFPOSX1 DFFPOSX1_1138 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf126), .D(_4522_), .Q(micro_hash_ucr_2_pipe33) );
DFFPOSX1 DFFPOSX1_1139 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf125), .D(_4523_), .Q(micro_hash_ucr_2_pipe34) );
DFFPOSX1 DFFPOSX1_1140 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf124), .D(_4524_), .Q(micro_hash_ucr_2_pipe35) );
DFFPOSX1 DFFPOSX1_1141 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf123), .D(_4525_), .Q(micro_hash_ucr_2_pipe36) );
DFFPOSX1 DFFPOSX1_1142 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf122), .D(_4526_), .Q(micro_hash_ucr_2_pipe37) );
DFFPOSX1 DFFPOSX1_1143 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf121), .D(_4527_), .Q(micro_hash_ucr_2_pipe38) );
DFFPOSX1 DFFPOSX1_1144 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf120), .D(_4528_), .Q(micro_hash_ucr_2_pipe39) );
DFFPOSX1 DFFPOSX1_1145 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf119), .D(_4530_), .Q(micro_hash_ucr_2_pipe40) );
DFFPOSX1 DFFPOSX1_1146 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf118), .D(_4531_), .Q(micro_hash_ucr_2_pipe41) );
DFFPOSX1 DFFPOSX1_1147 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf117), .D(_4532_), .Q(micro_hash_ucr_2_pipe42) );
DFFPOSX1 DFFPOSX1_1148 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf116), .D(_4533_), .Q(micro_hash_ucr_2_pipe43) );
DFFPOSX1 DFFPOSX1_1149 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf115), .D(_4534_), .Q(micro_hash_ucr_2_pipe44) );
DFFPOSX1 DFFPOSX1_1150 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf114), .D(_4535_), .Q(micro_hash_ucr_2_pipe45) );
DFFPOSX1 DFFPOSX1_1151 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf113), .D(_4536_), .Q(micro_hash_ucr_2_pipe46) );
DFFPOSX1 DFFPOSX1_1152 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf112), .D(_4537_), .Q(micro_hash_ucr_2_pipe47) );
DFFPOSX1 DFFPOSX1_1153 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf111), .D(_4538_), .Q(micro_hash_ucr_2_pipe48) );
DFFPOSX1 DFFPOSX1_1154 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf110), .D(_4539_), .Q(micro_hash_ucr_2_pipe49) );
DFFPOSX1 DFFPOSX1_1155 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf109), .D(_4541_), .Q(micro_hash_ucr_2_pipe50) );
DFFPOSX1 DFFPOSX1_1156 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf108), .D(_4542_), .Q(micro_hash_ucr_2_pipe51) );
DFFPOSX1 DFFPOSX1_1157 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf107), .D(_4543_), .Q(micro_hash_ucr_2_pipe52) );
DFFPOSX1 DFFPOSX1_1158 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(_4544_), .Q(micro_hash_ucr_2_pipe53) );
DFFPOSX1 DFFPOSX1_1159 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(_4545_), .Q(micro_hash_ucr_2_pipe54) );
DFFPOSX1 DFFPOSX1_1160 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(_4546_), .Q(micro_hash_ucr_2_pipe55) );
DFFPOSX1 DFFPOSX1_1161 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(_4547_), .Q(micro_hash_ucr_2_pipe56) );
DFFPOSX1 DFFPOSX1_1162 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(_4548_), .Q(micro_hash_ucr_2_pipe57) );
DFFPOSX1 DFFPOSX1_1163 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(_4549_), .Q(micro_hash_ucr_2_pipe58) );
DFFPOSX1 DFFPOSX1_1164 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(_4550_), .Q(micro_hash_ucr_2_pipe59) );
DFFPOSX1 DFFPOSX1_1165 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(_4552_), .Q(micro_hash_ucr_2_pipe60) );
DFFPOSX1 DFFPOSX1_1166 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_4553_), .Q(micro_hash_ucr_2_pipe61) );
DFFPOSX1 DFFPOSX1_1167 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_4554_), .Q(micro_hash_ucr_2_pipe62) );
DFFPOSX1 DFFPOSX1_1168 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_4555_), .Q(micro_hash_ucr_2_pipe63) );
DFFPOSX1 DFFPOSX1_1169 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_4556_), .Q(micro_hash_ucr_2_pipe64) );
DFFPOSX1 DFFPOSX1_1170 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_4557_), .Q(micro_hash_ucr_2_pipe65) );
DFFPOSX1 DFFPOSX1_1171 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_4558_), .Q(micro_hash_ucr_2_pipe66) );
DFFPOSX1 DFFPOSX1_1172 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_4559_), .Q(micro_hash_ucr_2_pipe67) );
DFFPOSX1 DFFPOSX1_1173 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_4560_), .Q(micro_hash_ucr_2_pipe68) );
DFFPOSX1 DFFPOSX1_1174 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_4561_), .Q(micro_hash_ucr_2_pipe69) );
DFFPOSX1 DFFPOSX1_1175 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_4563_), .Q(micro_hash_ucr_2_pipe70) );
DFFPOSX1 DFFPOSX1_1176 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_4564_), .Q(micro_hash_ucr_2_pipe71) );
INVX1 INVX1_573 ( .gnd(gnd), .vdd(vdd), .A(_0__bF_buf6), .Y(_12843_) );
NAND2X1 NAND2X1_1158 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf5), .B(_12843_), .Y(_12844_) );
NOR2X1 NOR2X1_1350 ( .gnd(gnd), .vdd(vdd), .A(comparador_next_bF_buf1), .B(_12844_), .Y(_8705_) );
NOR2X1 NOR2X1_1351 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe70_bF_buf3), .B(micro_hash_ucr_3_pipe5), .Y(_12845_) );
NAND2X1 NAND2X1_1159 ( .gnd(gnd), .vdd(vdd), .A(H_3_16_), .B(_12845_), .Y(_12846_) );
INVX2 INVX2_254 ( .gnd(gnd), .vdd(vdd), .A(H_3_16_), .Y(_12847_) );
INVX8 INVX8_194 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_0_), .Y(_12848_) );
OAI21X1 OAI21X1_2448 ( .gnd(gnd), .vdd(vdd), .A(_12847_), .B(_12848__bF_buf3), .C(micro_hash_ucr_3_pipe70_bF_buf2), .Y(_12849_) );
OAI21X1 OAI21X1_2449 ( .gnd(gnd), .vdd(vdd), .A(H_3_16_), .B(micro_hash_ucr_3_c_0_), .C(_8705__bF_buf13), .Y(_12850_) );
AOI21X1 AOI21X1_1524 ( .gnd(gnd), .vdd(vdd), .A(_12846_), .B(_12849_), .C(_12850_), .Y(_8703__16_) );
NOR2X1 NOR2X1_1352 ( .gnd(gnd), .vdd(vdd), .A(_12847_), .B(_12848__bF_buf2), .Y(_12851_) );
NOR2X1 NOR2X1_1353 ( .gnd(gnd), .vdd(vdd), .A(H_3_17_), .B(micro_hash_ucr_3_c_1_bF_buf3_), .Y(_12852_) );
NAND2X1 NAND2X1_1160 ( .gnd(gnd), .vdd(vdd), .A(H_3_17_), .B(micro_hash_ucr_3_c_1_bF_buf2_), .Y(_12853_) );
INVX1 INVX1_574 ( .gnd(gnd), .vdd(vdd), .A(_12853_), .Y(_12854_) );
NOR2X1 NOR2X1_1354 ( .gnd(gnd), .vdd(vdd), .A(_12852_), .B(_12854_), .Y(_12855_) );
XNOR2X1 XNOR2X1_375 ( .gnd(gnd), .vdd(vdd), .A(_12855_), .B(_12851_), .Y(_12856_) );
INVX8 INVX8_195 ( .gnd(gnd), .vdd(vdd), .A(_12845_), .Y(_12857_) );
OAI21X1 OAI21X1_2450 ( .gnd(gnd), .vdd(vdd), .A(H_3_17_), .B(_12857_), .C(_8705__bF_buf12), .Y(_12858_) );
AOI21X1 AOI21X1_1525 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe70_bF_buf1), .B(_12856_), .C(_12858_), .Y(_8703__17_) );
INVX1 INVX1_575 ( .gnd(gnd), .vdd(vdd), .A(_12851_), .Y(_12859_) );
OAI21X1 OAI21X1_2451 ( .gnd(gnd), .vdd(vdd), .A(_12859_), .B(_12852_), .C(_12853_), .Y(_12860_) );
XOR2X1 XOR2X1_154 ( .gnd(gnd), .vdd(vdd), .A(H_3_18_), .B(micro_hash_ucr_3_c_2_), .Y(_12861_) );
XNOR2X1 XNOR2X1_376 ( .gnd(gnd), .vdd(vdd), .A(_12860_), .B(_12861_), .Y(_12862_) );
OAI21X1 OAI21X1_2452 ( .gnd(gnd), .vdd(vdd), .A(H_3_18_), .B(_12857_), .C(_8705__bF_buf11), .Y(_12863_) );
AOI21X1 AOI21X1_1526 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe70_bF_buf0), .B(_12862_), .C(_12863_), .Y(_8703__18_) );
INVX1 INVX1_576 ( .gnd(gnd), .vdd(vdd), .A(_12860_), .Y(_12864_) );
INVX1 INVX1_577 ( .gnd(gnd), .vdd(vdd), .A(_12861_), .Y(_12865_) );
NOR2X1 NOR2X1_1355 ( .gnd(gnd), .vdd(vdd), .A(_12865_), .B(_12864_), .Y(_12866_) );
AOI21X1 AOI21X1_1527 ( .gnd(gnd), .vdd(vdd), .A(H_3_18_), .B(micro_hash_ucr_3_c_2_), .C(_12866_), .Y(_12867_) );
NOR2X1 NOR2X1_1356 ( .gnd(gnd), .vdd(vdd), .A(H_3_19_), .B(micro_hash_ucr_3_c_3_bF_buf3_), .Y(_12868_) );
INVX1 INVX1_578 ( .gnd(gnd), .vdd(vdd), .A(_12868_), .Y(_12869_) );
NAND2X1 NAND2X1_1161 ( .gnd(gnd), .vdd(vdd), .A(H_3_19_), .B(micro_hash_ucr_3_c_3_bF_buf2_), .Y(_12870_) );
NAND2X1 NAND2X1_1162 ( .gnd(gnd), .vdd(vdd), .A(_12870_), .B(_12869_), .Y(_12871_) );
XNOR2X1 XNOR2X1_377 ( .gnd(gnd), .vdd(vdd), .A(_12867_), .B(_12871_), .Y(_12872_) );
OAI21X1 OAI21X1_2453 ( .gnd(gnd), .vdd(vdd), .A(H_3_19_), .B(_12857_), .C(_8705__bF_buf10), .Y(_12873_) );
AOI21X1 AOI21X1_1528 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe70_bF_buf3), .B(_12872_), .C(_12873_), .Y(_8703__19_) );
NOR2X1 NOR2X1_1357 ( .gnd(gnd), .vdd(vdd), .A(H_3_20_), .B(micro_hash_ucr_3_c_4_), .Y(_12874_) );
AND2X2 AND2X2_511 ( .gnd(gnd), .vdd(vdd), .A(H_3_20_), .B(micro_hash_ucr_3_c_4_), .Y(_12875_) );
NOR2X1 NOR2X1_1358 ( .gnd(gnd), .vdd(vdd), .A(_12874_), .B(_12875_), .Y(_12876_) );
OAI21X1 OAI21X1_2454 ( .gnd(gnd), .vdd(vdd), .A(_12867_), .B(_12868_), .C(_12870_), .Y(_12877_) );
XNOR2X1 XNOR2X1_378 ( .gnd(gnd), .vdd(vdd), .A(_12877_), .B(_12876_), .Y(_12878_) );
OAI21X1 OAI21X1_2455 ( .gnd(gnd), .vdd(vdd), .A(H_3_20_), .B(_12857_), .C(_8705__bF_buf9), .Y(_12879_) );
AOI21X1 AOI21X1_1529 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe70_bF_buf2), .B(_12878_), .C(_12879_), .Y(_8703__20_) );
AOI21X1 AOI21X1_1530 ( .gnd(gnd), .vdd(vdd), .A(_12876_), .B(_12877_), .C(_12875_), .Y(_12880_) );
NOR2X1 NOR2X1_1359 ( .gnd(gnd), .vdd(vdd), .A(H_3_21_), .B(micro_hash_ucr_3_c_5_), .Y(_12881_) );
NAND2X1 NAND2X1_1163 ( .gnd(gnd), .vdd(vdd), .A(H_3_21_), .B(micro_hash_ucr_3_c_5_), .Y(_12882_) );
INVX1 INVX1_579 ( .gnd(gnd), .vdd(vdd), .A(_12882_), .Y(_12883_) );
NOR2X1 NOR2X1_1360 ( .gnd(gnd), .vdd(vdd), .A(_12881_), .B(_12883_), .Y(_12884_) );
OAI21X1 OAI21X1_2456 ( .gnd(gnd), .vdd(vdd), .A(_12880_), .B(_12884_), .C(micro_hash_ucr_3_pipe70_bF_buf1), .Y(_12885_) );
AOI21X1 AOI21X1_1531 ( .gnd(gnd), .vdd(vdd), .A(_12880_), .B(_12884_), .C(_12885_), .Y(_12886_) );
OAI21X1 OAI21X1_2457 ( .gnd(gnd), .vdd(vdd), .A(H_3_21_), .B(_12857_), .C(_8705__bF_buf8), .Y(_12887_) );
NOR2X1 NOR2X1_1361 ( .gnd(gnd), .vdd(vdd), .A(_12887_), .B(_12886_), .Y(_8703__21_) );
XOR2X1 XOR2X1_155 ( .gnd(gnd), .vdd(vdd), .A(H_3_22_), .B(micro_hash_ucr_3_c_6_), .Y(_12888_) );
OAI21X1 OAI21X1_2458 ( .gnd(gnd), .vdd(vdd), .A(_12880_), .B(_12881_), .C(_12882_), .Y(_12889_) );
XNOR2X1 XNOR2X1_379 ( .gnd(gnd), .vdd(vdd), .A(_12889_), .B(_12888_), .Y(_12890_) );
OAI21X1 OAI21X1_2459 ( .gnd(gnd), .vdd(vdd), .A(H_3_22_), .B(_12857_), .C(_8705__bF_buf7), .Y(_12891_) );
AOI21X1 AOI21X1_1532 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe70_bF_buf0), .B(_12890_), .C(_12891_), .Y(_8703__22_) );
INVX1 INVX1_580 ( .gnd(gnd), .vdd(vdd), .A(H_3_22_), .Y(_12892_) );
INVX2 INVX2_255 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_6_), .Y(_12893_) );
NAND2X1 NAND2X1_1164 ( .gnd(gnd), .vdd(vdd), .A(_12888_), .B(_12889_), .Y(_12894_) );
OAI21X1 OAI21X1_2460 ( .gnd(gnd), .vdd(vdd), .A(_12892_), .B(_12893_), .C(_12894_), .Y(_12895_) );
XOR2X1 XOR2X1_156 ( .gnd(gnd), .vdd(vdd), .A(H_3_23_), .B(micro_hash_ucr_3_c_7_), .Y(_12896_) );
XNOR2X1 XNOR2X1_380 ( .gnd(gnd), .vdd(vdd), .A(_12895_), .B(_12896_), .Y(_12897_) );
OAI21X1 OAI21X1_2461 ( .gnd(gnd), .vdd(vdd), .A(H_3_23_), .B(_12857_), .C(_8705__bF_buf6), .Y(_12898_) );
AOI21X1 AOI21X1_1533 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe70_bF_buf3), .B(_12897_), .C(_12898_), .Y(_8703__23_) );
INVX2 INVX2_256 ( .gnd(gnd), .vdd(vdd), .A(H_3_8_), .Y(_12899_) );
INVX8 INVX8_196 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe70_bF_buf2), .Y(_12900_) );
OAI21X1 OAI21X1_2462 ( .gnd(gnd), .vdd(vdd), .A(_12900__bF_buf3), .B(micro_hash_ucr_3_b_0_bF_buf3_), .C(_12857_), .Y(_12901_) );
INVX8 INVX8_197 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_0_bF_buf2_), .Y(_12902_) );
NOR2X1 NOR2X1_1362 ( .gnd(gnd), .vdd(vdd), .A(_12899_), .B(_12902_), .Y(_12903_) );
INVX1 INVX1_581 ( .gnd(gnd), .vdd(vdd), .A(_12903_), .Y(_12904_) );
OAI21X1 OAI21X1_2463 ( .gnd(gnd), .vdd(vdd), .A(_12904_), .B(_12900__bF_buf2), .C(_8705__bF_buf5), .Y(_12905_) );
AOI21X1 AOI21X1_1534 ( .gnd(gnd), .vdd(vdd), .A(_12899_), .B(_12901_), .C(_12905_), .Y(_8703__8_) );
INVX2 INVX2_257 ( .gnd(gnd), .vdd(vdd), .A(H_3_9_), .Y(_12906_) );
NOR2X1 NOR2X1_1363 ( .gnd(gnd), .vdd(vdd), .A(H_3_9_), .B(micro_hash_ucr_3_b_1_bF_buf3_), .Y(_12907_) );
INVX8 INVX8_198 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_1_bF_buf2_), .Y(_12908_) );
NOR2X1 NOR2X1_1364 ( .gnd(gnd), .vdd(vdd), .A(_12906_), .B(_12908__bF_buf3), .Y(_12909_) );
NOR2X1 NOR2X1_1365 ( .gnd(gnd), .vdd(vdd), .A(_12907_), .B(_12909_), .Y(_12910_) );
AOI21X1 AOI21X1_1535 ( .gnd(gnd), .vdd(vdd), .A(_12903_), .B(_12910_), .C(_12900__bF_buf1), .Y(_12911_) );
OAI21X1 OAI21X1_2464 ( .gnd(gnd), .vdd(vdd), .A(_12903_), .B(_12910_), .C(_12911_), .Y(_12912_) );
OAI21X1 OAI21X1_2465 ( .gnd(gnd), .vdd(vdd), .A(_12906_), .B(_12857_), .C(_12912_), .Y(_12913_) );
AND2X2 AND2X2_512 ( .gnd(gnd), .vdd(vdd), .A(_12913_), .B(_8705__bF_buf4), .Y(_8703__9_) );
INVX2 INVX2_258 ( .gnd(gnd), .vdd(vdd), .A(H_3_10_), .Y(_8779_) );
INVX1 INVX1_582 ( .gnd(gnd), .vdd(vdd), .A(_12909_), .Y(_8780_) );
OAI21X1 OAI21X1_2466 ( .gnd(gnd), .vdd(vdd), .A(_12904_), .B(_12907_), .C(_8780_), .Y(_8781_) );
XOR2X1 XOR2X1_157 ( .gnd(gnd), .vdd(vdd), .A(H_3_10_), .B(micro_hash_ucr_3_b_2_bF_buf3_), .Y(_8782_) );
INVX1 INVX1_583 ( .gnd(gnd), .vdd(vdd), .A(_8781_), .Y(_8783_) );
INVX1 INVX1_584 ( .gnd(gnd), .vdd(vdd), .A(_8782_), .Y(_8784_) );
NOR2X1 NOR2X1_1366 ( .gnd(gnd), .vdd(vdd), .A(_8784_), .B(_8783_), .Y(_8785_) );
NOR2X1 NOR2X1_1367 ( .gnd(gnd), .vdd(vdd), .A(_12900__bF_buf0), .B(_8785_), .Y(_8786_) );
OAI21X1 OAI21X1_2467 ( .gnd(gnd), .vdd(vdd), .A(_8781_), .B(_8782_), .C(_8786_), .Y(_8787_) );
OAI21X1 OAI21X1_2468 ( .gnd(gnd), .vdd(vdd), .A(_8779_), .B(_12857_), .C(_8787_), .Y(_8788_) );
AND2X2 AND2X2_513 ( .gnd(gnd), .vdd(vdd), .A(_8788_), .B(_8705__bF_buf3), .Y(_8703__10_) );
INVX8 INVX8_199 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_2_bF_buf2_), .Y(_8789_) );
INVX1 INVX1_585 ( .gnd(gnd), .vdd(vdd), .A(_8785_), .Y(_8790_) );
OAI21X1 OAI21X1_2469 ( .gnd(gnd), .vdd(vdd), .A(_8779_), .B(_8789__bF_buf3), .C(_8790_), .Y(_8791_) );
NOR2X1 NOR2X1_1368 ( .gnd(gnd), .vdd(vdd), .A(H_3_11_), .B(micro_hash_ucr_3_b_3_bF_buf3_), .Y(_8792_) );
INVX1 INVX1_586 ( .gnd(gnd), .vdd(vdd), .A(H_3_11_), .Y(_8793_) );
INVX8 INVX8_200 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_3_bF_buf2_), .Y(_8794_) );
NOR2X1 NOR2X1_1369 ( .gnd(gnd), .vdd(vdd), .A(_8793_), .B(_8794_), .Y(_8795_) );
OR2X2 OR2X2_65 ( .gnd(gnd), .vdd(vdd), .A(_8795_), .B(_8792_), .Y(_8796_) );
OAI21X1 OAI21X1_2470 ( .gnd(gnd), .vdd(vdd), .A(_8791_), .B(_8796_), .C(micro_hash_ucr_3_pipe70_bF_buf1), .Y(_8797_) );
AOI21X1 AOI21X1_1536 ( .gnd(gnd), .vdd(vdd), .A(_8791_), .B(_8796_), .C(_8797_), .Y(_8798_) );
OAI21X1 OAI21X1_2471 ( .gnd(gnd), .vdd(vdd), .A(H_3_11_), .B(_12857_), .C(_8705__bF_buf2), .Y(_8799_) );
NOR2X1 NOR2X1_1370 ( .gnd(gnd), .vdd(vdd), .A(_8799_), .B(_8798_), .Y(_8703__11_) );
INVX8 INVX8_201 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf1), .Y(_8800_) );
XOR2X1 XOR2X1_158 ( .gnd(gnd), .vdd(vdd), .A(H_3_12_), .B(micro_hash_ucr_3_b_4_bF_buf4_), .Y(_8801_) );
INVX1 INVX1_587 ( .gnd(gnd), .vdd(vdd), .A(_8792_), .Y(_8802_) );
AOI21X1 AOI21X1_1537 ( .gnd(gnd), .vdd(vdd), .A(_8802_), .B(_8791_), .C(_8795_), .Y(_8803_) );
XNOR2X1 XNOR2X1_381 ( .gnd(gnd), .vdd(vdd), .A(_8803_), .B(_8801_), .Y(_8804_) );
INVX1 INVX1_588 ( .gnd(gnd), .vdd(vdd), .A(H_3_12_), .Y(_8805_) );
OAI21X1 OAI21X1_2472 ( .gnd(gnd), .vdd(vdd), .A(_8805_), .B(micro_hash_ucr_3_pipe5), .C(_12900__bF_buf3), .Y(_8806_) );
OAI21X1 OAI21X1_2473 ( .gnd(gnd), .vdd(vdd), .A(_8804_), .B(_12900__bF_buf2), .C(_8806_), .Y(_8807_) );
NOR2X1 NOR2X1_1371 ( .gnd(gnd), .vdd(vdd), .A(_8800__bF_buf12), .B(_8807_), .Y(_8703__12_) );
NAND2X1 NAND2X1_1165 ( .gnd(gnd), .vdd(vdd), .A(H_3_12_), .B(micro_hash_ucr_3_b_4_bF_buf3_), .Y(_8808_) );
INVX1 INVX1_589 ( .gnd(gnd), .vdd(vdd), .A(_8801_), .Y(_8809_) );
OAI21X1 OAI21X1_2474 ( .gnd(gnd), .vdd(vdd), .A(_8803_), .B(_8809_), .C(_8808_), .Y(_8810_) );
INVX2 INVX2_259 ( .gnd(gnd), .vdd(vdd), .A(_8810_), .Y(_8811_) );
NOR2X1 NOR2X1_1372 ( .gnd(gnd), .vdd(vdd), .A(H_3_13_), .B(micro_hash_ucr_3_b_5_bF_buf3_), .Y(_8812_) );
INVX1 INVX1_590 ( .gnd(gnd), .vdd(vdd), .A(H_3_13_), .Y(_8813_) );
INVX8 INVX8_202 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_5_bF_buf2_), .Y(_8814_) );
NOR2X1 NOR2X1_1373 ( .gnd(gnd), .vdd(vdd), .A(_8813_), .B(_8814__bF_buf3), .Y(_8815_) );
NOR2X1 NOR2X1_1374 ( .gnd(gnd), .vdd(vdd), .A(_8812_), .B(_8815_), .Y(_8816_) );
AND2X2 AND2X2_514 ( .gnd(gnd), .vdd(vdd), .A(_8811_), .B(_8816_), .Y(_8817_) );
OAI21X1 OAI21X1_2475 ( .gnd(gnd), .vdd(vdd), .A(_8811_), .B(_8816_), .C(micro_hash_ucr_3_pipe70_bF_buf0), .Y(_8818_) );
OAI21X1 OAI21X1_2476 ( .gnd(gnd), .vdd(vdd), .A(_8813_), .B(micro_hash_ucr_3_pipe5), .C(_12900__bF_buf1), .Y(_8819_) );
OAI21X1 OAI21X1_2477 ( .gnd(gnd), .vdd(vdd), .A(_8817_), .B(_8818_), .C(_8819_), .Y(_8820_) );
NOR2X1 NOR2X1_1375 ( .gnd(gnd), .vdd(vdd), .A(_8800__bF_buf11), .B(_8820_), .Y(_8703__13_) );
XOR2X1 XOR2X1_159 ( .gnd(gnd), .vdd(vdd), .A(H_3_14_), .B(micro_hash_ucr_3_b_6_bF_buf3_), .Y(_8821_) );
INVX1 INVX1_591 ( .gnd(gnd), .vdd(vdd), .A(_8815_), .Y(_8822_) );
OAI21X1 OAI21X1_2478 ( .gnd(gnd), .vdd(vdd), .A(_8811_), .B(_8812_), .C(_8822_), .Y(_8823_) );
XNOR2X1 XNOR2X1_382 ( .gnd(gnd), .vdd(vdd), .A(_8823_), .B(_8821_), .Y(_8824_) );
INVX1 INVX1_592 ( .gnd(gnd), .vdd(vdd), .A(H_3_14_), .Y(_8825_) );
OAI21X1 OAI21X1_2479 ( .gnd(gnd), .vdd(vdd), .A(_8825_), .B(micro_hash_ucr_3_pipe5), .C(_12900__bF_buf0), .Y(_8826_) );
NAND2X1 NAND2X1_1166 ( .gnd(gnd), .vdd(vdd), .A(_8826_), .B(_8705__bF_buf0), .Y(_8827_) );
AOI21X1 AOI21X1_1538 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe70_bF_buf3), .B(_8824_), .C(_8827_), .Y(_8703__14_) );
INVX8 INVX8_203 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_6_bF_buf2_), .Y(_8828_) );
NAND2X1 NAND2X1_1167 ( .gnd(gnd), .vdd(vdd), .A(_8821_), .B(_8823_), .Y(_8829_) );
OAI21X1 OAI21X1_2480 ( .gnd(gnd), .vdd(vdd), .A(_8825_), .B(_8828_), .C(_8829_), .Y(_8830_) );
XOR2X1 XOR2X1_160 ( .gnd(gnd), .vdd(vdd), .A(H_3_15_), .B(micro_hash_ucr_3_b_7_bF_buf3_), .Y(_8831_) );
XNOR2X1 XNOR2X1_383 ( .gnd(gnd), .vdd(vdd), .A(_8830_), .B(_8831_), .Y(_8832_) );
OAI21X1 OAI21X1_2481 ( .gnd(gnd), .vdd(vdd), .A(H_3_15_), .B(_12857_), .C(_8705__bF_buf13), .Y(_8833_) );
AOI21X1 AOI21X1_1539 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe70_bF_buf2), .B(_8832_), .C(_8833_), .Y(_8703__15_) );
INVX1 INVX1_593 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_216_), .Y(_8834_) );
XNOR2X1 XNOR2X1_384 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_168_), .B(micro_hash_ucr_3_Wx_128_), .Y(_8835_) );
AOI21X1 AOI21X1_1540 ( .gnd(gnd), .vdd(vdd), .A(_8834_), .B(_8835_), .C(_8800__bF_buf10), .Y(_8699__240_) );
INVX2 INVX2_260 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_169_), .Y(_8836_) );
INVX1 INVX1_594 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_217_), .Y(_8837_) );
OAI21X1 OAI21X1_2482 ( .gnd(gnd), .vdd(vdd), .A(_8836_), .B(micro_hash_ucr_3_Wx_129_), .C(_8837_), .Y(_8838_) );
AOI21X1 AOI21X1_1541 ( .gnd(gnd), .vdd(vdd), .A(_8836_), .B(micro_hash_ucr_3_Wx_129_), .C(_8838_), .Y(_8839_) );
NOR2X1 NOR2X1_1376 ( .gnd(gnd), .vdd(vdd), .A(_8839_), .B(_8800__bF_buf9), .Y(_8699__241_) );
INVX4 INVX4_108 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_170_), .Y(_8840_) );
INVX2 INVX2_261 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_218_), .Y(_8841_) );
OAI21X1 OAI21X1_2483 ( .gnd(gnd), .vdd(vdd), .A(_8840_), .B(micro_hash_ucr_3_Wx_130_), .C(_8841_), .Y(_8842_) );
AOI21X1 AOI21X1_1542 ( .gnd(gnd), .vdd(vdd), .A(_8840_), .B(micro_hash_ucr_3_Wx_130_), .C(_8842_), .Y(_8843_) );
NOR2X1 NOR2X1_1377 ( .gnd(gnd), .vdd(vdd), .A(_8843_), .B(_8800__bF_buf8), .Y(_8699__242_) );
INVX2 INVX2_262 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_171_), .Y(_8844_) );
INVX1 INVX1_595 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_219_), .Y(_8845_) );
OAI21X1 OAI21X1_2484 ( .gnd(gnd), .vdd(vdd), .A(_8844_), .B(micro_hash_ucr_3_Wx_131_), .C(_8845_), .Y(_8846_) );
AOI21X1 AOI21X1_1543 ( .gnd(gnd), .vdd(vdd), .A(_8844_), .B(micro_hash_ucr_3_Wx_131_), .C(_8846_), .Y(_8847_) );
NOR2X1 NOR2X1_1378 ( .gnd(gnd), .vdd(vdd), .A(_8847_), .B(_8800__bF_buf7), .Y(_8699__243_) );
INVX2 INVX2_263 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_172_), .Y(_8848_) );
AOI21X1 AOI21X1_1544 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_132_), .B(_8848_), .C(micro_hash_ucr_3_Wx_220_), .Y(_8849_) );
OAI21X1 OAI21X1_2485 ( .gnd(gnd), .vdd(vdd), .A(_8848_), .B(micro_hash_ucr_3_Wx_132_), .C(_8849_), .Y(_8850_) );
AND2X2 AND2X2_515 ( .gnd(gnd), .vdd(vdd), .A(_8850_), .B(_8705__bF_buf12), .Y(_8699__244_) );
INVX2 INVX2_264 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_173_), .Y(_8851_) );
AOI21X1 AOI21X1_1545 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_133_), .B(_8851_), .C(micro_hash_ucr_3_Wx_221_), .Y(_8852_) );
OAI21X1 OAI21X1_2486 ( .gnd(gnd), .vdd(vdd), .A(_8851_), .B(micro_hash_ucr_3_Wx_133_), .C(_8852_), .Y(_8853_) );
AND2X2 AND2X2_516 ( .gnd(gnd), .vdd(vdd), .A(_8853_), .B(_8705__bF_buf11), .Y(_8699__245_) );
INVX4 INVX4_109 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_174_), .Y(_8854_) );
INVX2 INVX2_265 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_222_), .Y(_8855_) );
OAI21X1 OAI21X1_2487 ( .gnd(gnd), .vdd(vdd), .A(_8854_), .B(micro_hash_ucr_3_Wx_134_), .C(_8855_), .Y(_8856_) );
AOI21X1 AOI21X1_1546 ( .gnd(gnd), .vdd(vdd), .A(_8854_), .B(micro_hash_ucr_3_Wx_134_), .C(_8856_), .Y(_8857_) );
NOR2X1 NOR2X1_1379 ( .gnd(gnd), .vdd(vdd), .A(_8857_), .B(_8800__bF_buf6), .Y(_8699__246_) );
INVX1 INVX1_596 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_223_), .Y(_8858_) );
XNOR2X1 XNOR2X1_385 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_175_), .B(micro_hash_ucr_3_Wx_135_), .Y(_8859_) );
AOI21X1 AOI21X1_1547 ( .gnd(gnd), .vdd(vdd), .A(_8858_), .B(_8859_), .C(_8800__bF_buf5), .Y(_8699__247_) );
INVX1 INVX1_597 ( .gnd(gnd), .vdd(vdd), .A(H_3_0_), .Y(_8860_) );
OAI21X1 OAI21X1_2488 ( .gnd(gnd), .vdd(vdd), .A(_12900__bF_buf3), .B(micro_hash_ucr_3_a_0_bF_buf3_), .C(_12857_), .Y(_8861_) );
INVX8 INVX8_204 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_0_bF_buf2_), .Y(_8862_) );
NOR2X1 NOR2X1_1380 ( .gnd(gnd), .vdd(vdd), .A(_8860_), .B(_8862__bF_buf3), .Y(_8863_) );
INVX1 INVX1_598 ( .gnd(gnd), .vdd(vdd), .A(_8863_), .Y(_8864_) );
OAI21X1 OAI21X1_2489 ( .gnd(gnd), .vdd(vdd), .A(_8864_), .B(_12900__bF_buf2), .C(_8705__bF_buf10), .Y(_8865_) );
AOI21X1 AOI21X1_1548 ( .gnd(gnd), .vdd(vdd), .A(_8860_), .B(_8861_), .C(_8865_), .Y(_8703__0_) );
INVX2 INVX2_266 ( .gnd(gnd), .vdd(vdd), .A(H_3_1_), .Y(_8866_) );
NOR2X1 NOR2X1_1381 ( .gnd(gnd), .vdd(vdd), .A(H_3_1_), .B(micro_hash_ucr_3_a_1_bF_buf3_), .Y(_8867_) );
INVX8 INVX8_205 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_1_bF_buf2_), .Y(_8868_) );
NOR2X1 NOR2X1_1382 ( .gnd(gnd), .vdd(vdd), .A(_8866_), .B(_8868__bF_buf3), .Y(_8869_) );
NOR2X1 NOR2X1_1383 ( .gnd(gnd), .vdd(vdd), .A(_8867_), .B(_8869_), .Y(_8870_) );
AOI21X1 AOI21X1_1549 ( .gnd(gnd), .vdd(vdd), .A(_8863_), .B(_8870_), .C(_12900__bF_buf1), .Y(_8871_) );
OAI21X1 OAI21X1_2490 ( .gnd(gnd), .vdd(vdd), .A(_8863_), .B(_8870_), .C(_8871_), .Y(_8872_) );
OAI21X1 OAI21X1_2491 ( .gnd(gnd), .vdd(vdd), .A(_8866_), .B(_12857_), .C(_8872_), .Y(_8873_) );
AND2X2 AND2X2_517 ( .gnd(gnd), .vdd(vdd), .A(_8873_), .B(_8705__bF_buf9), .Y(_8703__1_) );
INVX2 INVX2_267 ( .gnd(gnd), .vdd(vdd), .A(H_3_2_), .Y(_8874_) );
INVX1 INVX1_599 ( .gnd(gnd), .vdd(vdd), .A(_8869_), .Y(_8875_) );
OAI21X1 OAI21X1_2492 ( .gnd(gnd), .vdd(vdd), .A(_8864_), .B(_8867_), .C(_8875_), .Y(_8876_) );
XOR2X1 XOR2X1_161 ( .gnd(gnd), .vdd(vdd), .A(H_3_2_), .B(micro_hash_ucr_3_a_2_), .Y(_8877_) );
INVX1 INVX1_600 ( .gnd(gnd), .vdd(vdd), .A(_8876_), .Y(_8878_) );
INVX1 INVX1_601 ( .gnd(gnd), .vdd(vdd), .A(_8877_), .Y(_8879_) );
NOR2X1 NOR2X1_1384 ( .gnd(gnd), .vdd(vdd), .A(_8879_), .B(_8878_), .Y(_8880_) );
NOR2X1 NOR2X1_1385 ( .gnd(gnd), .vdd(vdd), .A(_12900__bF_buf0), .B(_8880_), .Y(_8881_) );
OAI21X1 OAI21X1_2493 ( .gnd(gnd), .vdd(vdd), .A(_8876_), .B(_8877_), .C(_8881_), .Y(_8882_) );
OAI21X1 OAI21X1_2494 ( .gnd(gnd), .vdd(vdd), .A(_8874_), .B(_12857_), .C(_8882_), .Y(_8883_) );
AND2X2 AND2X2_518 ( .gnd(gnd), .vdd(vdd), .A(_8883_), .B(_8705__bF_buf8), .Y(_8703__2_) );
INVX8 INVX8_206 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_2_), .Y(_8884_) );
INVX1 INVX1_602 ( .gnd(gnd), .vdd(vdd), .A(_8880_), .Y(_8885_) );
OAI21X1 OAI21X1_2495 ( .gnd(gnd), .vdd(vdd), .A(_8874_), .B(_8884_), .C(_8885_), .Y(_8886_) );
NOR2X1 NOR2X1_1386 ( .gnd(gnd), .vdd(vdd), .A(H_3_3_), .B(micro_hash_ucr_3_a_3_), .Y(_8887_) );
INVX1 INVX1_603 ( .gnd(gnd), .vdd(vdd), .A(_8887_), .Y(_8888_) );
NAND2X1 NAND2X1_1168 ( .gnd(gnd), .vdd(vdd), .A(H_3_3_), .B(micro_hash_ucr_3_a_3_), .Y(_8889_) );
NAND2X1 NAND2X1_1169 ( .gnd(gnd), .vdd(vdd), .A(_8889_), .B(_8888_), .Y(_8890_) );
AND2X2 AND2X2_519 ( .gnd(gnd), .vdd(vdd), .A(_8886_), .B(_8890_), .Y(_8891_) );
OAI21X1 OAI21X1_2496 ( .gnd(gnd), .vdd(vdd), .A(_8886_), .B(_8890_), .C(micro_hash_ucr_3_pipe70_bF_buf1), .Y(_8892_) );
INVX1 INVX1_604 ( .gnd(gnd), .vdd(vdd), .A(H_3_3_), .Y(_8893_) );
OAI21X1 OAI21X1_2497 ( .gnd(gnd), .vdd(vdd), .A(_8893_), .B(micro_hash_ucr_3_pipe5), .C(_12900__bF_buf3), .Y(_8894_) );
OAI21X1 OAI21X1_2498 ( .gnd(gnd), .vdd(vdd), .A(_8891_), .B(_8892_), .C(_8894_), .Y(_8895_) );
NOR2X1 NOR2X1_1387 ( .gnd(gnd), .vdd(vdd), .A(_8800__bF_buf4), .B(_8895_), .Y(_8703__3_) );
XOR2X1 XOR2X1_162 ( .gnd(gnd), .vdd(vdd), .A(H_3_4_), .B(micro_hash_ucr_3_a_4_), .Y(_8896_) );
INVX1 INVX1_605 ( .gnd(gnd), .vdd(vdd), .A(_8886_), .Y(_8897_) );
OAI21X1 OAI21X1_2499 ( .gnd(gnd), .vdd(vdd), .A(_8897_), .B(_8887_), .C(_8889_), .Y(_8898_) );
XNOR2X1 XNOR2X1_386 ( .gnd(gnd), .vdd(vdd), .A(_8898_), .B(_8896_), .Y(_8899_) );
INVX1 INVX1_606 ( .gnd(gnd), .vdd(vdd), .A(H_3_4_), .Y(_8900_) );
OAI21X1 OAI21X1_2500 ( .gnd(gnd), .vdd(vdd), .A(_8900_), .B(micro_hash_ucr_3_pipe5), .C(_12900__bF_buf2), .Y(_8901_) );
NAND2X1 NAND2X1_1170 ( .gnd(gnd), .vdd(vdd), .A(_8901_), .B(_8705__bF_buf7), .Y(_8902_) );
AOI21X1 AOI21X1_1550 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe70_bF_buf0), .B(_8899_), .C(_8902_), .Y(_8703__4_) );
INVX8 INVX8_207 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_4_), .Y(_8903_) );
NAND2X1 NAND2X1_1171 ( .gnd(gnd), .vdd(vdd), .A(_8896_), .B(_8898_), .Y(_8904_) );
OAI21X1 OAI21X1_2501 ( .gnd(gnd), .vdd(vdd), .A(_8900_), .B(_8903__bF_buf3), .C(_8904_), .Y(_8905_) );
INVX2 INVX2_268 ( .gnd(gnd), .vdd(vdd), .A(_8905_), .Y(_8906_) );
NOR2X1 NOR2X1_1388 ( .gnd(gnd), .vdd(vdd), .A(H_3_5_), .B(micro_hash_ucr_3_a_5_bF_buf3_), .Y(_8907_) );
INVX1 INVX1_607 ( .gnd(gnd), .vdd(vdd), .A(H_3_5_), .Y(_8908_) );
INVX8 INVX8_208 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_5_bF_buf2_), .Y(_8909_) );
NOR2X1 NOR2X1_1389 ( .gnd(gnd), .vdd(vdd), .A(_8908_), .B(_8909_), .Y(_8910_) );
NOR2X1 NOR2X1_1390 ( .gnd(gnd), .vdd(vdd), .A(_8907_), .B(_8910_), .Y(_8911_) );
AND2X2 AND2X2_520 ( .gnd(gnd), .vdd(vdd), .A(_8906_), .B(_8911_), .Y(_8912_) );
OAI21X1 OAI21X1_2502 ( .gnd(gnd), .vdd(vdd), .A(_8906_), .B(_8911_), .C(micro_hash_ucr_3_pipe70_bF_buf3), .Y(_8913_) );
OAI21X1 OAI21X1_2503 ( .gnd(gnd), .vdd(vdd), .A(_8908_), .B(micro_hash_ucr_3_pipe5), .C(_12900__bF_buf1), .Y(_8914_) );
OAI21X1 OAI21X1_2504 ( .gnd(gnd), .vdd(vdd), .A(_8912_), .B(_8913_), .C(_8914_), .Y(_8915_) );
NOR2X1 NOR2X1_1391 ( .gnd(gnd), .vdd(vdd), .A(_8800__bF_buf3), .B(_8915_), .Y(_8703__5_) );
XOR2X1 XOR2X1_163 ( .gnd(gnd), .vdd(vdd), .A(H_3_6_), .B(micro_hash_ucr_3_a_6_bF_buf3_), .Y(_8916_) );
INVX1 INVX1_608 ( .gnd(gnd), .vdd(vdd), .A(_8910_), .Y(_8917_) );
OAI21X1 OAI21X1_2505 ( .gnd(gnd), .vdd(vdd), .A(_8906_), .B(_8907_), .C(_8917_), .Y(_8918_) );
XOR2X1 XOR2X1_164 ( .gnd(gnd), .vdd(vdd), .A(_8918_), .B(_8916_), .Y(_8919_) );
INVX2 INVX2_269 ( .gnd(gnd), .vdd(vdd), .A(H_3_6_), .Y(_8920_) );
OAI21X1 OAI21X1_2506 ( .gnd(gnd), .vdd(vdd), .A(_8920_), .B(micro_hash_ucr_3_pipe5), .C(_12900__bF_buf0), .Y(_8921_) );
OAI21X1 OAI21X1_2507 ( .gnd(gnd), .vdd(vdd), .A(_8919_), .B(_12900__bF_buf3), .C(_8921_), .Y(_8922_) );
NOR2X1 NOR2X1_1392 ( .gnd(gnd), .vdd(vdd), .A(_8800__bF_buf2), .B(_8922_), .Y(_8703__6_) );
INVX8 INVX8_209 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_6_bF_buf2_), .Y(_8923_) );
NAND2X1 NAND2X1_1172 ( .gnd(gnd), .vdd(vdd), .A(_8916_), .B(_8918_), .Y(_8924_) );
OAI21X1 OAI21X1_2508 ( .gnd(gnd), .vdd(vdd), .A(_8920_), .B(_8923_), .C(_8924_), .Y(_8925_) );
XNOR2X1 XNOR2X1_387 ( .gnd(gnd), .vdd(vdd), .A(H_3_7_), .B(micro_hash_ucr_3_a_7_bF_buf3_), .Y(_8926_) );
AND2X2 AND2X2_521 ( .gnd(gnd), .vdd(vdd), .A(_8925_), .B(_8926_), .Y(_8927_) );
OAI21X1 OAI21X1_2509 ( .gnd(gnd), .vdd(vdd), .A(_8925_), .B(_8926_), .C(micro_hash_ucr_3_pipe70_bF_buf2), .Y(_8928_) );
INVX1 INVX1_609 ( .gnd(gnd), .vdd(vdd), .A(H_3_7_), .Y(_8929_) );
OAI21X1 OAI21X1_2510 ( .gnd(gnd), .vdd(vdd), .A(_8929_), .B(micro_hash_ucr_3_pipe5), .C(_12900__bF_buf2), .Y(_8930_) );
OAI21X1 OAI21X1_2511 ( .gnd(gnd), .vdd(vdd), .A(_8927_), .B(_8928_), .C(_8930_), .Y(_8931_) );
NOR2X1 NOR2X1_1393 ( .gnd(gnd), .vdd(vdd), .A(_8800__bF_buf1), .B(_8931_), .Y(_8703__7_) );
INVX2 INVX2_270 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_144_), .Y(_8932_) );
INVX1 INVX1_610 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_192_), .Y(_8933_) );
OAI21X1 OAI21X1_2512 ( .gnd(gnd), .vdd(vdd), .A(_8932_), .B(micro_hash_ucr_3_Wx_104_), .C(_8933_), .Y(_8934_) );
AOI21X1 AOI21X1_1551 ( .gnd(gnd), .vdd(vdd), .A(_8932_), .B(micro_hash_ucr_3_Wx_104_), .C(_8934_), .Y(_8935_) );
NOR2X1 NOR2X1_1394 ( .gnd(gnd), .vdd(vdd), .A(_8935_), .B(_8800__bF_buf0), .Y(_8699__216_) );
INVX2 INVX2_271 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_145_), .Y(_8936_) );
INVX2 INVX2_272 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_193_), .Y(_8937_) );
OAI21X1 OAI21X1_2513 ( .gnd(gnd), .vdd(vdd), .A(_8936_), .B(micro_hash_ucr_3_Wx_105_), .C(_8937_), .Y(_8938_) );
AOI21X1 AOI21X1_1552 ( .gnd(gnd), .vdd(vdd), .A(_8936_), .B(micro_hash_ucr_3_Wx_105_), .C(_8938_), .Y(_8939_) );
NOR2X1 NOR2X1_1395 ( .gnd(gnd), .vdd(vdd), .A(_8939_), .B(_8800__bF_buf12), .Y(_8699__217_) );
INVX4 INVX4_110 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_146_), .Y(_8940_) );
INVX2 INVX2_273 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_194_), .Y(_8941_) );
OAI21X1 OAI21X1_2514 ( .gnd(gnd), .vdd(vdd), .A(_8940_), .B(micro_hash_ucr_3_Wx_106_), .C(_8941_), .Y(_8942_) );
AOI21X1 AOI21X1_1553 ( .gnd(gnd), .vdd(vdd), .A(_8940_), .B(micro_hash_ucr_3_Wx_106_), .C(_8942_), .Y(_8943_) );
NOR2X1 NOR2X1_1396 ( .gnd(gnd), .vdd(vdd), .A(_8943_), .B(_8800__bF_buf11), .Y(_8699__218_) );
INVX2 INVX2_274 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_147_), .Y(_8944_) );
INVX1 INVX1_611 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_195_), .Y(_8945_) );
OAI21X1 OAI21X1_2515 ( .gnd(gnd), .vdd(vdd), .A(_8944_), .B(micro_hash_ucr_3_Wx_107_), .C(_8945_), .Y(_8946_) );
AOI21X1 AOI21X1_1554 ( .gnd(gnd), .vdd(vdd), .A(_8944_), .B(micro_hash_ucr_3_Wx_107_), .C(_8946_), .Y(_8947_) );
NOR2X1 NOR2X1_1397 ( .gnd(gnd), .vdd(vdd), .A(_8947_), .B(_8800__bF_buf10), .Y(_8699__219_) );
INVX2 INVX2_275 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_148_), .Y(_8948_) );
AOI21X1 AOI21X1_1555 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_108_), .B(_8948_), .C(micro_hash_ucr_3_Wx_196_), .Y(_8949_) );
OAI21X1 OAI21X1_2516 ( .gnd(gnd), .vdd(vdd), .A(_8948_), .B(micro_hash_ucr_3_Wx_108_), .C(_8949_), .Y(_8950_) );
AND2X2 AND2X2_522 ( .gnd(gnd), .vdd(vdd), .A(_8950_), .B(_8705__bF_buf6), .Y(_8699__220_) );
INVX2 INVX2_276 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_149_), .Y(_8951_) );
INVX1 INVX1_612 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_197_), .Y(_8952_) );
OAI21X1 OAI21X1_2517 ( .gnd(gnd), .vdd(vdd), .A(_8951_), .B(micro_hash_ucr_3_Wx_109_), .C(_8952_), .Y(_8953_) );
AOI21X1 AOI21X1_1556 ( .gnd(gnd), .vdd(vdd), .A(_8951_), .B(micro_hash_ucr_3_Wx_109_), .C(_8953_), .Y(_8954_) );
NOR2X1 NOR2X1_1398 ( .gnd(gnd), .vdd(vdd), .A(_8954_), .B(_8800__bF_buf9), .Y(_8699__221_) );
INVX4 INVX4_111 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_150_), .Y(_8955_) );
INVX2 INVX2_277 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_198_), .Y(_8956_) );
OAI21X1 OAI21X1_2518 ( .gnd(gnd), .vdd(vdd), .A(_8955_), .B(micro_hash_ucr_3_Wx_110_), .C(_8956_), .Y(_8957_) );
AOI21X1 AOI21X1_1557 ( .gnd(gnd), .vdd(vdd), .A(_8955_), .B(micro_hash_ucr_3_Wx_110_), .C(_8957_), .Y(_8958_) );
NOR2X1 NOR2X1_1399 ( .gnd(gnd), .vdd(vdd), .A(_8958_), .B(_8800__bF_buf8), .Y(_8699__222_) );
INVX4 INVX4_112 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_111_), .Y(_8959_) );
AOI21X1 AOI21X1_1558 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_151_), .B(_8959_), .C(micro_hash_ucr_3_Wx_199_), .Y(_8960_) );
OAI21X1 OAI21X1_2519 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_151_), .B(_8959_), .C(_8960_), .Y(_8961_) );
AND2X2 AND2X2_523 ( .gnd(gnd), .vdd(vdd), .A(_8961_), .B(_8705__bF_buf5), .Y(_8699__223_) );
INVX2 INVX2_278 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_160_), .Y(_8962_) );
INVX1 INVX1_613 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_208_), .Y(_8963_) );
OAI21X1 OAI21X1_2520 ( .gnd(gnd), .vdd(vdd), .A(_8962_), .B(micro_hash_ucr_3_Wx_120_), .C(_8963_), .Y(_8964_) );
AOI21X1 AOI21X1_1559 ( .gnd(gnd), .vdd(vdd), .A(_8962_), .B(micro_hash_ucr_3_Wx_120_), .C(_8964_), .Y(_8965_) );
NOR2X1 NOR2X1_1400 ( .gnd(gnd), .vdd(vdd), .A(_8965_), .B(_8800__bF_buf7), .Y(_8699__232_) );
INVX2 INVX2_279 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_161_), .Y(_8966_) );
INVX2 INVX2_280 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_209_), .Y(_8967_) );
OAI21X1 OAI21X1_2521 ( .gnd(gnd), .vdd(vdd), .A(_8966_), .B(micro_hash_ucr_3_Wx_121_), .C(_8967_), .Y(_8968_) );
AOI21X1 AOI21X1_1560 ( .gnd(gnd), .vdd(vdd), .A(_8966_), .B(micro_hash_ucr_3_Wx_121_), .C(_8968_), .Y(_8969_) );
NOR2X1 NOR2X1_1401 ( .gnd(gnd), .vdd(vdd), .A(_8969_), .B(_8800__bF_buf6), .Y(_8699__233_) );
INVX4 INVX4_113 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_162_), .Y(_8970_) );
INVX2 INVX2_281 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_210_), .Y(_8971_) );
OAI21X1 OAI21X1_2522 ( .gnd(gnd), .vdd(vdd), .A(_8970_), .B(micro_hash_ucr_3_Wx_122_), .C(_8971_), .Y(_8972_) );
AOI21X1 AOI21X1_1561 ( .gnd(gnd), .vdd(vdd), .A(_8970_), .B(micro_hash_ucr_3_Wx_122_), .C(_8972_), .Y(_8973_) );
NOR2X1 NOR2X1_1402 ( .gnd(gnd), .vdd(vdd), .A(_8973_), .B(_8800__bF_buf5), .Y(_8699__234_) );
INVX2 INVX2_282 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_163_), .Y(_8974_) );
INVX1 INVX1_614 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_211_), .Y(_8975_) );
OAI21X1 OAI21X1_2523 ( .gnd(gnd), .vdd(vdd), .A(_8974_), .B(micro_hash_ucr_3_Wx_123_), .C(_8975_), .Y(_8976_) );
AOI21X1 AOI21X1_1562 ( .gnd(gnd), .vdd(vdd), .A(_8974_), .B(micro_hash_ucr_3_Wx_123_), .C(_8976_), .Y(_8977_) );
NOR2X1 NOR2X1_1403 ( .gnd(gnd), .vdd(vdd), .A(_8977_), .B(_8800__bF_buf4), .Y(_8699__235_) );
INVX4 INVX4_114 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_124_), .Y(_8978_) );
AOI21X1 AOI21X1_1563 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_164_), .B(_8978_), .C(micro_hash_ucr_3_Wx_212_), .Y(_8979_) );
OAI21X1 OAI21X1_2524 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_164_), .B(_8978_), .C(_8979_), .Y(_8980_) );
AND2X2 AND2X2_524 ( .gnd(gnd), .vdd(vdd), .A(_8980_), .B(_8705__bF_buf4), .Y(_8699__236_) );
INVX2 INVX2_283 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_165_), .Y(_8981_) );
INVX1 INVX1_615 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_213_), .Y(_8982_) );
OAI21X1 OAI21X1_2525 ( .gnd(gnd), .vdd(vdd), .A(_8981_), .B(micro_hash_ucr_3_Wx_125_), .C(_8982_), .Y(_8983_) );
AOI21X1 AOI21X1_1564 ( .gnd(gnd), .vdd(vdd), .A(_8981_), .B(micro_hash_ucr_3_Wx_125_), .C(_8983_), .Y(_8984_) );
NOR2X1 NOR2X1_1404 ( .gnd(gnd), .vdd(vdd), .A(_8984_), .B(_8800__bF_buf3), .Y(_8699__237_) );
INVX4 INVX4_115 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_126_), .Y(_8985_) );
AOI21X1 AOI21X1_1565 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_166_), .B(_8985_), .C(micro_hash_ucr_3_Wx_214_), .Y(_8986_) );
OAI21X1 OAI21X1_2526 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_166_), .B(_8985_), .C(_8986_), .Y(_8987_) );
AND2X2 AND2X2_525 ( .gnd(gnd), .vdd(vdd), .A(_8987_), .B(_8705__bF_buf3), .Y(_8699__238_) );
INVX4 INVX4_116 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_167_), .Y(_8988_) );
AOI21X1 AOI21X1_1566 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_127_), .B(_8988_), .C(micro_hash_ucr_3_Wx_215_), .Y(_8989_) );
OAI21X1 OAI21X1_2527 ( .gnd(gnd), .vdd(vdd), .A(_8988_), .B(micro_hash_ucr_3_Wx_127_), .C(_8989_), .Y(_8990_) );
AND2X2 AND2X2_526 ( .gnd(gnd), .vdd(vdd), .A(_8990_), .B(_8705__bF_buf2), .Y(_8699__239_) );
INVX2 INVX2_284 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_152_), .Y(_8991_) );
AOI21X1 AOI21X1_1567 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_112_), .B(_8991_), .C(micro_hash_ucr_3_Wx_200_), .Y(_8992_) );
OAI21X1 OAI21X1_2528 ( .gnd(gnd), .vdd(vdd), .A(_8991_), .B(micro_hash_ucr_3_Wx_112_), .C(_8992_), .Y(_8993_) );
AND2X2 AND2X2_527 ( .gnd(gnd), .vdd(vdd), .A(_8993_), .B(_8705__bF_buf1), .Y(_8699__224_) );
INVX2 INVX2_285 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_153_), .Y(_8994_) );
AOI21X1 AOI21X1_1568 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_113_), .B(_8994_), .C(micro_hash_ucr_3_Wx_201_), .Y(_8995_) );
OAI21X1 OAI21X1_2529 ( .gnd(gnd), .vdd(vdd), .A(_8994_), .B(micro_hash_ucr_3_Wx_113_), .C(_8995_), .Y(_8996_) );
AND2X2 AND2X2_528 ( .gnd(gnd), .vdd(vdd), .A(_8996_), .B(_8705__bF_buf0), .Y(_8699__225_) );
INVX4 INVX4_117 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_154_), .Y(_8997_) );
INVX2 INVX2_286 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_202_), .Y(_8998_) );
OAI21X1 OAI21X1_2530 ( .gnd(gnd), .vdd(vdd), .A(_8997_), .B(micro_hash_ucr_3_Wx_114_), .C(_8998_), .Y(_8999_) );
AOI21X1 AOI21X1_1569 ( .gnd(gnd), .vdd(vdd), .A(_8997_), .B(micro_hash_ucr_3_Wx_114_), .C(_8999_), .Y(_9000_) );
NOR2X1 NOR2X1_1405 ( .gnd(gnd), .vdd(vdd), .A(_9000_), .B(_8800__bF_buf2), .Y(_8699__226_) );
INVX2 INVX2_287 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_155_), .Y(_9001_) );
INVX1 INVX1_616 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_203_), .Y(_9002_) );
OAI21X1 OAI21X1_2531 ( .gnd(gnd), .vdd(vdd), .A(_9001_), .B(micro_hash_ucr_3_Wx_115_), .C(_9002_), .Y(_9003_) );
AOI21X1 AOI21X1_1570 ( .gnd(gnd), .vdd(vdd), .A(_9001_), .B(micro_hash_ucr_3_Wx_115_), .C(_9003_), .Y(_9004_) );
NOR2X1 NOR2X1_1406 ( .gnd(gnd), .vdd(vdd), .A(_9004_), .B(_8800__bF_buf1), .Y(_8699__227_) );
INVX2 INVX2_288 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_156_), .Y(_9005_) );
AOI21X1 AOI21X1_1571 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_116_), .B(_9005_), .C(micro_hash_ucr_3_Wx_204_), .Y(_9006_) );
OAI21X1 OAI21X1_2532 ( .gnd(gnd), .vdd(vdd), .A(_9005_), .B(micro_hash_ucr_3_Wx_116_), .C(_9006_), .Y(_9007_) );
AND2X2 AND2X2_529 ( .gnd(gnd), .vdd(vdd), .A(_9007_), .B(_8705__bF_buf13), .Y(_8699__228_) );
INVX2 INVX2_289 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_157_), .Y(_9008_) );
AOI21X1 AOI21X1_1572 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_117_), .B(_9008_), .C(micro_hash_ucr_3_Wx_205_), .Y(_9009_) );
OAI21X1 OAI21X1_2533 ( .gnd(gnd), .vdd(vdd), .A(_9008_), .B(micro_hash_ucr_3_Wx_117_), .C(_9009_), .Y(_9010_) );
AND2X2 AND2X2_530 ( .gnd(gnd), .vdd(vdd), .A(_9010_), .B(_8705__bF_buf12), .Y(_8699__229_) );
INVX2 INVX2_290 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_158_), .Y(_9011_) );
INVX2 INVX2_291 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_206_), .Y(_9012_) );
OAI21X1 OAI21X1_2534 ( .gnd(gnd), .vdd(vdd), .A(_9011_), .B(micro_hash_ucr_3_Wx_118_), .C(_9012_), .Y(_9013_) );
AOI21X1 AOI21X1_1573 ( .gnd(gnd), .vdd(vdd), .A(_9011_), .B(micro_hash_ucr_3_Wx_118_), .C(_9013_), .Y(_9014_) );
NOR2X1 NOR2X1_1407 ( .gnd(gnd), .vdd(vdd), .A(_9014_), .B(_8800__bF_buf0), .Y(_8699__230_) );
INVX4 INVX4_118 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_159_), .Y(_9015_) );
AOI21X1 AOI21X1_1574 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_119_), .B(_9015_), .C(micro_hash_ucr_3_Wx_207_), .Y(_9016_) );
OAI21X1 OAI21X1_2535 ( .gnd(gnd), .vdd(vdd), .A(_9015_), .B(micro_hash_ucr_3_Wx_119_), .C(_9016_), .Y(_9017_) );
AND2X2 AND2X2_531 ( .gnd(gnd), .vdd(vdd), .A(_9017_), .B(_8705__bF_buf11), .Y(_8699__231_) );
INVX2 INVX2_292 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_120_), .Y(_9018_) );
AOI21X1 AOI21X1_1575 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_80_), .B(_9018_), .C(micro_hash_ucr_3_Wx_168_), .Y(_9019_) );
OAI21X1 OAI21X1_2536 ( .gnd(gnd), .vdd(vdd), .A(_9018_), .B(micro_hash_ucr_3_Wx_80_), .C(_9019_), .Y(_9020_) );
AND2X2 AND2X2_532 ( .gnd(gnd), .vdd(vdd), .A(_9020_), .B(_8705__bF_buf10), .Y(_8699__192_) );
INVX2 INVX2_293 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_121_), .Y(_9021_) );
OAI21X1 OAI21X1_2537 ( .gnd(gnd), .vdd(vdd), .A(_9021_), .B(micro_hash_ucr_3_Wx_81_), .C(_8836_), .Y(_9022_) );
AOI21X1 AOI21X1_1576 ( .gnd(gnd), .vdd(vdd), .A(_9021_), .B(micro_hash_ucr_3_Wx_81_), .C(_9022_), .Y(_9023_) );
NOR2X1 NOR2X1_1408 ( .gnd(gnd), .vdd(vdd), .A(_9023_), .B(_8800__bF_buf12), .Y(_8699__193_) );
INVX4 INVX4_119 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_122_), .Y(_9024_) );
OAI21X1 OAI21X1_2538 ( .gnd(gnd), .vdd(vdd), .A(_9024_), .B(micro_hash_ucr_3_Wx_82_), .C(_8840_), .Y(_9025_) );
AOI21X1 AOI21X1_1577 ( .gnd(gnd), .vdd(vdd), .A(_9024_), .B(micro_hash_ucr_3_Wx_82_), .C(_9025_), .Y(_9026_) );
NOR2X1 NOR2X1_1409 ( .gnd(gnd), .vdd(vdd), .A(_9026_), .B(_8800__bF_buf11), .Y(_8699__194_) );
INVX2 INVX2_294 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_123_), .Y(_9027_) );
OAI21X1 OAI21X1_2539 ( .gnd(gnd), .vdd(vdd), .A(_9027_), .B(micro_hash_ucr_3_Wx_83_), .C(_8844_), .Y(_9028_) );
AOI21X1 AOI21X1_1578 ( .gnd(gnd), .vdd(vdd), .A(_9027_), .B(micro_hash_ucr_3_Wx_83_), .C(_9028_), .Y(_9029_) );
NOR2X1 NOR2X1_1410 ( .gnd(gnd), .vdd(vdd), .A(_9029_), .B(_8800__bF_buf10), .Y(_8699__195_) );
OAI21X1 OAI21X1_2540 ( .gnd(gnd), .vdd(vdd), .A(_8978_), .B(micro_hash_ucr_3_Wx_84_), .C(_8848_), .Y(_9030_) );
AOI21X1 AOI21X1_1579 ( .gnd(gnd), .vdd(vdd), .A(_8978_), .B(micro_hash_ucr_3_Wx_84_), .C(_9030_), .Y(_9031_) );
NOR2X1 NOR2X1_1411 ( .gnd(gnd), .vdd(vdd), .A(_9031_), .B(_8800__bF_buf9), .Y(_8699__196_) );
INVX2 INVX2_295 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_125_), .Y(_9032_) );
OAI21X1 OAI21X1_2541 ( .gnd(gnd), .vdd(vdd), .A(_9032_), .B(micro_hash_ucr_3_Wx_85_), .C(_8851_), .Y(_9033_) );
AOI21X1 AOI21X1_1580 ( .gnd(gnd), .vdd(vdd), .A(_9032_), .B(micro_hash_ucr_3_Wx_85_), .C(_9033_), .Y(_9034_) );
NOR2X1 NOR2X1_1412 ( .gnd(gnd), .vdd(vdd), .A(_9034_), .B(_8800__bF_buf8), .Y(_8699__197_) );
OAI21X1 OAI21X1_2542 ( .gnd(gnd), .vdd(vdd), .A(_8985_), .B(micro_hash_ucr_3_Wx_86_), .C(_8854_), .Y(_9035_) );
AOI21X1 AOI21X1_1581 ( .gnd(gnd), .vdd(vdd), .A(_8985_), .B(micro_hash_ucr_3_Wx_86_), .C(_9035_), .Y(_9036_) );
NOR2X1 NOR2X1_1413 ( .gnd(gnd), .vdd(vdd), .A(_9036_), .B(_8800__bF_buf7), .Y(_8699__198_) );
INVX2 INVX2_296 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_87_), .Y(_9037_) );
AOI21X1 AOI21X1_1582 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_127_), .B(_9037_), .C(micro_hash_ucr_3_Wx_175_), .Y(_9038_) );
OAI21X1 OAI21X1_2543 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_127_), .B(_9037_), .C(_9038_), .Y(_9039_) );
AND2X2 AND2X2_533 ( .gnd(gnd), .vdd(vdd), .A(_9039_), .B(_8705__bF_buf9), .Y(_8699__199_) );
INVX4 INVX4_120 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_96_), .Y(_9040_) );
AOI21X1 AOI21X1_1583 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_136_), .B(_9040_), .C(micro_hash_ucr_3_Wx_184_), .Y(_9041_) );
OAI21X1 OAI21X1_2544 ( .gnd(gnd), .vdd(vdd), .A(_9040_), .B(micro_hash_ucr_3_Wx_136_), .C(_9041_), .Y(_9042_) );
AND2X2 AND2X2_534 ( .gnd(gnd), .vdd(vdd), .A(_9042_), .B(_8705__bF_buf8), .Y(_8699__208_) );
INVX4 INVX4_121 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_97_), .Y(_9043_) );
INVX1 INVX1_617 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_185_), .Y(_9044_) );
OAI21X1 OAI21X1_2545 ( .gnd(gnd), .vdd(vdd), .A(_9043_), .B(micro_hash_ucr_3_Wx_137_), .C(_9044_), .Y(_9045_) );
AOI21X1 AOI21X1_1584 ( .gnd(gnd), .vdd(vdd), .A(_9043_), .B(micro_hash_ucr_3_Wx_137_), .C(_9045_), .Y(_9046_) );
NOR2X1 NOR2X1_1414 ( .gnd(gnd), .vdd(vdd), .A(_9046_), .B(_8800__bF_buf6), .Y(_8699__209_) );
INVX4 INVX4_122 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_98_), .Y(_9047_) );
INVX2 INVX2_297 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_186_), .Y(_9048_) );
OAI21X1 OAI21X1_2546 ( .gnd(gnd), .vdd(vdd), .A(_9047_), .B(micro_hash_ucr_3_Wx_138_), .C(_9048_), .Y(_9049_) );
AOI21X1 AOI21X1_1585 ( .gnd(gnd), .vdd(vdd), .A(_9047_), .B(micro_hash_ucr_3_Wx_138_), .C(_9049_), .Y(_9050_) );
NOR2X1 NOR2X1_1415 ( .gnd(gnd), .vdd(vdd), .A(_9050_), .B(_8800__bF_buf5), .Y(_8699__210_) );
INVX4 INVX4_123 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_99_), .Y(_9051_) );
INVX1 INVX1_618 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_187_), .Y(_9052_) );
OAI21X1 OAI21X1_2547 ( .gnd(gnd), .vdd(vdd), .A(_9051_), .B(micro_hash_ucr_3_Wx_139_), .C(_9052_), .Y(_9053_) );
AOI21X1 AOI21X1_1586 ( .gnd(gnd), .vdd(vdd), .A(_9051_), .B(micro_hash_ucr_3_Wx_139_), .C(_9053_), .Y(_9054_) );
NOR2X1 NOR2X1_1416 ( .gnd(gnd), .vdd(vdd), .A(_9054_), .B(_8800__bF_buf4), .Y(_8699__211_) );
INVX4 INVX4_124 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_100_), .Y(_9055_) );
AOI21X1 AOI21X1_1587 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_140_), .B(_9055_), .C(micro_hash_ucr_3_Wx_188_), .Y(_9056_) );
OAI21X1 OAI21X1_2548 ( .gnd(gnd), .vdd(vdd), .A(_9055_), .B(micro_hash_ucr_3_Wx_140_), .C(_9056_), .Y(_9057_) );
AND2X2 AND2X2_535 ( .gnd(gnd), .vdd(vdd), .A(_9057_), .B(_8705__bF_buf7), .Y(_8699__212_) );
INVX4 INVX4_125 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_101_), .Y(_9058_) );
AOI21X1 AOI21X1_1588 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_141_), .B(_9058_), .C(micro_hash_ucr_3_Wx_189_), .Y(_9059_) );
OAI21X1 OAI21X1_2549 ( .gnd(gnd), .vdd(vdd), .A(_9058_), .B(micro_hash_ucr_3_Wx_141_), .C(_9059_), .Y(_9060_) );
AND2X2 AND2X2_536 ( .gnd(gnd), .vdd(vdd), .A(_9060_), .B(_8705__bF_buf6), .Y(_8699__213_) );
INVX4 INVX4_126 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_102_), .Y(_9061_) );
INVX2 INVX2_298 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_190_), .Y(_9062_) );
OAI21X1 OAI21X1_2550 ( .gnd(gnd), .vdd(vdd), .A(_9061_), .B(micro_hash_ucr_3_Wx_142_), .C(_9062_), .Y(_9063_) );
AOI21X1 AOI21X1_1589 ( .gnd(gnd), .vdd(vdd), .A(_9061_), .B(micro_hash_ucr_3_Wx_142_), .C(_9063_), .Y(_9064_) );
NOR2X1 NOR2X1_1417 ( .gnd(gnd), .vdd(vdd), .A(_9064_), .B(_8800__bF_buf3), .Y(_8699__214_) );
INVX4 INVX4_127 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_103_), .Y(_9065_) );
AOI21X1 AOI21X1_1590 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_143_), .B(_9065_), .C(micro_hash_ucr_3_Wx_191_), .Y(_9066_) );
OAI21X1 OAI21X1_2551 ( .gnd(gnd), .vdd(vdd), .A(_9065_), .B(micro_hash_ucr_3_Wx_143_), .C(_9066_), .Y(_9067_) );
AND2X2 AND2X2_537 ( .gnd(gnd), .vdd(vdd), .A(_9067_), .B(_8705__bF_buf5), .Y(_8699__215_) );
INVX2 INVX2_299 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_128_), .Y(_9068_) );
INVX1 INVX1_619 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_176_), .Y(_9069_) );
OAI21X1 OAI21X1_2552 ( .gnd(gnd), .vdd(vdd), .A(_9068_), .B(micro_hash_ucr_3_Wx_88_), .C(_9069_), .Y(_9070_) );
AOI21X1 AOI21X1_1591 ( .gnd(gnd), .vdd(vdd), .A(_9068_), .B(micro_hash_ucr_3_Wx_88_), .C(_9070_), .Y(_9071_) );
NOR2X1 NOR2X1_1418 ( .gnd(gnd), .vdd(vdd), .A(_9071_), .B(_8800__bF_buf2), .Y(_8699__200_) );
INVX2 INVX2_300 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_129_), .Y(_9072_) );
INVX1 INVX1_620 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_177_), .Y(_9073_) );
OAI21X1 OAI21X1_2553 ( .gnd(gnd), .vdd(vdd), .A(_9072_), .B(micro_hash_ucr_3_Wx_89_), .C(_9073_), .Y(_9074_) );
AOI21X1 AOI21X1_1592 ( .gnd(gnd), .vdd(vdd), .A(_9072_), .B(micro_hash_ucr_3_Wx_89_), .C(_9074_), .Y(_9075_) );
NOR2X1 NOR2X1_1419 ( .gnd(gnd), .vdd(vdd), .A(_9075_), .B(_8800__bF_buf1), .Y(_8699__201_) );
INVX4 INVX4_128 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_130_), .Y(_9076_) );
INVX2 INVX2_301 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_178_), .Y(_9077_) );
OAI21X1 OAI21X1_2554 ( .gnd(gnd), .vdd(vdd), .A(_9076_), .B(micro_hash_ucr_3_Wx_90_), .C(_9077_), .Y(_9078_) );
AOI21X1 AOI21X1_1593 ( .gnd(gnd), .vdd(vdd), .A(_9076_), .B(micro_hash_ucr_3_Wx_90_), .C(_9078_), .Y(_9079_) );
NOR2X1 NOR2X1_1420 ( .gnd(gnd), .vdd(vdd), .A(_9079_), .B(_8800__bF_buf0), .Y(_8699__202_) );
INVX2 INVX2_302 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_131_), .Y(_9080_) );
INVX1 INVX1_621 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_179_), .Y(_9081_) );
OAI21X1 OAI21X1_2555 ( .gnd(gnd), .vdd(vdd), .A(_9080_), .B(micro_hash_ucr_3_Wx_91_), .C(_9081_), .Y(_9082_) );
AOI21X1 AOI21X1_1594 ( .gnd(gnd), .vdd(vdd), .A(_9080_), .B(micro_hash_ucr_3_Wx_91_), .C(_9082_), .Y(_9083_) );
NOR2X1 NOR2X1_1421 ( .gnd(gnd), .vdd(vdd), .A(_9083_), .B(_8800__bF_buf12), .Y(_8699__203_) );
INVX2 INVX2_303 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_132_), .Y(_9084_) );
INVX2 INVX2_304 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_180_), .Y(_9085_) );
OAI21X1 OAI21X1_2556 ( .gnd(gnd), .vdd(vdd), .A(_9084_), .B(micro_hash_ucr_3_Wx_92_), .C(_9085_), .Y(_9086_) );
AOI21X1 AOI21X1_1595 ( .gnd(gnd), .vdd(vdd), .A(_9084_), .B(micro_hash_ucr_3_Wx_92_), .C(_9086_), .Y(_9087_) );
NOR2X1 NOR2X1_1422 ( .gnd(gnd), .vdd(vdd), .A(_9087_), .B(_8800__bF_buf11), .Y(_8699__204_) );
INVX2 INVX2_305 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_133_), .Y(_9088_) );
INVX1 INVX1_622 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_181_), .Y(_9089_) );
OAI21X1 OAI21X1_2557 ( .gnd(gnd), .vdd(vdd), .A(_9088_), .B(micro_hash_ucr_3_Wx_93_), .C(_9089_), .Y(_9090_) );
AOI21X1 AOI21X1_1596 ( .gnd(gnd), .vdd(vdd), .A(_9088_), .B(micro_hash_ucr_3_Wx_93_), .C(_9090_), .Y(_9091_) );
NOR2X1 NOR2X1_1423 ( .gnd(gnd), .vdd(vdd), .A(_9091_), .B(_8800__bF_buf10), .Y(_8699__205_) );
INVX4 INVX4_129 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_134_), .Y(_9092_) );
INVX2 INVX2_306 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_182_), .Y(_9093_) );
OAI21X1 OAI21X1_2558 ( .gnd(gnd), .vdd(vdd), .A(_9092_), .B(micro_hash_ucr_3_Wx_94_), .C(_9093_), .Y(_9094_) );
AOI21X1 AOI21X1_1597 ( .gnd(gnd), .vdd(vdd), .A(_9092_), .B(micro_hash_ucr_3_Wx_94_), .C(_9094_), .Y(_9095_) );
NOR2X1 NOR2X1_1424 ( .gnd(gnd), .vdd(vdd), .A(_9095_), .B(_8800__bF_buf9), .Y(_8699__206_) );
INVX2 INVX2_307 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_183_), .Y(_9096_) );
XNOR2X1 XNOR2X1_388 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_135_), .B(micro_hash_ucr_3_Wx_95_), .Y(_9097_) );
AOI21X1 AOI21X1_1598 ( .gnd(gnd), .vdd(vdd), .A(_9096_), .B(_9097_), .C(_8800__bF_buf8), .Y(_8699__207_) );
OAI21X1 OAI21X1_2559 ( .gnd(gnd), .vdd(vdd), .A(_9040_), .B(micro_hash_ucr_3_Wx_56_), .C(_8932_), .Y(_9098_) );
AOI21X1 AOI21X1_1599 ( .gnd(gnd), .vdd(vdd), .A(_9040_), .B(micro_hash_ucr_3_Wx_56_), .C(_9098_), .Y(_9099_) );
NOR2X1 NOR2X1_1425 ( .gnd(gnd), .vdd(vdd), .A(_9099_), .B(_8800__bF_buf7), .Y(_8699__168_) );
OAI21X1 OAI21X1_2560 ( .gnd(gnd), .vdd(vdd), .A(_9043_), .B(micro_hash_ucr_3_Wx_57_), .C(_8936_), .Y(_9100_) );
AOI21X1 AOI21X1_1600 ( .gnd(gnd), .vdd(vdd), .A(_9043_), .B(micro_hash_ucr_3_Wx_57_), .C(_9100_), .Y(_9101_) );
NOR2X1 NOR2X1_1426 ( .gnd(gnd), .vdd(vdd), .A(_9101_), .B(_8800__bF_buf6), .Y(_8699__169_) );
OAI21X1 OAI21X1_2561 ( .gnd(gnd), .vdd(vdd), .A(_9047_), .B(micro_hash_ucr_3_Wx_58_), .C(_8940_), .Y(_9102_) );
AOI21X1 AOI21X1_1601 ( .gnd(gnd), .vdd(vdd), .A(_9047_), .B(micro_hash_ucr_3_Wx_58_), .C(_9102_), .Y(_9103_) );
NOR2X1 NOR2X1_1427 ( .gnd(gnd), .vdd(vdd), .A(_9103_), .B(_8800__bF_buf5), .Y(_8699__170_) );
OAI21X1 OAI21X1_2562 ( .gnd(gnd), .vdd(vdd), .A(_9051_), .B(micro_hash_ucr_3_Wx_59_), .C(_8944_), .Y(_9104_) );
AOI21X1 AOI21X1_1602 ( .gnd(gnd), .vdd(vdd), .A(_9051_), .B(micro_hash_ucr_3_Wx_59_), .C(_9104_), .Y(_9105_) );
NOR2X1 NOR2X1_1428 ( .gnd(gnd), .vdd(vdd), .A(_9105_), .B(_8800__bF_buf4), .Y(_8699__171_) );
OAI21X1 OAI21X1_2563 ( .gnd(gnd), .vdd(vdd), .A(_9055_), .B(micro_hash_ucr_3_Wx_60_), .C(_8948_), .Y(_9106_) );
AOI21X1 AOI21X1_1603 ( .gnd(gnd), .vdd(vdd), .A(_9055_), .B(micro_hash_ucr_3_Wx_60_), .C(_9106_), .Y(_9107_) );
NOR2X1 NOR2X1_1429 ( .gnd(gnd), .vdd(vdd), .A(_9107_), .B(_8800__bF_buf3), .Y(_8699__172_) );
OAI21X1 OAI21X1_2564 ( .gnd(gnd), .vdd(vdd), .A(_9058_), .B(micro_hash_ucr_3_Wx_61_), .C(_8951_), .Y(_9108_) );
AOI21X1 AOI21X1_1604 ( .gnd(gnd), .vdd(vdd), .A(_9058_), .B(micro_hash_ucr_3_Wx_61_), .C(_9108_), .Y(_9109_) );
NOR2X1 NOR2X1_1430 ( .gnd(gnd), .vdd(vdd), .A(_9109_), .B(_8800__bF_buf2), .Y(_8699__173_) );
OAI21X1 OAI21X1_2565 ( .gnd(gnd), .vdd(vdd), .A(_9061_), .B(micro_hash_ucr_3_Wx_62_), .C(_8955_), .Y(_9110_) );
AOI21X1 AOI21X1_1605 ( .gnd(gnd), .vdd(vdd), .A(_9061_), .B(micro_hash_ucr_3_Wx_62_), .C(_9110_), .Y(_9111_) );
NOR2X1 NOR2X1_1431 ( .gnd(gnd), .vdd(vdd), .A(_9111_), .B(_8800__bF_buf1), .Y(_8699__174_) );
AOI21X1 AOI21X1_1606 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_63_), .B(_9065_), .C(micro_hash_ucr_3_Wx_151_), .Y(_9112_) );
OAI21X1 OAI21X1_2566 ( .gnd(gnd), .vdd(vdd), .A(_9065_), .B(micro_hash_ucr_3_Wx_63_), .C(_9112_), .Y(_9113_) );
AND2X2 AND2X2_538 ( .gnd(gnd), .vdd(vdd), .A(_9113_), .B(_8705__bF_buf4), .Y(_8699__175_) );
INVX2 INVX2_308 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_112_), .Y(_9114_) );
OAI21X1 OAI21X1_2567 ( .gnd(gnd), .vdd(vdd), .A(_9114_), .B(micro_hash_ucr_3_Wx_72_), .C(_8962_), .Y(_9115_) );
AOI21X1 AOI21X1_1607 ( .gnd(gnd), .vdd(vdd), .A(_9114_), .B(micro_hash_ucr_3_Wx_72_), .C(_9115_), .Y(_9116_) );
NOR2X1 NOR2X1_1432 ( .gnd(gnd), .vdd(vdd), .A(_9116_), .B(_8800__bF_buf0), .Y(_8699__184_) );
INVX2 INVX2_309 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_113_), .Y(_9117_) );
OAI21X1 OAI21X1_2568 ( .gnd(gnd), .vdd(vdd), .A(_9117_), .B(micro_hash_ucr_3_Wx_73_), .C(_8966_), .Y(_9118_) );
AOI21X1 AOI21X1_1608 ( .gnd(gnd), .vdd(vdd), .A(_9117_), .B(micro_hash_ucr_3_Wx_73_), .C(_9118_), .Y(_9119_) );
NOR2X1 NOR2X1_1433 ( .gnd(gnd), .vdd(vdd), .A(_9119_), .B(_8800__bF_buf12), .Y(_8699__185_) );
INVX4 INVX4_130 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_114_), .Y(_9120_) );
OAI21X1 OAI21X1_2569 ( .gnd(gnd), .vdd(vdd), .A(_9120_), .B(micro_hash_ucr_3_Wx_74_), .C(_8970_), .Y(_9121_) );
AOI21X1 AOI21X1_1609 ( .gnd(gnd), .vdd(vdd), .A(_9120_), .B(micro_hash_ucr_3_Wx_74_), .C(_9121_), .Y(_9122_) );
NOR2X1 NOR2X1_1434 ( .gnd(gnd), .vdd(vdd), .A(_9122_), .B(_8800__bF_buf11), .Y(_8699__186_) );
INVX2 INVX2_310 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_115_), .Y(_9123_) );
OAI21X1 OAI21X1_2570 ( .gnd(gnd), .vdd(vdd), .A(_9123_), .B(micro_hash_ucr_3_Wx_75_), .C(_8974_), .Y(_9124_) );
AOI21X1 AOI21X1_1610 ( .gnd(gnd), .vdd(vdd), .A(_9123_), .B(micro_hash_ucr_3_Wx_75_), .C(_9124_), .Y(_9125_) );
NOR2X1 NOR2X1_1435 ( .gnd(gnd), .vdd(vdd), .A(_9125_), .B(_8800__bF_buf10), .Y(_8699__187_) );
INVX2 INVX2_311 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_116_), .Y(_9126_) );
AOI21X1 AOI21X1_1611 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_76_), .B(_9126_), .C(micro_hash_ucr_3_Wx_164_), .Y(_9127_) );
OAI21X1 OAI21X1_2571 ( .gnd(gnd), .vdd(vdd), .A(_9126_), .B(micro_hash_ucr_3_Wx_76_), .C(_9127_), .Y(_9128_) );
AND2X2 AND2X2_539 ( .gnd(gnd), .vdd(vdd), .A(_9128_), .B(_8705__bF_buf3), .Y(_8699__188_) );
INVX2 INVX2_312 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_117_), .Y(_9129_) );
OAI21X1 OAI21X1_2572 ( .gnd(gnd), .vdd(vdd), .A(_9129_), .B(micro_hash_ucr_3_Wx_77_), .C(_8981_), .Y(_9130_) );
AOI21X1 AOI21X1_1612 ( .gnd(gnd), .vdd(vdd), .A(_9129_), .B(micro_hash_ucr_3_Wx_77_), .C(_9130_), .Y(_9131_) );
NOR2X1 NOR2X1_1436 ( .gnd(gnd), .vdd(vdd), .A(_9131_), .B(_8800__bF_buf9), .Y(_8699__189_) );
INVX4 INVX4_131 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_118_), .Y(_9132_) );
AOI21X1 AOI21X1_1613 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_78_), .B(_9132_), .C(micro_hash_ucr_3_Wx_166_), .Y(_9133_) );
OAI21X1 OAI21X1_2573 ( .gnd(gnd), .vdd(vdd), .A(_9132_), .B(micro_hash_ucr_3_Wx_78_), .C(_9133_), .Y(_9134_) );
AND2X2 AND2X2_540 ( .gnd(gnd), .vdd(vdd), .A(_9134_), .B(_8705__bF_buf2), .Y(_8699__190_) );
INVX4 INVX4_132 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_79_), .Y(_9135_) );
OAI21X1 OAI21X1_2574 ( .gnd(gnd), .vdd(vdd), .A(_9135_), .B(micro_hash_ucr_3_Wx_119_), .C(_8988_), .Y(_9136_) );
AOI21X1 AOI21X1_1614 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_119_), .B(_9135_), .C(_9136_), .Y(_9137_) );
NOR2X1 NOR2X1_1437 ( .gnd(gnd), .vdd(vdd), .A(_9137_), .B(_8800__bF_buf8), .Y(_8699__191_) );
XNOR2X1 XNOR2X1_389 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_104_), .B(micro_hash_ucr_3_Wx_64_), .Y(_9138_) );
AOI21X1 AOI21X1_1615 ( .gnd(gnd), .vdd(vdd), .A(_8991_), .B(_9138_), .C(_8800__bF_buf7), .Y(_8699__176_) );
INVX2 INVX2_313 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_105_), .Y(_9139_) );
OAI21X1 OAI21X1_2575 ( .gnd(gnd), .vdd(vdd), .A(_9139_), .B(micro_hash_ucr_3_Wx_65_), .C(_8994_), .Y(_9140_) );
AOI21X1 AOI21X1_1616 ( .gnd(gnd), .vdd(vdd), .A(_9139_), .B(micro_hash_ucr_3_Wx_65_), .C(_9140_), .Y(_9141_) );
NOR2X1 NOR2X1_1438 ( .gnd(gnd), .vdd(vdd), .A(_9141_), .B(_8800__bF_buf6), .Y(_8699__177_) );
INVX4 INVX4_133 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_106_), .Y(_9142_) );
OAI21X1 OAI21X1_2576 ( .gnd(gnd), .vdd(vdd), .A(_9142_), .B(micro_hash_ucr_3_Wx_66_), .C(_8997_), .Y(_9143_) );
AOI21X1 AOI21X1_1617 ( .gnd(gnd), .vdd(vdd), .A(_9142_), .B(micro_hash_ucr_3_Wx_66_), .C(_9143_), .Y(_9144_) );
NOR2X1 NOR2X1_1439 ( .gnd(gnd), .vdd(vdd), .A(_9144_), .B(_8800__bF_buf5), .Y(_8699__178_) );
INVX2 INVX2_314 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_107_), .Y(_9145_) );
OAI21X1 OAI21X1_2577 ( .gnd(gnd), .vdd(vdd), .A(_9145_), .B(micro_hash_ucr_3_Wx_67_), .C(_9001_), .Y(_9146_) );
AOI21X1 AOI21X1_1618 ( .gnd(gnd), .vdd(vdd), .A(_9145_), .B(micro_hash_ucr_3_Wx_67_), .C(_9146_), .Y(_9147_) );
NOR2X1 NOR2X1_1440 ( .gnd(gnd), .vdd(vdd), .A(_9147_), .B(_8800__bF_buf4), .Y(_8699__179_) );
INVX2 INVX2_315 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_68_), .Y(_9148_) );
OAI21X1 OAI21X1_2578 ( .gnd(gnd), .vdd(vdd), .A(_9148_), .B(micro_hash_ucr_3_Wx_108_), .C(_9005_), .Y(_9149_) );
AOI21X1 AOI21X1_1619 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_108_), .B(_9148_), .C(_9149_), .Y(_9150_) );
NOR2X1 NOR2X1_1441 ( .gnd(gnd), .vdd(vdd), .A(_9150_), .B(_8800__bF_buf3), .Y(_8699__180_) );
INVX2 INVX2_316 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_109_), .Y(_9151_) );
OAI21X1 OAI21X1_2579 ( .gnd(gnd), .vdd(vdd), .A(_9151_), .B(micro_hash_ucr_3_Wx_69_), .C(_9008_), .Y(_9152_) );
AOI21X1 AOI21X1_1620 ( .gnd(gnd), .vdd(vdd), .A(_9151_), .B(micro_hash_ucr_3_Wx_69_), .C(_9152_), .Y(_9153_) );
NOR2X1 NOR2X1_1442 ( .gnd(gnd), .vdd(vdd), .A(_9153_), .B(_8800__bF_buf2), .Y(_8699__181_) );
INVX2 INVX2_317 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_110_), .Y(_9154_) );
OAI21X1 OAI21X1_2580 ( .gnd(gnd), .vdd(vdd), .A(_9154_), .B(micro_hash_ucr_3_Wx_70_), .C(_9011_), .Y(_9155_) );
AOI21X1 AOI21X1_1621 ( .gnd(gnd), .vdd(vdd), .A(_9154_), .B(micro_hash_ucr_3_Wx_70_), .C(_9155_), .Y(_9156_) );
NOR2X1 NOR2X1_1443 ( .gnd(gnd), .vdd(vdd), .A(_9156_), .B(_8800__bF_buf1), .Y(_8699__182_) );
OAI21X1 OAI21X1_2581 ( .gnd(gnd), .vdd(vdd), .A(_8959_), .B(micro_hash_ucr_3_Wx_71_), .C(_9015_), .Y(_9157_) );
AOI21X1 AOI21X1_1622 ( .gnd(gnd), .vdd(vdd), .A(_8959_), .B(micro_hash_ucr_3_Wx_71_), .C(_9157_), .Y(_9158_) );
NOR2X1 NOR2X1_1444 ( .gnd(gnd), .vdd(vdd), .A(_9158_), .B(_8800__bF_buf0), .Y(_8699__183_) );
INVX2 INVX2_318 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_72_), .Y(_9159_) );
OAI21X1 OAI21X1_2582 ( .gnd(gnd), .vdd(vdd), .A(_9159_), .B(micro_hash_ucr_3_Wx_32_), .C(_9018_), .Y(_9160_) );
AOI21X1 AOI21X1_1623 ( .gnd(gnd), .vdd(vdd), .A(_9159_), .B(micro_hash_ucr_3_Wx_32_), .C(_9160_), .Y(_9161_) );
NOR2X1 NOR2X1_1445 ( .gnd(gnd), .vdd(vdd), .A(_9161_), .B(_8800__bF_buf12), .Y(_8699__144_) );
INVX2 INVX2_319 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_73_), .Y(_9162_) );
OAI21X1 OAI21X1_2583 ( .gnd(gnd), .vdd(vdd), .A(_9162_), .B(micro_hash_ucr_3_Wx_33_), .C(_9021_), .Y(_9163_) );
AOI21X1 AOI21X1_1624 ( .gnd(gnd), .vdd(vdd), .A(_9162_), .B(micro_hash_ucr_3_Wx_33_), .C(_9163_), .Y(_9164_) );
NOR2X1 NOR2X1_1446 ( .gnd(gnd), .vdd(vdd), .A(_9164_), .B(_8800__bF_buf11), .Y(_8699__145_) );
INVX4 INVX4_134 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_74_), .Y(_9165_) );
OAI21X1 OAI21X1_2584 ( .gnd(gnd), .vdd(vdd), .A(_9165_), .B(micro_hash_ucr_3_Wx_34_), .C(_9024_), .Y(_9166_) );
AOI21X1 AOI21X1_1625 ( .gnd(gnd), .vdd(vdd), .A(_9165_), .B(micro_hash_ucr_3_Wx_34_), .C(_9166_), .Y(_9167_) );
NOR2X1 NOR2X1_1447 ( .gnd(gnd), .vdd(vdd), .A(_9167_), .B(_8800__bF_buf10), .Y(_8699__146_) );
INVX2 INVX2_320 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_75_), .Y(_9168_) );
OAI21X1 OAI21X1_2585 ( .gnd(gnd), .vdd(vdd), .A(_9168_), .B(micro_hash_ucr_3_Wx_35_), .C(_9027_), .Y(_9169_) );
AOI21X1 AOI21X1_1626 ( .gnd(gnd), .vdd(vdd), .A(_9168_), .B(micro_hash_ucr_3_Wx_35_), .C(_9169_), .Y(_9170_) );
NOR2X1 NOR2X1_1448 ( .gnd(gnd), .vdd(vdd), .A(_9170_), .B(_8800__bF_buf9), .Y(_8699__147_) );
INVX2 INVX2_321 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_76_), .Y(_9171_) );
OAI21X1 OAI21X1_2586 ( .gnd(gnd), .vdd(vdd), .A(_9171_), .B(micro_hash_ucr_3_Wx_36_), .C(_8978_), .Y(_9172_) );
AOI21X1 AOI21X1_1627 ( .gnd(gnd), .vdd(vdd), .A(_9171_), .B(micro_hash_ucr_3_Wx_36_), .C(_9172_), .Y(_9173_) );
NOR2X1 NOR2X1_1449 ( .gnd(gnd), .vdd(vdd), .A(_9173_), .B(_8800__bF_buf8), .Y(_8699__148_) );
INVX2 INVX2_322 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_77_), .Y(_9174_) );
OAI21X1 OAI21X1_2587 ( .gnd(gnd), .vdd(vdd), .A(_9174_), .B(micro_hash_ucr_3_Wx_37_), .C(_9032_), .Y(_9175_) );
AOI21X1 AOI21X1_1628 ( .gnd(gnd), .vdd(vdd), .A(_9174_), .B(micro_hash_ucr_3_Wx_37_), .C(_9175_), .Y(_9176_) );
NOR2X1 NOR2X1_1450 ( .gnd(gnd), .vdd(vdd), .A(_9176_), .B(_8800__bF_buf7), .Y(_8699__149_) );
INVX2 INVX2_323 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_78_), .Y(_9177_) );
OAI21X1 OAI21X1_2588 ( .gnd(gnd), .vdd(vdd), .A(_9177_), .B(micro_hash_ucr_3_Wx_38_), .C(_8985_), .Y(_9178_) );
AOI21X1 AOI21X1_1629 ( .gnd(gnd), .vdd(vdd), .A(_9177_), .B(micro_hash_ucr_3_Wx_38_), .C(_9178_), .Y(_9179_) );
NOR2X1 NOR2X1_1451 ( .gnd(gnd), .vdd(vdd), .A(_9179_), .B(_8800__bF_buf6), .Y(_8699__150_) );
AOI21X1 AOI21X1_1630 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_39_), .B(_9135_), .C(micro_hash_ucr_3_Wx_127_), .Y(_9180_) );
OAI21X1 OAI21X1_2589 ( .gnd(gnd), .vdd(vdd), .A(_9135_), .B(micro_hash_ucr_3_Wx_39_), .C(_9180_), .Y(_9181_) );
AND2X2 AND2X2_541 ( .gnd(gnd), .vdd(vdd), .A(_9181_), .B(_8705__bF_buf1), .Y(_8699__151_) );
INVX2 INVX2_324 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_88_), .Y(_9182_) );
INVX2 INVX2_325 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_136_), .Y(_9183_) );
OAI21X1 OAI21X1_2590 ( .gnd(gnd), .vdd(vdd), .A(_9182_), .B(micro_hash_ucr_3_Wx_48_), .C(_9183_), .Y(_9184_) );
AOI21X1 AOI21X1_1631 ( .gnd(gnd), .vdd(vdd), .A(_9182_), .B(micro_hash_ucr_3_Wx_48_), .C(_9184_), .Y(_9185_) );
NOR2X1 NOR2X1_1452 ( .gnd(gnd), .vdd(vdd), .A(_9185_), .B(_8800__bF_buf5), .Y(_8699__160_) );
INVX2 INVX2_326 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_89_), .Y(_9186_) );
INVX2 INVX2_327 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_137_), .Y(_9187_) );
OAI21X1 OAI21X1_2591 ( .gnd(gnd), .vdd(vdd), .A(_9186_), .B(micro_hash_ucr_3_Wx_49_), .C(_9187_), .Y(_9188_) );
AOI21X1 AOI21X1_1632 ( .gnd(gnd), .vdd(vdd), .A(_9186_), .B(micro_hash_ucr_3_Wx_49_), .C(_9188_), .Y(_9189_) );
NOR2X1 NOR2X1_1453 ( .gnd(gnd), .vdd(vdd), .A(_9189_), .B(_8800__bF_buf4), .Y(_8699__161_) );
INVX2 INVX2_328 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_90_), .Y(_9190_) );
INVX4 INVX4_135 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_138_), .Y(_9191_) );
OAI21X1 OAI21X1_2592 ( .gnd(gnd), .vdd(vdd), .A(_9190_), .B(micro_hash_ucr_3_Wx_50_), .C(_9191_), .Y(_9192_) );
AOI21X1 AOI21X1_1633 ( .gnd(gnd), .vdd(vdd), .A(_9190_), .B(micro_hash_ucr_3_Wx_50_), .C(_9192_), .Y(_9193_) );
NOR2X1 NOR2X1_1454 ( .gnd(gnd), .vdd(vdd), .A(_9193_), .B(_8800__bF_buf3), .Y(_8699__162_) );
INVX2 INVX2_329 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_91_), .Y(_9194_) );
INVX2 INVX2_330 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_139_), .Y(_9195_) );
OAI21X1 OAI21X1_2593 ( .gnd(gnd), .vdd(vdd), .A(_9194_), .B(micro_hash_ucr_3_Wx_51_), .C(_9195_), .Y(_9196_) );
AOI21X1 AOI21X1_1634 ( .gnd(gnd), .vdd(vdd), .A(_9194_), .B(micro_hash_ucr_3_Wx_51_), .C(_9196_), .Y(_9197_) );
NOR2X1 NOR2X1_1455 ( .gnd(gnd), .vdd(vdd), .A(_9197_), .B(_8800__bF_buf2), .Y(_8699__163_) );
INVX2 INVX2_331 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_92_), .Y(_9198_) );
INVX2 INVX2_332 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_140_), .Y(_9199_) );
OAI21X1 OAI21X1_2594 ( .gnd(gnd), .vdd(vdd), .A(_9198_), .B(micro_hash_ucr_3_Wx_52_), .C(_9199_), .Y(_9200_) );
AOI21X1 AOI21X1_1635 ( .gnd(gnd), .vdd(vdd), .A(_9198_), .B(micro_hash_ucr_3_Wx_52_), .C(_9200_), .Y(_9201_) );
NOR2X1 NOR2X1_1456 ( .gnd(gnd), .vdd(vdd), .A(_9201_), .B(_8800__bF_buf1), .Y(_8699__164_) );
INVX2 INVX2_333 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_93_), .Y(_9202_) );
INVX2 INVX2_334 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_141_), .Y(_9203_) );
OAI21X1 OAI21X1_2595 ( .gnd(gnd), .vdd(vdd), .A(_9202_), .B(micro_hash_ucr_3_Wx_53_), .C(_9203_), .Y(_9204_) );
AOI21X1 AOI21X1_1636 ( .gnd(gnd), .vdd(vdd), .A(_9202_), .B(micro_hash_ucr_3_Wx_53_), .C(_9204_), .Y(_9205_) );
NOR2X1 NOR2X1_1457 ( .gnd(gnd), .vdd(vdd), .A(_9205_), .B(_8800__bF_buf0), .Y(_8699__165_) );
INVX4 INVX4_136 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_94_), .Y(_9206_) );
INVX4 INVX4_137 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_142_), .Y(_9207_) );
OAI21X1 OAI21X1_2596 ( .gnd(gnd), .vdd(vdd), .A(_9206_), .B(micro_hash_ucr_3_Wx_54_), .C(_9207_), .Y(_9208_) );
AOI21X1 AOI21X1_1637 ( .gnd(gnd), .vdd(vdd), .A(_9206_), .B(micro_hash_ucr_3_Wx_54_), .C(_9208_), .Y(_9209_) );
NOR2X1 NOR2X1_1458 ( .gnd(gnd), .vdd(vdd), .A(_9209_), .B(_8800__bF_buf12), .Y(_8699__166_) );
INVX1 INVX1_623 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_95_), .Y(_9210_) );
INVX2 INVX2_335 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_143_), .Y(_9211_) );
OAI21X1 OAI21X1_2597 ( .gnd(gnd), .vdd(vdd), .A(_9210_), .B(micro_hash_ucr_3_Wx_55_), .C(_9211_), .Y(_9212_) );
AOI21X1 AOI21X1_1638 ( .gnd(gnd), .vdd(vdd), .A(_9210_), .B(micro_hash_ucr_3_Wx_55_), .C(_9212_), .Y(_9213_) );
NOR2X1 NOR2X1_1459 ( .gnd(gnd), .vdd(vdd), .A(_9213_), .B(_8800__bF_buf11), .Y(_8699__167_) );
INVX2 INVX2_336 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_80_), .Y(_9214_) );
OAI21X1 OAI21X1_2598 ( .gnd(gnd), .vdd(vdd), .A(_9214_), .B(micro_hash_ucr_3_Wx_40_), .C(_9068_), .Y(_9215_) );
AOI21X1 AOI21X1_1639 ( .gnd(gnd), .vdd(vdd), .A(_9214_), .B(micro_hash_ucr_3_Wx_40_), .C(_9215_), .Y(_9216_) );
NOR2X1 NOR2X1_1460 ( .gnd(gnd), .vdd(vdd), .A(_9216_), .B(_8800__bF_buf10), .Y(_8699__152_) );
INVX2 INVX2_337 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_81_), .Y(_9217_) );
OAI21X1 OAI21X1_2599 ( .gnd(gnd), .vdd(vdd), .A(_9217_), .B(micro_hash_ucr_3_Wx_41_), .C(_9072_), .Y(_9218_) );
AOI21X1 AOI21X1_1640 ( .gnd(gnd), .vdd(vdd), .A(_9217_), .B(micro_hash_ucr_3_Wx_41_), .C(_9218_), .Y(_9219_) );
NOR2X1 NOR2X1_1461 ( .gnd(gnd), .vdd(vdd), .A(_9219_), .B(_8800__bF_buf9), .Y(_8699__153_) );
INVX2 INVX2_338 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_82_), .Y(_9220_) );
OAI21X1 OAI21X1_2600 ( .gnd(gnd), .vdd(vdd), .A(_9220_), .B(micro_hash_ucr_3_Wx_42_), .C(_9076_), .Y(_9221_) );
AOI21X1 AOI21X1_1641 ( .gnd(gnd), .vdd(vdd), .A(_9220_), .B(micro_hash_ucr_3_Wx_42_), .C(_9221_), .Y(_9222_) );
NOR2X1 NOR2X1_1462 ( .gnd(gnd), .vdd(vdd), .A(_9222_), .B(_8800__bF_buf8), .Y(_8699__154_) );
INVX2 INVX2_339 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_83_), .Y(_9223_) );
OAI21X1 OAI21X1_2601 ( .gnd(gnd), .vdd(vdd), .A(_9223_), .B(micro_hash_ucr_3_Wx_43_), .C(_9080_), .Y(_9224_) );
AOI21X1 AOI21X1_1642 ( .gnd(gnd), .vdd(vdd), .A(_9223_), .B(micro_hash_ucr_3_Wx_43_), .C(_9224_), .Y(_9225_) );
NOR2X1 NOR2X1_1463 ( .gnd(gnd), .vdd(vdd), .A(_9225_), .B(_8800__bF_buf7), .Y(_8699__155_) );
INVX2 INVX2_340 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_84_), .Y(_9226_) );
OAI21X1 OAI21X1_2602 ( .gnd(gnd), .vdd(vdd), .A(_9226_), .B(micro_hash_ucr_3_Wx_44_), .C(_9084_), .Y(_9227_) );
AOI21X1 AOI21X1_1643 ( .gnd(gnd), .vdd(vdd), .A(_9226_), .B(micro_hash_ucr_3_Wx_44_), .C(_9227_), .Y(_9228_) );
NOR2X1 NOR2X1_1464 ( .gnd(gnd), .vdd(vdd), .A(_9228_), .B(_8800__bF_buf6), .Y(_8699__156_) );
INVX2 INVX2_341 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_85_), .Y(_9229_) );
OAI21X1 OAI21X1_2603 ( .gnd(gnd), .vdd(vdd), .A(_9229_), .B(micro_hash_ucr_3_Wx_45_), .C(_9088_), .Y(_9230_) );
AOI21X1 AOI21X1_1644 ( .gnd(gnd), .vdd(vdd), .A(_9229_), .B(micro_hash_ucr_3_Wx_45_), .C(_9230_), .Y(_9231_) );
NOR2X1 NOR2X1_1465 ( .gnd(gnd), .vdd(vdd), .A(_9231_), .B(_8800__bF_buf5), .Y(_8699__157_) );
INVX4 INVX4_138 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_86_), .Y(_9232_) );
OAI21X1 OAI21X1_2604 ( .gnd(gnd), .vdd(vdd), .A(_9232_), .B(micro_hash_ucr_3_Wx_46_), .C(_9092_), .Y(_9233_) );
AOI21X1 AOI21X1_1645 ( .gnd(gnd), .vdd(vdd), .A(_9232_), .B(micro_hash_ucr_3_Wx_46_), .C(_9233_), .Y(_9234_) );
NOR2X1 NOR2X1_1466 ( .gnd(gnd), .vdd(vdd), .A(_9234_), .B(_8800__bF_buf4), .Y(_8699__158_) );
AOI21X1 AOI21X1_1646 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_47_), .B(_9037_), .C(micro_hash_ucr_3_Wx_135_), .Y(_9235_) );
OAI21X1 OAI21X1_2605 ( .gnd(gnd), .vdd(vdd), .A(_9037_), .B(micro_hash_ucr_3_Wx_47_), .C(_9235_), .Y(_9236_) );
AND2X2 AND2X2_542 ( .gnd(gnd), .vdd(vdd), .A(_9236_), .B(_8705__bF_buf0), .Y(_8699__159_) );
AND2X2 AND2X2_543 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf13), .B(concatenador_3_data_out_120_), .Y(_8699__120_) );
AND2X2 AND2X2_544 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf12), .B(concatenador_3_data_out_121_), .Y(_8699__121_) );
AND2X2 AND2X2_545 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf11), .B(concatenador_3_data_out_122_), .Y(_8699__122_) );
AND2X2 AND2X2_546 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf10), .B(concatenador_3_data_out_123_), .Y(_8699__123_) );
AND2X2 AND2X2_547 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf9), .B(concatenador_3_data_out_124_), .Y(_8699__124_) );
AND2X2 AND2X2_548 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf8), .B(concatenador_3_data_out_125_), .Y(_8699__125_) );
AND2X2 AND2X2_549 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf7), .B(concatenador_3_data_out_126_), .Y(_8699__126_) );
AND2X2 AND2X2_550 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf6), .B(concatenador_3_data_out_127_), .Y(_8699__127_) );
INVX2 INVX2_342 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_64_), .Y(_9237_) );
OAI21X1 OAI21X1_2606 ( .gnd(gnd), .vdd(vdd), .A(_9237_), .B(micro_hash_ucr_3_Wx_24_), .C(_9114_), .Y(_9238_) );
AOI21X1 AOI21X1_1647 ( .gnd(gnd), .vdd(vdd), .A(_9237_), .B(micro_hash_ucr_3_Wx_24_), .C(_9238_), .Y(_9239_) );
NOR2X1 NOR2X1_1467 ( .gnd(gnd), .vdd(vdd), .A(_9239_), .B(_8800__bF_buf3), .Y(_8699__136_) );
INVX2 INVX2_343 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_65_), .Y(_9240_) );
OAI21X1 OAI21X1_2607 ( .gnd(gnd), .vdd(vdd), .A(_9240_), .B(micro_hash_ucr_3_Wx_25_), .C(_9117_), .Y(_9241_) );
AOI21X1 AOI21X1_1648 ( .gnd(gnd), .vdd(vdd), .A(_9240_), .B(micro_hash_ucr_3_Wx_25_), .C(_9241_), .Y(_9242_) );
NOR2X1 NOR2X1_1468 ( .gnd(gnd), .vdd(vdd), .A(_9242_), .B(_8800__bF_buf2), .Y(_8699__137_) );
INVX2 INVX2_344 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_66_), .Y(_9243_) );
OAI21X1 OAI21X1_2608 ( .gnd(gnd), .vdd(vdd), .A(_9243_), .B(micro_hash_ucr_3_Wx_26_), .C(_9120_), .Y(_9244_) );
AOI21X1 AOI21X1_1649 ( .gnd(gnd), .vdd(vdd), .A(_9243_), .B(micro_hash_ucr_3_Wx_26_), .C(_9244_), .Y(_9245_) );
NOR2X1 NOR2X1_1469 ( .gnd(gnd), .vdd(vdd), .A(_9245_), .B(_8800__bF_buf1), .Y(_8699__138_) );
INVX2 INVX2_345 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_67_), .Y(_9246_) );
OAI21X1 OAI21X1_2609 ( .gnd(gnd), .vdd(vdd), .A(_9246_), .B(micro_hash_ucr_3_Wx_27_), .C(_9123_), .Y(_9247_) );
AOI21X1 AOI21X1_1650 ( .gnd(gnd), .vdd(vdd), .A(_9246_), .B(micro_hash_ucr_3_Wx_27_), .C(_9247_), .Y(_9248_) );
NOR2X1 NOR2X1_1470 ( .gnd(gnd), .vdd(vdd), .A(_9248_), .B(_8800__bF_buf0), .Y(_8699__139_) );
OAI21X1 OAI21X1_2610 ( .gnd(gnd), .vdd(vdd), .A(_9148_), .B(micro_hash_ucr_3_Wx_28_), .C(_9126_), .Y(_9249_) );
AOI21X1 AOI21X1_1651 ( .gnd(gnd), .vdd(vdd), .A(_9148_), .B(micro_hash_ucr_3_Wx_28_), .C(_9249_), .Y(_9250_) );
NOR2X1 NOR2X1_1471 ( .gnd(gnd), .vdd(vdd), .A(_9250_), .B(_8800__bF_buf12), .Y(_8699__140_) );
INVX2 INVX2_346 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_69_), .Y(_9251_) );
OAI21X1 OAI21X1_2611 ( .gnd(gnd), .vdd(vdd), .A(_9251_), .B(micro_hash_ucr_3_Wx_29_), .C(_9129_), .Y(_9252_) );
AOI21X1 AOI21X1_1652 ( .gnd(gnd), .vdd(vdd), .A(_9251_), .B(micro_hash_ucr_3_Wx_29_), .C(_9252_), .Y(_9253_) );
NOR2X1 NOR2X1_1472 ( .gnd(gnd), .vdd(vdd), .A(_9253_), .B(_8800__bF_buf11), .Y(_8699__141_) );
INVX1 INVX1_624 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_70_), .Y(_9254_) );
OAI21X1 OAI21X1_2612 ( .gnd(gnd), .vdd(vdd), .A(_9254_), .B(micro_hash_ucr_3_Wx_30_), .C(_9132_), .Y(_9255_) );
AOI21X1 AOI21X1_1653 ( .gnd(gnd), .vdd(vdd), .A(_9254_), .B(micro_hash_ucr_3_Wx_30_), .C(_9255_), .Y(_9256_) );
NOR2X1 NOR2X1_1473 ( .gnd(gnd), .vdd(vdd), .A(_9256_), .B(_8800__bF_buf10), .Y(_8699__142_) );
INVX2 INVX2_347 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_71_), .Y(_9257_) );
AOI21X1 AOI21X1_1654 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_31_), .B(_9257_), .C(micro_hash_ucr_3_Wx_119_), .Y(_9258_) );
OAI21X1 OAI21X1_2613 ( .gnd(gnd), .vdd(vdd), .A(_9257_), .B(micro_hash_ucr_3_Wx_31_), .C(_9258_), .Y(_9259_) );
AND2X2 AND2X2_551 ( .gnd(gnd), .vdd(vdd), .A(_9259_), .B(_8705__bF_buf5), .Y(_8699__143_) );
INVX2 INVX2_348 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_56_), .Y(_9260_) );
AOI21X1 AOI21X1_1655 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_16_), .B(_9260_), .C(micro_hash_ucr_3_Wx_104_), .Y(_9261_) );
OAI21X1 OAI21X1_2614 ( .gnd(gnd), .vdd(vdd), .A(_9260_), .B(micro_hash_ucr_3_Wx_16_), .C(_9261_), .Y(_9262_) );
AND2X2 AND2X2_552 ( .gnd(gnd), .vdd(vdd), .A(_9262_), .B(_8705__bF_buf4), .Y(_8699__128_) );
INVX2 INVX2_349 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_57_), .Y(_9263_) );
OAI21X1 OAI21X1_2615 ( .gnd(gnd), .vdd(vdd), .A(_9263_), .B(micro_hash_ucr_3_Wx_17_), .C(_9139_), .Y(_9264_) );
AOI21X1 AOI21X1_1656 ( .gnd(gnd), .vdd(vdd), .A(_9263_), .B(micro_hash_ucr_3_Wx_17_), .C(_9264_), .Y(_9265_) );
NOR2X1 NOR2X1_1474 ( .gnd(gnd), .vdd(vdd), .A(_9265_), .B(_8800__bF_buf9), .Y(_8699__129_) );
INVX2 INVX2_350 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_58_), .Y(_9266_) );
OAI21X1 OAI21X1_2616 ( .gnd(gnd), .vdd(vdd), .A(_9266_), .B(micro_hash_ucr_3_Wx_18_), .C(_9142_), .Y(_9267_) );
AOI21X1 AOI21X1_1657 ( .gnd(gnd), .vdd(vdd), .A(_9266_), .B(micro_hash_ucr_3_Wx_18_), .C(_9267_), .Y(_9268_) );
NOR2X1 NOR2X1_1475 ( .gnd(gnd), .vdd(vdd), .A(_9268_), .B(_8800__bF_buf8), .Y(_8699__130_) );
INVX2 INVX2_351 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_59_), .Y(_9269_) );
OAI21X1 OAI21X1_2617 ( .gnd(gnd), .vdd(vdd), .A(_9269_), .B(micro_hash_ucr_3_Wx_19_), .C(_9145_), .Y(_9270_) );
AOI21X1 AOI21X1_1658 ( .gnd(gnd), .vdd(vdd), .A(_9269_), .B(micro_hash_ucr_3_Wx_19_), .C(_9270_), .Y(_9271_) );
NOR2X1 NOR2X1_1476 ( .gnd(gnd), .vdd(vdd), .A(_9271_), .B(_8800__bF_buf7), .Y(_8699__131_) );
INVX2 INVX2_352 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_60_), .Y(_9272_) );
AOI21X1 AOI21X1_1659 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_20_), .B(_9272_), .C(micro_hash_ucr_3_Wx_108_), .Y(_9273_) );
OAI21X1 OAI21X1_2618 ( .gnd(gnd), .vdd(vdd), .A(_9272_), .B(micro_hash_ucr_3_Wx_20_), .C(_9273_), .Y(_9274_) );
AND2X2 AND2X2_553 ( .gnd(gnd), .vdd(vdd), .A(_9274_), .B(_8705__bF_buf3), .Y(_8699__132_) );
INVX2 INVX2_353 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_61_), .Y(_9275_) );
OAI21X1 OAI21X1_2619 ( .gnd(gnd), .vdd(vdd), .A(_9275_), .B(micro_hash_ucr_3_Wx_21_), .C(_9151_), .Y(_9276_) );
AOI21X1 AOI21X1_1660 ( .gnd(gnd), .vdd(vdd), .A(_9275_), .B(micro_hash_ucr_3_Wx_21_), .C(_9276_), .Y(_9277_) );
NOR2X1 NOR2X1_1477 ( .gnd(gnd), .vdd(vdd), .A(_9277_), .B(_8800__bF_buf6), .Y(_8699__133_) );
INVX4 INVX4_139 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_62_), .Y(_9278_) );
OAI21X1 OAI21X1_2620 ( .gnd(gnd), .vdd(vdd), .A(_9278_), .B(micro_hash_ucr_3_Wx_22_), .C(_9154_), .Y(_9279_) );
AOI21X1 AOI21X1_1661 ( .gnd(gnd), .vdd(vdd), .A(_9278_), .B(micro_hash_ucr_3_Wx_22_), .C(_9279_), .Y(_9280_) );
NOR2X1 NOR2X1_1478 ( .gnd(gnd), .vdd(vdd), .A(_9280_), .B(_8800__bF_buf5), .Y(_8699__134_) );
XNOR2X1 XNOR2X1_390 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_63_), .B(micro_hash_ucr_3_Wx_23_), .Y(_9281_) );
AOI21X1 AOI21X1_1662 ( .gnd(gnd), .vdd(vdd), .A(_8959_), .B(_9281_), .C(_8800__bF_buf4), .Y(_8699__135_) );
AND2X2 AND2X2_554 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf2), .B(concatenador_3_data_out_96_), .Y(_8699__96_) );
AND2X2 AND2X2_555 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf1), .B(concatenador_3_data_out_97_), .Y(_8699__97_) );
AND2X2 AND2X2_556 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf0), .B(concatenador_3_data_out_98_), .Y(_8699__98_) );
AND2X2 AND2X2_557 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf13), .B(concatenador_3_data_out_99_), .Y(_8699__99_) );
AND2X2 AND2X2_558 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf12), .B(concatenador_3_data_out_100_), .Y(_8699__100_) );
AND2X2 AND2X2_559 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf11), .B(concatenador_3_data_out_101_), .Y(_8699__101_) );
AND2X2 AND2X2_560 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf10), .B(concatenador_3_data_out_102_), .Y(_8699__102_) );
AND2X2 AND2X2_561 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf9), .B(concatenador_3_data_out_103_), .Y(_8699__103_) );
AND2X2 AND2X2_562 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf8), .B(concatenador_3_data_out_112_), .Y(_8699__112_) );
AND2X2 AND2X2_563 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf7), .B(concatenador_3_data_out_113_), .Y(_8699__113_) );
AND2X2 AND2X2_564 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf6), .B(concatenador_3_data_out_114_), .Y(_8699__114_) );
AND2X2 AND2X2_565 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf5), .B(concatenador_3_data_out_115_), .Y(_8699__115_) );
AND2X2 AND2X2_566 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf4), .B(concatenador_3_data_out_116_), .Y(_8699__116_) );
AND2X2 AND2X2_567 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf3), .B(concatenador_3_data_out_117_), .Y(_8699__117_) );
AND2X2 AND2X2_568 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf2), .B(concatenador_3_data_out_118_), .Y(_8699__118_) );
AND2X2 AND2X2_569 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf1), .B(concatenador_3_data_out_119_), .Y(_8699__119_) );
AND2X2 AND2X2_570 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf0), .B(concatenador_3_data_out_104_), .Y(_8699__104_) );
AND2X2 AND2X2_571 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf13), .B(concatenador_3_data_out_105_), .Y(_8699__105_) );
AND2X2 AND2X2_572 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf12), .B(concatenador_3_data_out_106_), .Y(_8699__106_) );
AND2X2 AND2X2_573 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf11), .B(concatenador_3_data_out_107_), .Y(_8699__107_) );
AND2X2 AND2X2_574 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf10), .B(concatenador_3_data_out_108_), .Y(_8699__108_) );
AND2X2 AND2X2_575 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf9), .B(concatenador_3_data_out_109_), .Y(_8699__109_) );
AND2X2 AND2X2_576 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf8), .B(concatenador_3_data_out_110_), .Y(_8699__110_) );
AND2X2 AND2X2_577 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf7), .B(concatenador_3_data_out_111_), .Y(_8699__111_) );
AND2X2 AND2X2_578 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf6), .B(concatenador_3_data_out_72_), .Y(_8699__72_) );
AND2X2 AND2X2_579 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf5), .B(concatenador_3_data_out_73_), .Y(_8699__73_) );
AND2X2 AND2X2_580 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf4), .B(concatenador_3_data_out_74_), .Y(_8699__74_) );
AND2X2 AND2X2_581 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf3), .B(concatenador_3_data_out_75_), .Y(_8699__75_) );
AND2X2 AND2X2_582 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf2), .B(concatenador_3_data_out_76_), .Y(_8699__76_) );
AND2X2 AND2X2_583 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf1), .B(concatenador_3_data_out_77_), .Y(_8699__77_) );
AND2X2 AND2X2_584 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf0), .B(concatenador_3_data_out_78_), .Y(_8699__78_) );
AND2X2 AND2X2_585 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf13), .B(concatenador_3_data_out_79_), .Y(_8699__79_) );
AND2X2 AND2X2_586 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf12), .B(concatenador_3_data_out_88_), .Y(_8699__88_) );
AND2X2 AND2X2_587 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf11), .B(concatenador_3_data_out_89_), .Y(_8699__89_) );
AND2X2 AND2X2_588 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf10), .B(concatenador_3_data_out_90_), .Y(_8699__90_) );
AND2X2 AND2X2_589 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf9), .B(concatenador_3_data_out_91_), .Y(_8699__91_) );
AND2X2 AND2X2_590 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf8), .B(concatenador_3_data_out_92_), .Y(_8699__92_) );
AND2X2 AND2X2_591 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf7), .B(concatenador_3_data_out_93_), .Y(_8699__93_) );
AND2X2 AND2X2_592 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf6), .B(concatenador_3_data_out_94_), .Y(_8699__94_) );
AND2X2 AND2X2_593 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf5), .B(concatenador_3_data_out_95_), .Y(_8699__95_) );
AND2X2 AND2X2_594 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf4), .B(concatenador_3_data_out_80_), .Y(_8699__80_) );
AND2X2 AND2X2_595 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf3), .B(concatenador_3_data_out_81_), .Y(_8699__81_) );
AND2X2 AND2X2_596 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf2), .B(concatenador_3_data_out_82_), .Y(_8699__82_) );
AND2X2 AND2X2_597 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf1), .B(concatenador_3_data_out_83_), .Y(_8699__83_) );
AND2X2 AND2X2_598 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf0), .B(concatenador_3_data_out_84_), .Y(_8699__84_) );
AND2X2 AND2X2_599 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf13), .B(concatenador_3_data_out_85_), .Y(_8699__85_) );
AND2X2 AND2X2_600 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf12), .B(concatenador_3_data_out_86_), .Y(_8699__86_) );
AND2X2 AND2X2_601 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf11), .B(concatenador_3_data_out_87_), .Y(_8699__87_) );
AND2X2 AND2X2_602 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf10), .B(concatenador_3_data_out_48_), .Y(_8699__48_) );
AND2X2 AND2X2_603 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf9), .B(concatenador_3_data_out_49_), .Y(_8699__49_) );
AND2X2 AND2X2_604 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf8), .B(concatenador_3_data_out_50_), .Y(_8699__50_) );
AND2X2 AND2X2_605 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf7), .B(concatenador_3_data_out_51_), .Y(_8699__51_) );
AND2X2 AND2X2_606 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf6), .B(concatenador_3_data_out_52_), .Y(_8699__52_) );
AND2X2 AND2X2_607 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf5), .B(concatenador_3_data_out_53_), .Y(_8699__53_) );
AND2X2 AND2X2_608 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf4), .B(concatenador_3_data_out_54_), .Y(_8699__54_) );
AND2X2 AND2X2_609 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf3), .B(concatenador_3_data_out_55_), .Y(_8699__55_) );
AND2X2 AND2X2_610 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf2), .B(concatenador_3_data_out_64_), .Y(_8699__64_) );
AND2X2 AND2X2_611 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf1), .B(concatenador_3_data_out_65_), .Y(_8699__65_) );
AND2X2 AND2X2_612 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf0), .B(concatenador_3_data_out_66_), .Y(_8699__66_) );
AND2X2 AND2X2_613 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf13), .B(concatenador_3_data_out_67_), .Y(_8699__67_) );
AND2X2 AND2X2_614 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf12), .B(concatenador_3_data_out_68_), .Y(_8699__68_) );
AND2X2 AND2X2_615 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf11), .B(concatenador_3_data_out_69_), .Y(_8699__69_) );
AND2X2 AND2X2_616 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf10), .B(concatenador_3_data_out_70_), .Y(_8699__70_) );
AND2X2 AND2X2_617 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf9), .B(concatenador_3_data_out_71_), .Y(_8699__71_) );
AND2X2 AND2X2_618 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf8), .B(concatenador_3_data_out_56_), .Y(_8699__56_) );
AND2X2 AND2X2_619 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf7), .B(concatenador_3_data_out_57_), .Y(_8699__57_) );
AND2X2 AND2X2_620 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf6), .B(concatenador_3_data_out_58_), .Y(_8699__58_) );
AND2X2 AND2X2_621 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf5), .B(concatenador_3_data_out_59_), .Y(_8699__59_) );
AND2X2 AND2X2_622 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf4), .B(concatenador_3_data_out_60_), .Y(_8699__60_) );
AND2X2 AND2X2_623 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf3), .B(concatenador_3_data_out_61_), .Y(_8699__61_) );
AND2X2 AND2X2_624 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf2), .B(concatenador_3_data_out_62_), .Y(_8699__62_) );
AND2X2 AND2X2_625 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf1), .B(concatenador_3_data_out_63_), .Y(_8699__63_) );
AND2X2 AND2X2_626 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf0), .B(concatenador_3_data_out_24_), .Y(_8699__24_) );
AND2X2 AND2X2_627 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf13), .B(concatenador_3_data_out_25_), .Y(_8699__25_) );
AND2X2 AND2X2_628 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf12), .B(concatenador_3_data_out_26_), .Y(_8699__26_) );
AND2X2 AND2X2_629 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf11), .B(concatenador_3_data_out_27_), .Y(_8699__27_) );
AND2X2 AND2X2_630 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf10), .B(concatenador_3_data_out_28_), .Y(_8699__28_) );
AND2X2 AND2X2_631 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf9), .B(concatenador_3_data_out_29_), .Y(_8699__29_) );
AND2X2 AND2X2_632 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf8), .B(concatenador_3_data_out_30_), .Y(_8699__30_) );
AND2X2 AND2X2_633 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf7), .B(concatenador_3_data_out_31_), .Y(_8699__31_) );
AND2X2 AND2X2_634 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf6), .B(concatenador_3_data_out_40_), .Y(_8699__40_) );
AND2X2 AND2X2_635 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf5), .B(concatenador_3_data_out_41_), .Y(_8699__41_) );
AND2X2 AND2X2_636 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf4), .B(concatenador_3_data_out_42_), .Y(_8699__42_) );
AND2X2 AND2X2_637 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf3), .B(concatenador_3_data_out_43_), .Y(_8699__43_) );
AND2X2 AND2X2_638 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf2), .B(concatenador_3_data_out_44_), .Y(_8699__44_) );
AND2X2 AND2X2_639 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf1), .B(concatenador_3_data_out_45_), .Y(_8699__45_) );
AND2X2 AND2X2_640 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf0), .B(concatenador_3_data_out_46_), .Y(_8699__46_) );
AND2X2 AND2X2_641 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf13), .B(concatenador_3_data_out_47_), .Y(_8699__47_) );
AND2X2 AND2X2_642 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf12), .B(concatenador_3_data_out_32_), .Y(_8699__32_) );
AND2X2 AND2X2_643 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf11), .B(concatenador_3_data_out_33_), .Y(_8699__33_) );
AND2X2 AND2X2_644 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf10), .B(concatenador_3_data_out_34_), .Y(_8699__34_) );
AND2X2 AND2X2_645 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf9), .B(concatenador_3_data_out_35_), .Y(_8699__35_) );
AND2X2 AND2X2_646 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf8), .B(concatenador_3_data_out_36_), .Y(_8699__36_) );
AND2X2 AND2X2_647 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf7), .B(concatenador_3_data_out_37_), .Y(_8699__37_) );
AND2X2 AND2X2_648 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf6), .B(concatenador_3_data_out_38_), .Y(_8699__38_) );
AND2X2 AND2X2_649 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf5), .B(concatenador_3_data_out_39_), .Y(_8699__39_) );
AND2X2 AND2X2_650 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf4), .B(concatenador_3_data_out_0_), .Y(_8699__0_) );
AND2X2 AND2X2_651 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf3), .B(concatenador_3_data_out_1_), .Y(_8699__1_) );
AND2X2 AND2X2_652 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf2), .B(concatenador_3_data_out_2_), .Y(_8699__2_) );
AND2X2 AND2X2_653 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf1), .B(concatenador_3_data_out_3_), .Y(_8699__3_) );
AND2X2 AND2X2_654 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf0), .B(concatenador_3_data_out_4_), .Y(_8699__4_) );
AND2X2 AND2X2_655 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf13), .B(concatenador_3_data_out_5_), .Y(_8699__5_) );
AND2X2 AND2X2_656 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf12), .B(concatenador_3_data_out_6_), .Y(_8699__6_) );
AND2X2 AND2X2_657 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf11), .B(concatenador_3_data_out_7_), .Y(_8699__7_) );
AND2X2 AND2X2_658 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf10), .B(concatenador_3_data_out_16_), .Y(_8699__16_) );
AND2X2 AND2X2_659 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf9), .B(concatenador_3_data_out_17_), .Y(_8699__17_) );
AND2X2 AND2X2_660 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf8), .B(concatenador_3_data_out_18_), .Y(_8699__18_) );
AND2X2 AND2X2_661 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf7), .B(concatenador_3_data_out_19_), .Y(_8699__19_) );
AND2X2 AND2X2_662 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf6), .B(concatenador_3_data_out_20_), .Y(_8699__20_) );
AND2X2 AND2X2_663 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf5), .B(concatenador_3_data_out_21_), .Y(_8699__21_) );
AND2X2 AND2X2_664 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf4), .B(concatenador_3_data_out_22_), .Y(_8699__22_) );
AND2X2 AND2X2_665 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf3), .B(concatenador_3_data_out_23_), .Y(_8699__23_) );
AND2X2 AND2X2_666 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf2), .B(concatenador_3_data_out_8_), .Y(_8699__8_) );
AND2X2 AND2X2_667 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf1), .B(concatenador_3_data_out_9_), .Y(_8699__9_) );
AND2X2 AND2X2_668 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf0), .B(concatenador_3_data_out_10_), .Y(_8699__10_) );
AND2X2 AND2X2_669 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf13), .B(concatenador_3_data_out_11_), .Y(_8699__11_) );
AND2X2 AND2X2_670 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf12), .B(concatenador_3_data_out_12_), .Y(_8699__12_) );
AND2X2 AND2X2_671 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf11), .B(concatenador_3_data_out_13_), .Y(_8699__13_) );
AND2X2 AND2X2_672 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf10), .B(concatenador_3_data_out_14_), .Y(_8699__14_) );
AND2X2 AND2X2_673 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf9), .B(concatenador_3_data_out_15_), .Y(_8699__15_) );
INVX8 INVX8_210 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe68_bF_buf3), .Y(_9282_) );
NOR2X1 NOR2X1_1479 ( .gnd(gnd), .vdd(vdd), .A(_9282__bF_buf4), .B(_8800__bF_buf3), .Y(_8770_) );
NOR2X1 NOR2X1_1480 ( .gnd(gnd), .vdd(vdd), .A(_12900__bF_buf1), .B(_8800__bF_buf2), .Y(_8773_) );
INVX8 INVX8_211 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe69), .Y(_9283_) );
NOR2X1 NOR2X1_1481 ( .gnd(gnd), .vdd(vdd), .A(_9283__bF_buf3), .B(_8800__bF_buf1), .Y(_8772_) );
INVX8 INVX8_212 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe65_bF_buf3), .Y(_9284_) );
NOR2X1 NOR2X1_1482 ( .gnd(gnd), .vdd(vdd), .A(_9284_), .B(_8800__bF_buf0), .Y(_8767_) );
INVX8 INVX8_213 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe67), .Y(_9285_) );
NOR2X1 NOR2X1_1483 ( .gnd(gnd), .vdd(vdd), .A(_9285__bF_buf3), .B(_8800__bF_buf12), .Y(_8769_) );
INVX8 INVX8_214 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe66_bF_buf4), .Y(_9286_) );
NOR2X1 NOR2X1_1484 ( .gnd(gnd), .vdd(vdd), .A(_9286__bF_buf3), .B(_8800__bF_buf11), .Y(_8768_) );
INVX8 INVX8_215 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe62_bF_buf3), .Y(_9287_) );
NOR2X1 NOR2X1_1485 ( .gnd(gnd), .vdd(vdd), .A(_9287__bF_buf4), .B(_8800__bF_buf10), .Y(_8764_) );
INVX8 INVX8_216 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe64_bF_buf4), .Y(_9288_) );
NOR2X1 NOR2X1_1486 ( .gnd(gnd), .vdd(vdd), .A(_9288__bF_buf3), .B(_8800__bF_buf9), .Y(_8766_) );
INVX8 INVX8_217 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe63), .Y(_9289_) );
NOR2X1 NOR2X1_1487 ( .gnd(gnd), .vdd(vdd), .A(_9289__bF_buf3), .B(_8800__bF_buf8), .Y(_8765_) );
INVX8 INVX8_218 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe59), .Y(_9290_) );
NOR2X1 NOR2X1_1488 ( .gnd(gnd), .vdd(vdd), .A(_9290__bF_buf3), .B(_8800__bF_buf7), .Y(_8761_) );
INVX8 INVX8_219 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe61_bF_buf3), .Y(_9291_) );
NOR2X1 NOR2X1_1489 ( .gnd(gnd), .vdd(vdd), .A(_9291_), .B(_8800__bF_buf6), .Y(_8763_) );
INVX8 INVX8_220 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe60_bF_buf4), .Y(_9292_) );
NOR2X1 NOR2X1_1490 ( .gnd(gnd), .vdd(vdd), .A(_9292__bF_buf3), .B(_8800__bF_buf5), .Y(_8762_) );
INVX8 INVX8_221 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe56_bF_buf4), .Y(_9293_) );
NOR2X1 NOR2X1_1491 ( .gnd(gnd), .vdd(vdd), .A(_9293__bF_buf3), .B(_8800__bF_buf4), .Y(_8757_) );
INVX8 INVX8_222 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe58_bF_buf3), .Y(_9294_) );
NOR2X1 NOR2X1_1492 ( .gnd(gnd), .vdd(vdd), .A(_9294__bF_buf4), .B(_8800__bF_buf3), .Y(_8759_) );
INVX8 INVX8_223 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe57_bF_buf3), .Y(_9295_) );
NOR2X1 NOR2X1_1493 ( .gnd(gnd), .vdd(vdd), .A(_9295_), .B(_8800__bF_buf2), .Y(_8758_) );
INVX8 INVX8_224 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe53), .Y(_9296_) );
NOR2X1 NOR2X1_1494 ( .gnd(gnd), .vdd(vdd), .A(_9296_), .B(_8800__bF_buf1), .Y(_8754_) );
INVX8 INVX8_225 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe55), .Y(_9297_) );
NOR2X1 NOR2X1_1495 ( .gnd(gnd), .vdd(vdd), .A(_9297_), .B(_8800__bF_buf0), .Y(_8756_) );
INVX8 INVX8_226 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe54_bF_buf3), .Y(_9298_) );
NOR2X1 NOR2X1_1496 ( .gnd(gnd), .vdd(vdd), .A(_9298__bF_buf4), .B(_8800__bF_buf12), .Y(_8755_) );
INVX8 INVX8_227 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe50_bF_buf4), .Y(_9299_) );
NOR2X1 NOR2X1_1497 ( .gnd(gnd), .vdd(vdd), .A(_9299__bF_buf3), .B(_8800__bF_buf11), .Y(_8751_) );
INVX8 INVX8_228 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe52_bF_buf4), .Y(_9300_) );
NOR2X1 NOR2X1_1498 ( .gnd(gnd), .vdd(vdd), .A(_9300__bF_buf3), .B(_8800__bF_buf10), .Y(_8753_) );
INVX8 INVX8_229 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe51), .Y(_9301_) );
NOR2X1 NOR2X1_1499 ( .gnd(gnd), .vdd(vdd), .A(_9301__bF_buf3), .B(_8800__bF_buf9), .Y(_8752_) );
INVX8 INVX8_230 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe47), .Y(_9302_) );
NOR2X1 NOR2X1_1500 ( .gnd(gnd), .vdd(vdd), .A(_9302_), .B(_8800__bF_buf8), .Y(_8747_) );
INVX4 INVX4_140 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe49_bF_buf3), .Y(_9303_) );
NOR2X1 NOR2X1_1501 ( .gnd(gnd), .vdd(vdd), .A(_9303_), .B(_8800__bF_buf7), .Y(_8750_) );
INVX8 INVX8_231 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe48_bF_buf4), .Y(_9304_) );
NOR2X1 NOR2X1_1502 ( .gnd(gnd), .vdd(vdd), .A(_9304__bF_buf3), .B(_8800__bF_buf6), .Y(_8748_) );
INVX8 INVX8_232 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe44_bF_buf3), .Y(_9305_) );
NOR2X1 NOR2X1_1503 ( .gnd(gnd), .vdd(vdd), .A(_9305__bF_buf4), .B(_8800__bF_buf5), .Y(_8744_) );
INVX8 INVX8_233 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe46_bF_buf4), .Y(_9306_) );
NOR2X1 NOR2X1_1504 ( .gnd(gnd), .vdd(vdd), .A(_9306__bF_buf3), .B(_8800__bF_buf4), .Y(_8746_) );
INVX8 INVX8_234 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe45_bF_buf3), .Y(_9307_) );
NOR2X1 NOR2X1_1505 ( .gnd(gnd), .vdd(vdd), .A(_9307_), .B(_8800__bF_buf3), .Y(_8745_) );
INVX8 INVX8_235 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe41_bF_buf3), .Y(_9308_) );
NOR2X1 NOR2X1_1506 ( .gnd(gnd), .vdd(vdd), .A(_9308_), .B(_8800__bF_buf2), .Y(_8741_) );
INVX8 INVX8_236 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe43), .Y(_9309_) );
NOR2X1 NOR2X1_1507 ( .gnd(gnd), .vdd(vdd), .A(_9309__bF_buf3), .B(_8800__bF_buf1), .Y(_8743_) );
INVX8 INVX8_237 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe42_bF_buf3), .Y(_9310_) );
NOR2X1 NOR2X1_1508 ( .gnd(gnd), .vdd(vdd), .A(_9310__bF_buf4), .B(_8800__bF_buf0), .Y(_8742_) );
INVX8 INVX8_238 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe38_bF_buf3), .Y(_9311_) );
NOR2X1 NOR2X1_1509 ( .gnd(gnd), .vdd(vdd), .A(_9311__bF_buf4), .B(_8800__bF_buf12), .Y(_8737_) );
INVX8 INVX8_239 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe40_bF_buf4), .Y(_9312_) );
NOR2X1 NOR2X1_1510 ( .gnd(gnd), .vdd(vdd), .A(_9312__bF_buf3), .B(_8800__bF_buf11), .Y(_8740_) );
INVX4 INVX4_141 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe39_bF_buf3), .Y(_9313_) );
NOR2X1 NOR2X1_1511 ( .gnd(gnd), .vdd(vdd), .A(_9313_), .B(_8800__bF_buf10), .Y(_8739_) );
INVX8 INVX8_240 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe35_bF_buf3), .Y(_9314_) );
NOR2X1 NOR2X1_1512 ( .gnd(gnd), .vdd(vdd), .A(_9314_), .B(_8800__bF_buf9), .Y(_8734_) );
INVX8 INVX8_241 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe37_bF_buf3), .Y(_9315_) );
NOR2X1 NOR2X1_1513 ( .gnd(gnd), .vdd(vdd), .A(_9315_), .B(_8800__bF_buf8), .Y(_8736_) );
INVX8 INVX8_242 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe36_bF_buf4), .Y(_9316_) );
NOR2X1 NOR2X1_1514 ( .gnd(gnd), .vdd(vdd), .A(_9316__bF_buf3), .B(_8800__bF_buf7), .Y(_8735_) );
INVX8 INVX8_243 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe32_bF_buf3), .Y(_9317_) );
NOR2X1 NOR2X1_1515 ( .gnd(gnd), .vdd(vdd), .A(_9317__bF_buf4), .B(_8800__bF_buf6), .Y(_8731_) );
INVX8 INVX8_244 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe34_bF_buf4), .Y(_9318_) );
NOR2X1 NOR2X1_1516 ( .gnd(gnd), .vdd(vdd), .A(_9318__bF_buf4), .B(_8800__bF_buf5), .Y(_8733_) );
INVX8 INVX8_245 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe33_bF_buf3), .Y(_9319_) );
NOR2X1 NOR2X1_1517 ( .gnd(gnd), .vdd(vdd), .A(_9319_), .B(_8800__bF_buf4), .Y(_8732_) );
INVX8 INVX8_246 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe29_bF_buf3), .Y(_9320_) );
NOR2X1 NOR2X1_1518 ( .gnd(gnd), .vdd(vdd), .A(_9320_), .B(_8800__bF_buf3), .Y(_8728_) );
INVX8 INVX8_247 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe31), .Y(_9321_) );
NOR2X1 NOR2X1_1519 ( .gnd(gnd), .vdd(vdd), .A(_9321__bF_buf3), .B(_8800__bF_buf2), .Y(_8730_) );
INVX8 INVX8_248 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe30_bF_buf4), .Y(_9322_) );
NOR2X1 NOR2X1_1520 ( .gnd(gnd), .vdd(vdd), .A(_9322__bF_buf3), .B(_8800__bF_buf1), .Y(_8729_) );
INVX8 INVX8_249 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe26_bF_buf4), .Y(_9323_) );
NOR2X1 NOR2X1_1521 ( .gnd(gnd), .vdd(vdd), .A(_9323__bF_buf3), .B(_8800__bF_buf0), .Y(_8724_) );
INVX8 INVX8_250 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe28_bF_buf4), .Y(_9324_) );
NOR2X1 NOR2X1_1522 ( .gnd(gnd), .vdd(vdd), .A(_9324__bF_buf4), .B(_8800__bF_buf12), .Y(_8726_) );
INVX8 INVX8_251 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe27), .Y(_9325_) );
NOR2X1 NOR2X1_1523 ( .gnd(gnd), .vdd(vdd), .A(_9325__bF_buf3), .B(_8800__bF_buf11), .Y(_8725_) );
INVX8 INVX8_252 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe23), .Y(_9326_) );
NOR2X1 NOR2X1_1524 ( .gnd(gnd), .vdd(vdd), .A(_9326__bF_buf3), .B(_8800__bF_buf10), .Y(_8721_) );
INVX8 INVX8_253 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe25_bF_buf3), .Y(_9327_) );
NOR2X1 NOR2X1_1525 ( .gnd(gnd), .vdd(vdd), .A(_9327_), .B(_8800__bF_buf9), .Y(_8723_) );
INVX8 INVX8_254 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe24_bF_buf4), .Y(_9328_) );
NOR2X1 NOR2X1_1526 ( .gnd(gnd), .vdd(vdd), .A(_9328__bF_buf3), .B(_8800__bF_buf8), .Y(_8722_) );
INVX8 INVX8_255 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe20_bF_buf4), .Y(_9329_) );
NOR2X1 NOR2X1_1527 ( .gnd(gnd), .vdd(vdd), .A(_9329__bF_buf4), .B(_8800__bF_buf7), .Y(_8718_) );
INVX8 INVX8_256 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe22_bF_buf4), .Y(_9330_) );
NOR2X1 NOR2X1_1528 ( .gnd(gnd), .vdd(vdd), .A(_9330__bF_buf4), .B(_8800__bF_buf6), .Y(_8720_) );
INVX8 INVX8_257 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe21_bF_buf3), .Y(_9331_) );
NOR2X1 NOR2X1_1529 ( .gnd(gnd), .vdd(vdd), .A(_9331_), .B(_8800__bF_buf5), .Y(_8719_) );
INVX4 INVX4_142 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe17_bF_buf3), .Y(_9332_) );
NOR2X1 NOR2X1_1530 ( .gnd(gnd), .vdd(vdd), .A(_9332_), .B(_8800__bF_buf4), .Y(_8714_) );
INVX8 INVX8_258 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe19), .Y(_9333_) );
NOR2X1 NOR2X1_1531 ( .gnd(gnd), .vdd(vdd), .A(_9333__bF_buf3), .B(_8800__bF_buf3), .Y(_8717_) );
INVX8 INVX8_259 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe18_bF_buf4), .Y(_9334_) );
NOR2X1 NOR2X1_1532 ( .gnd(gnd), .vdd(vdd), .A(_9334__bF_buf3), .B(_8800__bF_buf2), .Y(_8715_) );
INVX8 INVX8_260 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe14_bF_buf3), .Y(_9335_) );
NOR2X1 NOR2X1_1533 ( .gnd(gnd), .vdd(vdd), .A(_9335__bF_buf3), .B(_8800__bF_buf1), .Y(_8711_) );
INVX8 INVX8_261 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe16_bF_buf4), .Y(_9336_) );
NOR2X1 NOR2X1_1534 ( .gnd(gnd), .vdd(vdd), .A(_9336__bF_buf3), .B(_8800__bF_buf0), .Y(_8713_) );
INVX8 INVX8_262 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe15_bF_buf3), .Y(_9337_) );
NOR2X1 NOR2X1_1535 ( .gnd(gnd), .vdd(vdd), .A(_9337_), .B(_8800__bF_buf12), .Y(_8712_) );
INVX2 INVX2_354 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe11), .Y(_9338_) );
NOR2X1 NOR2X1_1536 ( .gnd(gnd), .vdd(vdd), .A(_9338_), .B(_8800__bF_buf11), .Y(_8708_) );
INVX4 INVX4_143 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe13), .Y(_9339_) );
NOR2X1 NOR2X1_1537 ( .gnd(gnd), .vdd(vdd), .A(_9339_), .B(_8800__bF_buf10), .Y(_8710_) );
INVX8 INVX8_263 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe12), .Y(_9340_) );
NOR2X1 NOR2X1_1538 ( .gnd(gnd), .vdd(vdd), .A(_9340_), .B(_8800__bF_buf9), .Y(_8709_) );
INVX8 INVX8_264 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe8), .Y(_9341_) );
NOR2X1 NOR2X1_1539 ( .gnd(gnd), .vdd(vdd), .A(_9341_), .B(_8800__bF_buf8), .Y(_8776_) );
INVX8 INVX8_265 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe10_bF_buf3), .Y(_9342_) );
NOR2X1 NOR2X1_1540 ( .gnd(gnd), .vdd(vdd), .A(_9342_), .B(_8800__bF_buf7), .Y(_8707_) );
INVX4 INVX4_144 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe9), .Y(_9343_) );
NOR2X1 NOR2X1_1541 ( .gnd(gnd), .vdd(vdd), .A(_9343_), .B(_8800__bF_buf6), .Y(_8706_) );
AND2X2 AND2X2_674 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf8), .B(micro_hash_ucr_3_pipe5), .Y(_8771_) );
INVX4 INVX4_145 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe7), .Y(_9344_) );
NOR2X1 NOR2X1_1542 ( .gnd(gnd), .vdd(vdd), .A(_9344_), .B(_8800__bF_buf5), .Y(_8775_) );
INVX4 INVX4_146 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe6_bF_buf3), .Y(_9345_) );
NOR2X1 NOR2X1_1543 ( .gnd(gnd), .vdd(vdd), .A(_9345_), .B(_8800__bF_buf4), .Y(_8774_) );
AND2X2 AND2X2_675 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf7), .B(micro_hash_ucr_3_pipe2), .Y(_8738_) );
AND2X2 AND2X2_676 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf6), .B(micro_hash_ucr_3_pipe4), .Y(_8760_) );
AND2X2 AND2X2_677 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf5), .B(micro_hash_ucr_3_pipe3), .Y(_8749_) );
AND2X2 AND2X2_678 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf4), .B(micro_hash_ucr_3_pipe1), .Y(_8727_) );
AND2X2 AND2X2_679 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf3), .B(micro_hash_ucr_3_pipe0), .Y(_8716_) );
NAND2X1 NAND2X1_1173 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe64_bF_buf3), .B(_8862__bF_buf2), .Y(_9346_) );
NAND2X1 NAND2X1_1174 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe62_bF_buf2), .B(_8862__bF_buf1), .Y(_9347_) );
NAND2X1 NAND2X1_1175 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe60_bF_buf3), .B(_8862__bF_buf0), .Y(_9348_) );
NAND2X1 NAND2X1_1176 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_0_bF_buf1_), .B(micro_hash_ucr_3_pipe54_bF_buf2), .Y(_9349_) );
NAND2X1 NAND2X1_1177 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_0_bF_buf0_), .B(micro_hash_ucr_3_pipe52_bF_buf3), .Y(_9350_) );
NAND2X1 NAND2X1_1178 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_0_bF_buf3_), .B(micro_hash_ucr_3_pipe50_bF_buf3), .Y(_9351_) );
NAND2X1 NAND2X1_1179 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_0_bF_buf2_), .B(micro_hash_ucr_3_pipe48_bF_buf3), .Y(_9352_) );
NAND2X1 NAND2X1_1180 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_0_bF_buf1_), .B(micro_hash_ucr_3_pipe38_bF_buf2), .Y(_9353_) );
NAND2X1 NAND2X1_1181 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_0_bF_buf0_), .B(micro_hash_ucr_3_pipe36_bF_buf3), .Y(_9354_) );
NAND2X1 NAND2X1_1182 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_0_bF_buf3_), .B(micro_hash_ucr_3_pipe30_bF_buf3), .Y(_9355_) );
NAND2X1 NAND2X1_1183 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_0_bF_buf2_), .B(micro_hash_ucr_3_pipe28_bF_buf3), .Y(_9356_) );
NAND2X1 NAND2X1_1184 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe22_bF_buf3), .B(_8862__bF_buf3), .Y(_9357_) );
NAND2X1 NAND2X1_1185 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe20_bF_buf3), .B(_8862__bF_buf2), .Y(_9358_) );
NAND2X1 NAND2X1_1186 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe18_bF_buf3), .B(_8862__bF_buf1), .Y(_9359_) );
NAND2X1 NAND2X1_1187 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe16_bF_buf3), .B(_8862__bF_buf0), .Y(_9360_) );
NOR2X1 NOR2X1_1544 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_0_), .B(micro_hash_ucr_3_b_0_bF_buf1_), .Y(_9361_) );
NOR2X1 NOR2X1_1545 ( .gnd(gnd), .vdd(vdd), .A(_12848__bF_buf1), .B(_12902_), .Y(_9362_) );
NOR2X1 NOR2X1_1546 ( .gnd(gnd), .vdd(vdd), .A(_9361_), .B(_9362_), .Y(_9363_) );
NAND2X1 NAND2X1_1188 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe15_bF_buf2), .B(_9363_), .Y(_9364_) );
NOR2X1 NOR2X1_1547 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe8), .B(micro_hash_ucr_3_pipe10_bF_buf2), .Y(_9365_) );
NOR2X1 NOR2X1_1548 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe11), .B(micro_hash_ucr_3_pipe13), .Y(_9366_) );
OAI21X1 OAI21X1_2621 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe10_bF_buf1), .B(_9343_), .C(_9366_), .Y(_9367_) );
AOI21X1 AOI21X1_1663 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe7), .B(_9365_), .C(_9367_), .Y(_9368_) );
NOR2X1 NOR2X1_1549 ( .gnd(gnd), .vdd(vdd), .A(_9363_), .B(_9368_), .Y(_9369_) );
OR2X2 OR2X2_66 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe7), .B(micro_hash_ucr_3_pipe6_bF_buf2), .Y(_9370_) );
AOI22X1 AOI22X1_64 ( .gnd(gnd), .vdd(vdd), .A(_9342_), .B(micro_hash_ucr_3_pipe9), .C(_9370_), .D(_9365_), .Y(_9371_) );
NAND2X1 NAND2X1_1189 ( .gnd(gnd), .vdd(vdd), .A(_9343_), .B(_9344_), .Y(_9372_) );
INVX2 INVX2_355 ( .gnd(gnd), .vdd(vdd), .A(_9372_), .Y(_9373_) );
OR2X2 OR2X2_67 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe8), .B(micro_hash_ucr_3_pipe10_bF_buf0), .Y(_9374_) );
NOR3X1 NOR3X1_7 ( .gnd(gnd), .vdd(vdd), .A(H_3_0_), .B(_9345_), .C(_9374_), .Y(_9375_) );
AOI22X1 AOI22X1_65 ( .gnd(gnd), .vdd(vdd), .A(_8862__bF_buf3), .B(_9371_), .C(_9375_), .D(_9373_), .Y(_9376_) );
OAI21X1 OAI21X1_2622 ( .gnd(gnd), .vdd(vdd), .A(_9376_), .B(micro_hash_ucr_3_pipe11), .C(_9340_), .Y(_9377_) );
AOI21X1 AOI21X1_1664 ( .gnd(gnd), .vdd(vdd), .A(_9339_), .B(_9377_), .C(_9369_), .Y(_9378_) );
NAND2X1 NAND2X1_1190 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe12), .B(_9339_), .Y(_9379_) );
OAI21X1 OAI21X1_2623 ( .gnd(gnd), .vdd(vdd), .A(_9379_), .B(_8862__bF_buf2), .C(_9335__bF_buf2), .Y(_9380_) );
AOI21X1 AOI21X1_1665 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe14_bF_buf2), .B(_8862__bF_buf1), .C(micro_hash_ucr_3_pipe15_bF_buf1), .Y(_9381_) );
OAI21X1 OAI21X1_2624 ( .gnd(gnd), .vdd(vdd), .A(_9378_), .B(_9380_), .C(_9381_), .Y(_9382_) );
NAND3X1 NAND3X1_417 ( .gnd(gnd), .vdd(vdd), .A(_9336__bF_buf2), .B(_9364_), .C(_9382_), .Y(_9383_) );
NAND3X1 NAND3X1_418 ( .gnd(gnd), .vdd(vdd), .A(_9332_), .B(_9360_), .C(_9383_), .Y(_9384_) );
NAND2X1 NAND2X1_1191 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe17_bF_buf2), .B(_9363_), .Y(_9385_) );
NAND3X1 NAND3X1_419 ( .gnd(gnd), .vdd(vdd), .A(_9334__bF_buf2), .B(_9385_), .C(_9384_), .Y(_9386_) );
NAND3X1 NAND3X1_420 ( .gnd(gnd), .vdd(vdd), .A(_9333__bF_buf2), .B(_9359_), .C(_9386_), .Y(_9387_) );
NAND2X1 NAND2X1_1192 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe19), .B(_9363_), .Y(_9388_) );
NAND3X1 NAND3X1_421 ( .gnd(gnd), .vdd(vdd), .A(_9329__bF_buf3), .B(_9388_), .C(_9387_), .Y(_9389_) );
NAND3X1 NAND3X1_422 ( .gnd(gnd), .vdd(vdd), .A(_9331_), .B(_9358_), .C(_9389_), .Y(_9390_) );
NAND2X1 NAND2X1_1193 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe21_bF_buf2), .B(_9363_), .Y(_9391_) );
NAND3X1 NAND3X1_423 ( .gnd(gnd), .vdd(vdd), .A(_9330__bF_buf3), .B(_9391_), .C(_9390_), .Y(_9392_) );
NAND3X1 NAND3X1_424 ( .gnd(gnd), .vdd(vdd), .A(_9326__bF_buf2), .B(_9357_), .C(_9392_), .Y(_9393_) );
NAND2X1 NAND2X1_1194 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe23), .B(_9363_), .Y(_9394_) );
AOI21X1 AOI21X1_1666 ( .gnd(gnd), .vdd(vdd), .A(_9394_), .B(_9393_), .C(micro_hash_ucr_3_pipe24_bF_buf3), .Y(_9395_) );
OAI21X1 OAI21X1_2625 ( .gnd(gnd), .vdd(vdd), .A(_8862__bF_buf0), .B(_9328__bF_buf2), .C(_9327_), .Y(_9396_) );
INVX4 INVX4_147 ( .gnd(gnd), .vdd(vdd), .A(_9363_), .Y(_9397_) );
AOI21X1 AOI21X1_1667 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe25_bF_buf2), .B(_9397_), .C(micro_hash_ucr_3_pipe26_bF_buf3), .Y(_9398_) );
OAI21X1 OAI21X1_2626 ( .gnd(gnd), .vdd(vdd), .A(_9395_), .B(_9396_), .C(_9398_), .Y(_9399_) );
NAND2X1 NAND2X1_1195 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_0_bF_buf1_), .B(micro_hash_ucr_3_pipe26_bF_buf2), .Y(_9400_) );
NAND3X1 NAND3X1_425 ( .gnd(gnd), .vdd(vdd), .A(_9325__bF_buf2), .B(_9400_), .C(_9399_), .Y(_9401_) );
OAI21X1 OAI21X1_2627 ( .gnd(gnd), .vdd(vdd), .A(_9362_), .B(_9361_), .C(micro_hash_ucr_3_pipe27), .Y(_9402_) );
NAND3X1 NAND3X1_426 ( .gnd(gnd), .vdd(vdd), .A(_9324__bF_buf3), .B(_9402_), .C(_9401_), .Y(_9403_) );
NAND3X1 NAND3X1_427 ( .gnd(gnd), .vdd(vdd), .A(_9320_), .B(_9356_), .C(_9403_), .Y(_9404_) );
OAI21X1 OAI21X1_2628 ( .gnd(gnd), .vdd(vdd), .A(_9362_), .B(_9361_), .C(micro_hash_ucr_3_pipe29_bF_buf2), .Y(_9405_) );
NAND3X1 NAND3X1_428 ( .gnd(gnd), .vdd(vdd), .A(_9322__bF_buf2), .B(_9405_), .C(_9404_), .Y(_9406_) );
AOI21X1 AOI21X1_1668 ( .gnd(gnd), .vdd(vdd), .A(_9355_), .B(_9406_), .C(micro_hash_ucr_3_pipe31), .Y(_9407_) );
OAI21X1 OAI21X1_2629 ( .gnd(gnd), .vdd(vdd), .A(_9397_), .B(_9321__bF_buf2), .C(_9317__bF_buf3), .Y(_9408_) );
AOI21X1 AOI21X1_1669 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe32_bF_buf2), .B(_8862__bF_buf3), .C(micro_hash_ucr_3_pipe33_bF_buf2), .Y(_9409_) );
OAI21X1 OAI21X1_2630 ( .gnd(gnd), .vdd(vdd), .A(_9407_), .B(_9408_), .C(_9409_), .Y(_9410_) );
AOI21X1 AOI21X1_1670 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe33_bF_buf1), .B(_9363_), .C(micro_hash_ucr_3_pipe34_bF_buf3), .Y(_9411_) );
NOR2X1 NOR2X1_1550 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_0_bF_buf0_), .B(_9318__bF_buf3), .Y(_9412_) );
AOI21X1 AOI21X1_1671 ( .gnd(gnd), .vdd(vdd), .A(_9411_), .B(_9410_), .C(_9412_), .Y(_9413_) );
OAI21X1 OAI21X1_2631 ( .gnd(gnd), .vdd(vdd), .A(_9362_), .B(_9361_), .C(micro_hash_ucr_3_pipe35_bF_buf2), .Y(_9414_) );
OAI21X1 OAI21X1_2632 ( .gnd(gnd), .vdd(vdd), .A(_9413_), .B(micro_hash_ucr_3_pipe35_bF_buf1), .C(_9414_), .Y(_9415_) );
OAI21X1 OAI21X1_2633 ( .gnd(gnd), .vdd(vdd), .A(_9415_), .B(micro_hash_ucr_3_pipe36_bF_buf2), .C(_9354_), .Y(_9416_) );
OAI21X1 OAI21X1_2634 ( .gnd(gnd), .vdd(vdd), .A(_9362_), .B(_9361_), .C(micro_hash_ucr_3_pipe37_bF_buf2), .Y(_9417_) );
OAI21X1 OAI21X1_2635 ( .gnd(gnd), .vdd(vdd), .A(_9416_), .B(micro_hash_ucr_3_pipe37_bF_buf1), .C(_9417_), .Y(_9418_) );
OAI21X1 OAI21X1_2636 ( .gnd(gnd), .vdd(vdd), .A(_9418_), .B(micro_hash_ucr_3_pipe38_bF_buf1), .C(_9353_), .Y(_9419_) );
OAI21X1 OAI21X1_2637 ( .gnd(gnd), .vdd(vdd), .A(_9362_), .B(_9361_), .C(micro_hash_ucr_3_pipe39_bF_buf2), .Y(_9420_) );
OAI21X1 OAI21X1_2638 ( .gnd(gnd), .vdd(vdd), .A(_9419_), .B(micro_hash_ucr_3_pipe39_bF_buf1), .C(_9420_), .Y(_9421_) );
AOI21X1 AOI21X1_1672 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_0_bF_buf3_), .B(micro_hash_ucr_3_pipe40_bF_buf3), .C(micro_hash_ucr_3_pipe41_bF_buf2), .Y(_9422_) );
OAI21X1 OAI21X1_2639 ( .gnd(gnd), .vdd(vdd), .A(_9421_), .B(micro_hash_ucr_3_pipe40_bF_buf2), .C(_9422_), .Y(_9423_) );
AOI21X1 AOI21X1_1673 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe41_bF_buf1), .B(_9397_), .C(micro_hash_ucr_3_pipe42_bF_buf2), .Y(_9424_) );
NOR2X1 NOR2X1_1551 ( .gnd(gnd), .vdd(vdd), .A(_8862__bF_buf2), .B(_9310__bF_buf3), .Y(_9425_) );
AOI21X1 AOI21X1_1674 ( .gnd(gnd), .vdd(vdd), .A(_9424_), .B(_9423_), .C(_9425_), .Y(_9426_) );
AOI21X1 AOI21X1_1675 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe43), .B(_9363_), .C(micro_hash_ucr_3_pipe44_bF_buf2), .Y(_9427_) );
OAI21X1 OAI21X1_2640 ( .gnd(gnd), .vdd(vdd), .A(_9426_), .B(micro_hash_ucr_3_pipe43), .C(_9427_), .Y(_9428_) );
AOI21X1 AOI21X1_1676 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe44_bF_buf1), .B(_8862__bF_buf1), .C(micro_hash_ucr_3_pipe45_bF_buf2), .Y(_9429_) );
OAI21X1 OAI21X1_2641 ( .gnd(gnd), .vdd(vdd), .A(_9397_), .B(_9307_), .C(_9306__bF_buf2), .Y(_9430_) );
AOI21X1 AOI21X1_1677 ( .gnd(gnd), .vdd(vdd), .A(_9429_), .B(_9428_), .C(_9430_), .Y(_9431_) );
NOR2X1 NOR2X1_1552 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_0_bF_buf2_), .B(_9306__bF_buf1), .Y(_9432_) );
OAI21X1 OAI21X1_2642 ( .gnd(gnd), .vdd(vdd), .A(_9431_), .B(_9432_), .C(_9302_), .Y(_9433_) );
OAI21X1 OAI21X1_2643 ( .gnd(gnd), .vdd(vdd), .A(_9362_), .B(_9361_), .C(micro_hash_ucr_3_pipe47), .Y(_9434_) );
NAND3X1 NAND3X1_429 ( .gnd(gnd), .vdd(vdd), .A(_9304__bF_buf2), .B(_9434_), .C(_9433_), .Y(_9435_) );
NAND3X1 NAND3X1_430 ( .gnd(gnd), .vdd(vdd), .A(_9303_), .B(_9352_), .C(_9435_), .Y(_9436_) );
OAI21X1 OAI21X1_2644 ( .gnd(gnd), .vdd(vdd), .A(_9362_), .B(_9361_), .C(micro_hash_ucr_3_pipe49_bF_buf2), .Y(_9437_) );
NAND3X1 NAND3X1_431 ( .gnd(gnd), .vdd(vdd), .A(_9299__bF_buf2), .B(_9437_), .C(_9436_), .Y(_9438_) );
NAND3X1 NAND3X1_432 ( .gnd(gnd), .vdd(vdd), .A(_9301__bF_buf2), .B(_9351_), .C(_9438_), .Y(_9439_) );
OAI21X1 OAI21X1_2645 ( .gnd(gnd), .vdd(vdd), .A(_9362_), .B(_9361_), .C(micro_hash_ucr_3_pipe51), .Y(_9440_) );
NAND3X1 NAND3X1_433 ( .gnd(gnd), .vdd(vdd), .A(_9300__bF_buf2), .B(_9440_), .C(_9439_), .Y(_9441_) );
NAND3X1 NAND3X1_434 ( .gnd(gnd), .vdd(vdd), .A(_9296_), .B(_9350_), .C(_9441_), .Y(_9442_) );
OAI21X1 OAI21X1_2646 ( .gnd(gnd), .vdd(vdd), .A(_9362_), .B(_9361_), .C(micro_hash_ucr_3_pipe53), .Y(_9443_) );
NAND3X1 NAND3X1_435 ( .gnd(gnd), .vdd(vdd), .A(_9298__bF_buf3), .B(_9443_), .C(_9442_), .Y(_9444_) );
NAND3X1 NAND3X1_436 ( .gnd(gnd), .vdd(vdd), .A(_9297_), .B(_9349_), .C(_9444_), .Y(_9445_) );
OAI21X1 OAI21X1_2647 ( .gnd(gnd), .vdd(vdd), .A(_9362_), .B(_9361_), .C(micro_hash_ucr_3_pipe55), .Y(_9446_) );
NAND3X1 NAND3X1_437 ( .gnd(gnd), .vdd(vdd), .A(_9293__bF_buf2), .B(_9446_), .C(_9445_), .Y(_9447_) );
AOI21X1 AOI21X1_1678 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_0_bF_buf1_), .B(micro_hash_ucr_3_pipe56_bF_buf3), .C(micro_hash_ucr_3_pipe57_bF_buf2), .Y(_9448_) );
OAI21X1 OAI21X1_2648 ( .gnd(gnd), .vdd(vdd), .A(_9363_), .B(_9295_), .C(_9294__bF_buf3), .Y(_9449_) );
AOI21X1 AOI21X1_1679 ( .gnd(gnd), .vdd(vdd), .A(_9448_), .B(_9447_), .C(_9449_), .Y(_9450_) );
NOR2X1 NOR2X1_1553 ( .gnd(gnd), .vdd(vdd), .A(_8862__bF_buf0), .B(_9294__bF_buf2), .Y(_9451_) );
OAI21X1 OAI21X1_2649 ( .gnd(gnd), .vdd(vdd), .A(_9450_), .B(_9451_), .C(_9290__bF_buf2), .Y(_9452_) );
NAND2X1 NAND2X1_1196 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe59), .B(_9363_), .Y(_9453_) );
NAND3X1 NAND3X1_438 ( .gnd(gnd), .vdd(vdd), .A(_9292__bF_buf2), .B(_9453_), .C(_9452_), .Y(_9454_) );
NAND3X1 NAND3X1_439 ( .gnd(gnd), .vdd(vdd), .A(_9291_), .B(_9348_), .C(_9454_), .Y(_9455_) );
NAND2X1 NAND2X1_1197 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe61_bF_buf2), .B(_9363_), .Y(_9456_) );
NAND3X1 NAND3X1_440 ( .gnd(gnd), .vdd(vdd), .A(_9287__bF_buf3), .B(_9456_), .C(_9455_), .Y(_9457_) );
NAND3X1 NAND3X1_441 ( .gnd(gnd), .vdd(vdd), .A(_9289__bF_buf2), .B(_9347_), .C(_9457_), .Y(_9458_) );
NAND2X1 NAND2X1_1198 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe63), .B(_9363_), .Y(_9459_) );
NAND3X1 NAND3X1_442 ( .gnd(gnd), .vdd(vdd), .A(_9288__bF_buf2), .B(_9459_), .C(_9458_), .Y(_9460_) );
NAND3X1 NAND3X1_443 ( .gnd(gnd), .vdd(vdd), .A(_9284_), .B(_9346_), .C(_9460_), .Y(_9461_) );
AOI21X1 AOI21X1_1680 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe65_bF_buf2), .B(_9363_), .C(micro_hash_ucr_3_pipe66_bF_buf3), .Y(_9462_) );
OAI21X1 OAI21X1_2650 ( .gnd(gnd), .vdd(vdd), .A(_9286__bF_buf2), .B(micro_hash_ucr_3_a_0_bF_buf0_), .C(_9285__bF_buf2), .Y(_9463_) );
AOI21X1 AOI21X1_1681 ( .gnd(gnd), .vdd(vdd), .A(_9462_), .B(_9461_), .C(_9463_), .Y(_9464_) );
OAI21X1 OAI21X1_2651 ( .gnd(gnd), .vdd(vdd), .A(_9397_), .B(_9285__bF_buf1), .C(_9282__bF_buf3), .Y(_9465_) );
NAND2X1 NAND2X1_1199 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe68_bF_buf2), .B(_8862__bF_buf3), .Y(_9466_) );
OAI21X1 OAI21X1_2652 ( .gnd(gnd), .vdd(vdd), .A(_9464_), .B(_9465_), .C(_9466_), .Y(_9467_) );
OAI21X1 OAI21X1_2653 ( .gnd(gnd), .vdd(vdd), .A(_9363_), .B(_9283__bF_buf2), .C(_8705__bF_buf2), .Y(_9468_) );
AOI21X1 AOI21X1_1682 ( .gnd(gnd), .vdd(vdd), .A(_9283__bF_buf1), .B(_9467_), .C(_9468_), .Y(_8700__0_) );
NAND2X1 NAND2X1_1200 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_1_bF_buf1_), .B(micro_hash_ucr_3_pipe66_bF_buf2), .Y(_9469_) );
NAND2X1 NAND2X1_1201 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_1_bF_buf0_), .B(micro_hash_ucr_3_pipe64_bF_buf2), .Y(_9470_) );
NAND2X1 NAND2X1_1202 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_1_bF_buf3_), .B(micro_hash_ucr_3_pipe62_bF_buf1), .Y(_9471_) );
NAND2X1 NAND2X1_1203 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_1_bF_buf2_), .B(micro_hash_ucr_3_pipe52_bF_buf2), .Y(_9472_) );
NAND2X1 NAND2X1_1204 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe46_bF_buf3), .B(_8868__bF_buf2), .Y(_9473_) );
NAND2X1 NAND2X1_1205 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_1_bF_buf1_), .B(micro_hash_ucr_3_pipe40_bF_buf1), .Y(_9474_) );
NAND2X1 NAND2X1_1206 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_1_bF_buf0_), .B(micro_hash_ucr_3_pipe38_bF_buf0), .Y(_9475_) );
NAND2X1 NAND2X1_1207 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_1_bF_buf3_), .B(micro_hash_ucr_3_pipe36_bF_buf1), .Y(_9476_) );
NAND2X1 NAND2X1_1208 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_1_bF_buf2_), .B(micro_hash_ucr_3_pipe34_bF_buf2), .Y(_9477_) );
NAND2X1 NAND2X1_1209 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_1_bF_buf1_), .B(micro_hash_ucr_3_pipe32_bF_buf1), .Y(_9478_) );
NAND2X1 NAND2X1_1210 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe26_bF_buf1), .B(_8868__bF_buf1), .Y(_9479_) );
NAND2X1 NAND2X1_1211 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe24_bF_buf2), .B(_8868__bF_buf0), .Y(_9480_) );
NAND2X1 NAND2X1_1212 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_1_bF_buf0_), .B(micro_hash_ucr_3_pipe18_bF_buf2), .Y(_9481_) );
NOR2X1 NOR2X1_1554 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_1_bF_buf1_), .B(micro_hash_ucr_3_b_1_bF_buf1_), .Y(_9482_) );
INVX8 INVX8_266 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_1_bF_buf0_), .Y(_9483_) );
NOR2X1 NOR2X1_1555 ( .gnd(gnd), .vdd(vdd), .A(_9483_), .B(_12908__bF_buf2), .Y(_9484_) );
NOR2X1 NOR2X1_1556 ( .gnd(gnd), .vdd(vdd), .A(_9482_), .B(_9484_), .Y(_9485_) );
OAI21X1 OAI21X1_2654 ( .gnd(gnd), .vdd(vdd), .A(_9344_), .B(micro_hash_ucr_3_pipe8), .C(_9343_), .Y(_9486_) );
AOI21X1 AOI21X1_1683 ( .gnd(gnd), .vdd(vdd), .A(_9342_), .B(_9486_), .C(micro_hash_ucr_3_pipe11), .Y(_9487_) );
OAI21X1 OAI21X1_2655 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe7), .B(micro_hash_ucr_3_pipe6_bF_buf1), .C(_9341_), .Y(_9488_) );
NOR2X1 NOR2X1_1557 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe7), .B(micro_hash_ucr_3_pipe6_bF_buf0), .Y(_9489_) );
OAI21X1 OAI21X1_2656 ( .gnd(gnd), .vdd(vdd), .A(_9489_), .B(micro_hash_ucr_3_pipe8), .C(_8868__bF_buf3), .Y(_9490_) );
NAND3X1 NAND3X1_444 ( .gnd(gnd), .vdd(vdd), .A(_8866_), .B(_9342_), .C(_9344_), .Y(_9491_) );
OAI21X1 OAI21X1_2657 ( .gnd(gnd), .vdd(vdd), .A(_9488_), .B(_9491_), .C(_9490_), .Y(_9492_) );
AOI22X1 AOI22X1_66 ( .gnd(gnd), .vdd(vdd), .A(_8868__bF_buf2), .B(micro_hash_ucr_3_pipe10_bF_buf3), .C(_9492_), .D(_9343_), .Y(_9493_) );
OAI22X1 OAI22X1_112 ( .gnd(gnd), .vdd(vdd), .A(_9485_), .B(_9487_), .C(_9493_), .D(micro_hash_ucr_3_pipe11), .Y(_9494_) );
NOR2X1 NOR2X1_1558 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe13), .B(micro_hash_ucr_3_pipe12), .Y(_9495_) );
OAI22X1 OAI22X1_113 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_1_bF_buf3_), .B(_9379_), .C(_9485_), .D(_9339_), .Y(_9496_) );
AOI21X1 AOI21X1_1684 ( .gnd(gnd), .vdd(vdd), .A(_9495_), .B(_9494_), .C(_9496_), .Y(_9497_) );
AOI21X1 AOI21X1_1685 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe14_bF_buf1), .B(_8868__bF_buf1), .C(micro_hash_ucr_3_pipe15_bF_buf0), .Y(_9498_) );
OAI21X1 OAI21X1_2658 ( .gnd(gnd), .vdd(vdd), .A(_9497_), .B(micro_hash_ucr_3_pipe14_bF_buf0), .C(_9498_), .Y(_9499_) );
AOI21X1 AOI21X1_1686 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe15_bF_buf3), .B(_9485_), .C(micro_hash_ucr_3_pipe16_bF_buf2), .Y(_9500_) );
AOI22X1 AOI22X1_67 ( .gnd(gnd), .vdd(vdd), .A(_8868__bF_buf0), .B(micro_hash_ucr_3_pipe16_bF_buf1), .C(_9499_), .D(_9500_), .Y(_9501_) );
OAI21X1 OAI21X1_2659 ( .gnd(gnd), .vdd(vdd), .A(_9484_), .B(_9482_), .C(micro_hash_ucr_3_pipe17_bF_buf1), .Y(_9502_) );
OAI21X1 OAI21X1_2660 ( .gnd(gnd), .vdd(vdd), .A(_9501_), .B(micro_hash_ucr_3_pipe17_bF_buf0), .C(_9502_), .Y(_9503_) );
OAI21X1 OAI21X1_2661 ( .gnd(gnd), .vdd(vdd), .A(_9503_), .B(micro_hash_ucr_3_pipe18_bF_buf1), .C(_9481_), .Y(_9504_) );
INVX4 INVX4_148 ( .gnd(gnd), .vdd(vdd), .A(_9485_), .Y(_9505_) );
OAI21X1 OAI21X1_2662 ( .gnd(gnd), .vdd(vdd), .A(_9505_), .B(_9333__bF_buf1), .C(_9329__bF_buf2), .Y(_9506_) );
AOI21X1 AOI21X1_1687 ( .gnd(gnd), .vdd(vdd), .A(_9333__bF_buf0), .B(_9504_), .C(_9506_), .Y(_9507_) );
OAI21X1 OAI21X1_2663 ( .gnd(gnd), .vdd(vdd), .A(_9329__bF_buf1), .B(micro_hash_ucr_3_a_1_bF_buf2_), .C(_9331_), .Y(_9508_) );
AOI21X1 AOI21X1_1688 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe21_bF_buf1), .B(_9485_), .C(micro_hash_ucr_3_pipe22_bF_buf2), .Y(_9509_) );
OAI21X1 OAI21X1_2664 ( .gnd(gnd), .vdd(vdd), .A(_9507_), .B(_9508_), .C(_9509_), .Y(_9510_) );
NAND2X1 NAND2X1_1213 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe22_bF_buf1), .B(_8868__bF_buf3), .Y(_9511_) );
NAND3X1 NAND3X1_445 ( .gnd(gnd), .vdd(vdd), .A(_9326__bF_buf1), .B(_9511_), .C(_9510_), .Y(_9512_) );
NAND2X1 NAND2X1_1214 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe23), .B(_9485_), .Y(_9513_) );
NAND3X1 NAND3X1_446 ( .gnd(gnd), .vdd(vdd), .A(_9328__bF_buf1), .B(_9513_), .C(_9512_), .Y(_9514_) );
NAND3X1 NAND3X1_447 ( .gnd(gnd), .vdd(vdd), .A(_9327_), .B(_9480_), .C(_9514_), .Y(_9515_) );
NAND2X1 NAND2X1_1215 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe25_bF_buf1), .B(_9485_), .Y(_9516_) );
NAND3X1 NAND3X1_448 ( .gnd(gnd), .vdd(vdd), .A(_9323__bF_buf2), .B(_9516_), .C(_9515_), .Y(_9517_) );
NAND3X1 NAND3X1_449 ( .gnd(gnd), .vdd(vdd), .A(_9325__bF_buf1), .B(_9479_), .C(_9517_), .Y(_9518_) );
NAND2X1 NAND2X1_1216 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe27), .B(_9485_), .Y(_9519_) );
AOI21X1 AOI21X1_1689 ( .gnd(gnd), .vdd(vdd), .A(_9519_), .B(_9518_), .C(micro_hash_ucr_3_pipe28_bF_buf2), .Y(_9520_) );
OAI21X1 OAI21X1_2665 ( .gnd(gnd), .vdd(vdd), .A(_8868__bF_buf2), .B(_9324__bF_buf2), .C(_9320_), .Y(_9521_) );
AOI21X1 AOI21X1_1690 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe29_bF_buf1), .B(_9505_), .C(micro_hash_ucr_3_pipe30_bF_buf2), .Y(_9522_) );
OAI21X1 OAI21X1_2666 ( .gnd(gnd), .vdd(vdd), .A(_9520_), .B(_9521_), .C(_9522_), .Y(_9523_) );
NAND2X1 NAND2X1_1217 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_1_bF_buf1_), .B(micro_hash_ucr_3_pipe30_bF_buf1), .Y(_9524_) );
NAND3X1 NAND3X1_450 ( .gnd(gnd), .vdd(vdd), .A(_9321__bF_buf1), .B(_9524_), .C(_9523_), .Y(_9525_) );
OAI21X1 OAI21X1_2667 ( .gnd(gnd), .vdd(vdd), .A(_9484_), .B(_9482_), .C(micro_hash_ucr_3_pipe31), .Y(_9526_) );
NAND3X1 NAND3X1_451 ( .gnd(gnd), .vdd(vdd), .A(_9317__bF_buf2), .B(_9526_), .C(_9525_), .Y(_9527_) );
NAND3X1 NAND3X1_452 ( .gnd(gnd), .vdd(vdd), .A(_9319_), .B(_9478_), .C(_9527_), .Y(_9528_) );
OAI21X1 OAI21X1_2668 ( .gnd(gnd), .vdd(vdd), .A(_9484_), .B(_9482_), .C(micro_hash_ucr_3_pipe33_bF_buf0), .Y(_9529_) );
NAND3X1 NAND3X1_453 ( .gnd(gnd), .vdd(vdd), .A(_9318__bF_buf2), .B(_9529_), .C(_9528_), .Y(_9530_) );
NAND3X1 NAND3X1_454 ( .gnd(gnd), .vdd(vdd), .A(_9314_), .B(_9477_), .C(_9530_), .Y(_9531_) );
OAI21X1 OAI21X1_2669 ( .gnd(gnd), .vdd(vdd), .A(_9484_), .B(_9482_), .C(micro_hash_ucr_3_pipe35_bF_buf0), .Y(_9532_) );
NAND3X1 NAND3X1_455 ( .gnd(gnd), .vdd(vdd), .A(_9316__bF_buf2), .B(_9532_), .C(_9531_), .Y(_9533_) );
NAND3X1 NAND3X1_456 ( .gnd(gnd), .vdd(vdd), .A(_9315_), .B(_9476_), .C(_9533_), .Y(_9534_) );
OAI21X1 OAI21X1_2670 ( .gnd(gnd), .vdd(vdd), .A(_9484_), .B(_9482_), .C(micro_hash_ucr_3_pipe37_bF_buf0), .Y(_9535_) );
NAND3X1 NAND3X1_457 ( .gnd(gnd), .vdd(vdd), .A(_9311__bF_buf3), .B(_9535_), .C(_9534_), .Y(_9536_) );
NAND3X1 NAND3X1_458 ( .gnd(gnd), .vdd(vdd), .A(_9313_), .B(_9475_), .C(_9536_), .Y(_9537_) );
OAI21X1 OAI21X1_2671 ( .gnd(gnd), .vdd(vdd), .A(_9484_), .B(_9482_), .C(micro_hash_ucr_3_pipe39_bF_buf0), .Y(_9538_) );
NAND3X1 NAND3X1_459 ( .gnd(gnd), .vdd(vdd), .A(_9312__bF_buf2), .B(_9538_), .C(_9537_), .Y(_9539_) );
AOI21X1 AOI21X1_1691 ( .gnd(gnd), .vdd(vdd), .A(_9474_), .B(_9539_), .C(micro_hash_ucr_3_pipe41_bF_buf0), .Y(_9540_) );
OAI21X1 OAI21X1_2672 ( .gnd(gnd), .vdd(vdd), .A(_9505_), .B(_9308_), .C(_9310__bF_buf2), .Y(_9541_) );
AOI21X1 AOI21X1_1692 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe42_bF_buf1), .B(_8868__bF_buf1), .C(micro_hash_ucr_3_pipe43), .Y(_9542_) );
OAI21X1 OAI21X1_2673 ( .gnd(gnd), .vdd(vdd), .A(_9540_), .B(_9541_), .C(_9542_), .Y(_9543_) );
AOI21X1 AOI21X1_1693 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe43), .B(_9485_), .C(micro_hash_ucr_3_pipe44_bF_buf0), .Y(_9544_) );
NAND2X1 NAND2X1_1218 ( .gnd(gnd), .vdd(vdd), .A(_9544_), .B(_9543_), .Y(_9545_) );
NAND2X1 NAND2X1_1219 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe44_bF_buf3), .B(_8868__bF_buf0), .Y(_9546_) );
NAND3X1 NAND3X1_460 ( .gnd(gnd), .vdd(vdd), .A(_9307_), .B(_9546_), .C(_9545_), .Y(_9547_) );
NAND2X1 NAND2X1_1220 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe45_bF_buf1), .B(_9485_), .Y(_9548_) );
NAND3X1 NAND3X1_461 ( .gnd(gnd), .vdd(vdd), .A(_9306__bF_buf0), .B(_9548_), .C(_9547_), .Y(_9549_) );
NAND3X1 NAND3X1_462 ( .gnd(gnd), .vdd(vdd), .A(_9302_), .B(_9473_), .C(_9549_), .Y(_9550_) );
NAND2X1 NAND2X1_1221 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe47), .B(_9485_), .Y(_9551_) );
AOI21X1 AOI21X1_1694 ( .gnd(gnd), .vdd(vdd), .A(_9551_), .B(_9550_), .C(micro_hash_ucr_3_pipe48_bF_buf2), .Y(_9552_) );
OAI21X1 OAI21X1_2674 ( .gnd(gnd), .vdd(vdd), .A(_8868__bF_buf3), .B(_9304__bF_buf1), .C(_9303_), .Y(_9553_) );
AOI21X1 AOI21X1_1695 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe49_bF_buf1), .B(_9505_), .C(micro_hash_ucr_3_pipe50_bF_buf2), .Y(_9554_) );
OAI21X1 OAI21X1_2675 ( .gnd(gnd), .vdd(vdd), .A(_9552_), .B(_9553_), .C(_9554_), .Y(_9555_) );
NAND2X1 NAND2X1_1222 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_1_bF_buf0_), .B(micro_hash_ucr_3_pipe50_bF_buf1), .Y(_9556_) );
NAND3X1 NAND3X1_463 ( .gnd(gnd), .vdd(vdd), .A(_9301__bF_buf1), .B(_9556_), .C(_9555_), .Y(_9557_) );
OAI21X1 OAI21X1_2676 ( .gnd(gnd), .vdd(vdd), .A(_9484_), .B(_9482_), .C(micro_hash_ucr_3_pipe51), .Y(_9558_) );
NAND3X1 NAND3X1_464 ( .gnd(gnd), .vdd(vdd), .A(_9300__bF_buf1), .B(_9558_), .C(_9557_), .Y(_9559_) );
AOI21X1 AOI21X1_1696 ( .gnd(gnd), .vdd(vdd), .A(_9472_), .B(_9559_), .C(micro_hash_ucr_3_pipe53), .Y(_9560_) );
OAI21X1 OAI21X1_2677 ( .gnd(gnd), .vdd(vdd), .A(_9505_), .B(_9296_), .C(_9298__bF_buf2), .Y(_9561_) );
AOI21X1 AOI21X1_1697 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe54_bF_buf1), .B(_8868__bF_buf2), .C(micro_hash_ucr_3_pipe55), .Y(_9562_) );
OAI21X1 OAI21X1_2678 ( .gnd(gnd), .vdd(vdd), .A(_9560_), .B(_9561_), .C(_9562_), .Y(_9563_) );
AOI21X1 AOI21X1_1698 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe55), .B(_9485_), .C(micro_hash_ucr_3_pipe56_bF_buf2), .Y(_9564_) );
NAND2X1 NAND2X1_1223 ( .gnd(gnd), .vdd(vdd), .A(_9564_), .B(_9563_), .Y(_9565_) );
NAND2X1 NAND2X1_1224 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe56_bF_buf1), .B(_8868__bF_buf1), .Y(_9566_) );
NAND3X1 NAND3X1_465 ( .gnd(gnd), .vdd(vdd), .A(_9295_), .B(_9566_), .C(_9565_), .Y(_9567_) );
NAND2X1 NAND2X1_1225 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe57_bF_buf1), .B(_9485_), .Y(_9568_) );
AOI21X1 AOI21X1_1699 ( .gnd(gnd), .vdd(vdd), .A(_9568_), .B(_9567_), .C(micro_hash_ucr_3_pipe58_bF_buf2), .Y(_9569_) );
OAI21X1 OAI21X1_2679 ( .gnd(gnd), .vdd(vdd), .A(_8868__bF_buf0), .B(_9294__bF_buf1), .C(_9290__bF_buf1), .Y(_9570_) );
AOI21X1 AOI21X1_1700 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe59), .B(_9505_), .C(micro_hash_ucr_3_pipe60_bF_buf2), .Y(_9571_) );
OAI21X1 OAI21X1_2680 ( .gnd(gnd), .vdd(vdd), .A(_9569_), .B(_9570_), .C(_9571_), .Y(_9572_) );
NAND2X1 NAND2X1_1226 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_1_bF_buf3_), .B(micro_hash_ucr_3_pipe60_bF_buf1), .Y(_9573_) );
NAND3X1 NAND3X1_466 ( .gnd(gnd), .vdd(vdd), .A(_9291_), .B(_9573_), .C(_9572_), .Y(_9574_) );
OAI21X1 OAI21X1_2681 ( .gnd(gnd), .vdd(vdd), .A(_9484_), .B(_9482_), .C(micro_hash_ucr_3_pipe61_bF_buf1), .Y(_9575_) );
NAND3X1 NAND3X1_467 ( .gnd(gnd), .vdd(vdd), .A(_9287__bF_buf2), .B(_9575_), .C(_9574_), .Y(_9576_) );
NAND3X1 NAND3X1_468 ( .gnd(gnd), .vdd(vdd), .A(_9289__bF_buf1), .B(_9471_), .C(_9576_), .Y(_9577_) );
OAI21X1 OAI21X1_2682 ( .gnd(gnd), .vdd(vdd), .A(_9484_), .B(_9482_), .C(micro_hash_ucr_3_pipe63), .Y(_9578_) );
NAND3X1 NAND3X1_469 ( .gnd(gnd), .vdd(vdd), .A(_9288__bF_buf1), .B(_9578_), .C(_9577_), .Y(_9579_) );
NAND3X1 NAND3X1_470 ( .gnd(gnd), .vdd(vdd), .A(_9284_), .B(_9470_), .C(_9579_), .Y(_9580_) );
OAI21X1 OAI21X1_2683 ( .gnd(gnd), .vdd(vdd), .A(_9484_), .B(_9482_), .C(micro_hash_ucr_3_pipe65_bF_buf1), .Y(_9581_) );
NAND3X1 NAND3X1_471 ( .gnd(gnd), .vdd(vdd), .A(_9286__bF_buf1), .B(_9581_), .C(_9580_), .Y(_9582_) );
NAND3X1 NAND3X1_472 ( .gnd(gnd), .vdd(vdd), .A(_9285__bF_buf0), .B(_9469_), .C(_9582_), .Y(_9583_) );
OAI21X1 OAI21X1_2684 ( .gnd(gnd), .vdd(vdd), .A(_9484_), .B(_9482_), .C(micro_hash_ucr_3_pipe67), .Y(_9584_) );
NAND3X1 NAND3X1_473 ( .gnd(gnd), .vdd(vdd), .A(_9282__bF_buf2), .B(_9584_), .C(_9583_), .Y(_9585_) );
AOI21X1 AOI21X1_1701 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_1_bF_buf2_), .B(micro_hash_ucr_3_pipe68_bF_buf1), .C(micro_hash_ucr_3_pipe69), .Y(_9586_) );
OAI21X1 OAI21X1_2685 ( .gnd(gnd), .vdd(vdd), .A(_9485_), .B(_9283__bF_buf0), .C(_8705__bF_buf1), .Y(_9587_) );
AOI21X1 AOI21X1_1702 ( .gnd(gnd), .vdd(vdd), .A(_9586_), .B(_9585_), .C(_9587_), .Y(_8700__1_) );
NOR2X1 NOR2X1_1559 ( .gnd(gnd), .vdd(vdd), .A(_8884_), .B(_9287__bF_buf1), .Y(_9588_) );
NOR2X1 NOR2X1_1560 ( .gnd(gnd), .vdd(vdd), .A(_8884_), .B(_9292__bF_buf1), .Y(_9589_) );
NOR2X1 NOR2X1_1561 ( .gnd(gnd), .vdd(vdd), .A(_8884_), .B(_9294__bF_buf0), .Y(_9590_) );
NOR2X1 NOR2X1_1562 ( .gnd(gnd), .vdd(vdd), .A(_8884_), .B(_9293__bF_buf1), .Y(_9591_) );
NOR2X1 NOR2X1_1563 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_2_), .B(micro_hash_ucr_3_b_2_bF_buf1_), .Y(_9592_) );
INVX8 INVX8_267 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_2_), .Y(_9593_) );
NOR2X1 NOR2X1_1564 ( .gnd(gnd), .vdd(vdd), .A(_9593__bF_buf3), .B(_8789__bF_buf2), .Y(_9594_) );
NOR2X1 NOR2X1_1565 ( .gnd(gnd), .vdd(vdd), .A(_9592_), .B(_9594_), .Y(_9595_) );
INVX8 INVX8_268 ( .gnd(gnd), .vdd(vdd), .A(_9595_), .Y(_9596_) );
NOR2X1 NOR2X1_1566 ( .gnd(gnd), .vdd(vdd), .A(_8884_), .B(_9306__bF_buf3), .Y(_9597_) );
NAND2X1 NAND2X1_1227 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_2_), .B(micro_hash_ucr_3_pipe34_bF_buf1), .Y(_9598_) );
OAI21X1 OAI21X1_2686 ( .gnd(gnd), .vdd(vdd), .A(_9487_), .B(micro_hash_ucr_3_pipe12), .C(_9339_), .Y(_9599_) );
AOI21X1 AOI21X1_1703 ( .gnd(gnd), .vdd(vdd), .A(_9335__bF_buf1), .B(_9599_), .C(micro_hash_ucr_3_pipe15_bF_buf2), .Y(_9600_) );
OAI21X1 OAI21X1_2687 ( .gnd(gnd), .vdd(vdd), .A(_9600_), .B(micro_hash_ucr_3_pipe16_bF_buf0), .C(_9332_), .Y(_9601_) );
INVX1 INVX1_625 ( .gnd(gnd), .vdd(vdd), .A(_9601_), .Y(_9602_) );
OAI21X1 OAI21X1_2688 ( .gnd(gnd), .vdd(vdd), .A(_9602_), .B(micro_hash_ucr_3_pipe18_bF_buf0), .C(_9333__bF_buf3), .Y(_9603_) );
AOI21X1 AOI21X1_1704 ( .gnd(gnd), .vdd(vdd), .A(_9329__bF_buf0), .B(_9603_), .C(micro_hash_ucr_3_pipe21_bF_buf0), .Y(_9604_) );
OAI21X1 OAI21X1_2689 ( .gnd(gnd), .vdd(vdd), .A(_9604_), .B(micro_hash_ucr_3_pipe22_bF_buf0), .C(_9326__bF_buf0), .Y(_9605_) );
AOI21X1 AOI21X1_1705 ( .gnd(gnd), .vdd(vdd), .A(_9328__bF_buf0), .B(_9605_), .C(micro_hash_ucr_3_pipe25_bF_buf0), .Y(_9606_) );
OAI21X1 OAI21X1_2690 ( .gnd(gnd), .vdd(vdd), .A(_9606_), .B(micro_hash_ucr_3_pipe26_bF_buf0), .C(_9325__bF_buf0), .Y(_9607_) );
OAI21X1 OAI21X1_2691 ( .gnd(gnd), .vdd(vdd), .A(_9592_), .B(_9594_), .C(_9607_), .Y(_9608_) );
NOR2X1 NOR2X1_1567 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe11), .B(micro_hash_ucr_3_pipe10_bF_buf2), .Y(_9609_) );
NAND2X1 NAND2X1_1228 ( .gnd(gnd), .vdd(vdd), .A(_9495_), .B(_9609_), .Y(_9610_) );
NOR2X1 NOR2X1_1568 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe19), .B(micro_hash_ucr_3_pipe18_bF_buf4), .Y(_9611_) );
NAND3X1 NAND3X1_474 ( .gnd(gnd), .vdd(vdd), .A(_9335__bF_buf0), .B(_9344_), .C(_9611_), .Y(_9612_) );
NOR2X1 NOR2X1_1569 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe20_bF_buf2), .B(micro_hash_ucr_3_pipe22_bF_buf4), .Y(_9613_) );
NAND3X1 NAND3X1_475 ( .gnd(gnd), .vdd(vdd), .A(_9331_), .B(_9332_), .C(_9613_), .Y(_9614_) );
OR2X2 OR2X2_68 ( .gnd(gnd), .vdd(vdd), .A(_9612_), .B(_9614_), .Y(_9615_) );
NOR2X1 NOR2X1_1570 ( .gnd(gnd), .vdd(vdd), .A(_9610_), .B(_9615_), .Y(_9616_) );
NOR2X1 NOR2X1_1571 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe9), .B(_9488_), .Y(_9617_) );
NOR2X1 NOR2X1_1572 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe27), .B(micro_hash_ucr_3_pipe23), .Y(_9618_) );
NAND3X1 NAND3X1_476 ( .gnd(gnd), .vdd(vdd), .A(_9327_), .B(_9328__bF_buf3), .C(_9618_), .Y(_9619_) );
NOR2X1 NOR2X1_1573 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe16_bF_buf4), .B(micro_hash_ucr_3_pipe15_bF_buf1), .Y(_9620_) );
NAND3X1 NAND3X1_477 ( .gnd(gnd), .vdd(vdd), .A(_8874_), .B(_9323__bF_buf1), .C(_9620_), .Y(_9621_) );
NOR2X1 NOR2X1_1574 ( .gnd(gnd), .vdd(vdd), .A(_9619_), .B(_9621_), .Y(_9622_) );
NAND3X1 NAND3X1_478 ( .gnd(gnd), .vdd(vdd), .A(_9617_), .B(_9622_), .C(_9616_), .Y(_9623_) );
AOI21X1 AOI21X1_1706 ( .gnd(gnd), .vdd(vdd), .A(_9623_), .B(_9608_), .C(micro_hash_ucr_3_pipe28_bF_buf1), .Y(_9624_) );
AOI21X1 AOI21X1_1707 ( .gnd(gnd), .vdd(vdd), .A(_9338_), .B(_9371_), .C(micro_hash_ucr_3_pipe12), .Y(_9625_) );
OAI21X1 OAI21X1_2692 ( .gnd(gnd), .vdd(vdd), .A(_9625_), .B(micro_hash_ucr_3_pipe13), .C(_9335__bF_buf3), .Y(_9626_) );
AOI21X1 AOI21X1_1708 ( .gnd(gnd), .vdd(vdd), .A(_9337_), .B(_9626_), .C(micro_hash_ucr_3_pipe16_bF_buf3), .Y(_9627_) );
OAI21X1 OAI21X1_2693 ( .gnd(gnd), .vdd(vdd), .A(_9627_), .B(micro_hash_ucr_3_pipe17_bF_buf3), .C(_9334__bF_buf1), .Y(_9628_) );
AOI21X1 AOI21X1_1709 ( .gnd(gnd), .vdd(vdd), .A(_9333__bF_buf2), .B(_9628_), .C(micro_hash_ucr_3_pipe20_bF_buf1), .Y(_9629_) );
OAI21X1 OAI21X1_2694 ( .gnd(gnd), .vdd(vdd), .A(_9629_), .B(micro_hash_ucr_3_pipe21_bF_buf3), .C(_9330__bF_buf2), .Y(_9630_) );
AOI21X1 AOI21X1_1710 ( .gnd(gnd), .vdd(vdd), .A(_9326__bF_buf3), .B(_9630_), .C(micro_hash_ucr_3_pipe24_bF_buf1), .Y(_9631_) );
OAI21X1 OAI21X1_2695 ( .gnd(gnd), .vdd(vdd), .A(_9631_), .B(micro_hash_ucr_3_pipe25_bF_buf3), .C(_9323__bF_buf0), .Y(_9632_) );
AOI21X1 AOI21X1_1711 ( .gnd(gnd), .vdd(vdd), .A(_9325__bF_buf3), .B(_9632_), .C(micro_hash_ucr_3_pipe28_bF_buf0), .Y(_9633_) );
OAI21X1 OAI21X1_2696 ( .gnd(gnd), .vdd(vdd), .A(_9633_), .B(micro_hash_ucr_3_a_2_), .C(_9320_), .Y(_9634_) );
AOI21X1 AOI21X1_1712 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe29_bF_buf0), .B(_9595_), .C(micro_hash_ucr_3_pipe30_bF_buf0), .Y(_9635_) );
OAI21X1 OAI21X1_2697 ( .gnd(gnd), .vdd(vdd), .A(_9624_), .B(_9634_), .C(_9635_), .Y(_9636_) );
AOI21X1 AOI21X1_1713 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe30_bF_buf4), .B(_8884_), .C(micro_hash_ucr_3_pipe31), .Y(_9637_) );
OAI21X1 OAI21X1_2698 ( .gnd(gnd), .vdd(vdd), .A(_9596_), .B(_9321__bF_buf0), .C(_9317__bF_buf1), .Y(_9638_) );
AOI21X1 AOI21X1_1714 ( .gnd(gnd), .vdd(vdd), .A(_9637_), .B(_9636_), .C(_9638_), .Y(_9639_) );
NOR2X1 NOR2X1_1575 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_2_), .B(_9317__bF_buf0), .Y(_9640_) );
OAI21X1 OAI21X1_2699 ( .gnd(gnd), .vdd(vdd), .A(_9639_), .B(_9640_), .C(_9319_), .Y(_9641_) );
OAI21X1 OAI21X1_2700 ( .gnd(gnd), .vdd(vdd), .A(_9319_), .B(_9595_), .C(_9641_), .Y(_9642_) );
OAI21X1 OAI21X1_2701 ( .gnd(gnd), .vdd(vdd), .A(_9642_), .B(micro_hash_ucr_3_pipe34_bF_buf0), .C(_9598_), .Y(_9643_) );
NAND2X1 NAND2X1_1229 ( .gnd(gnd), .vdd(vdd), .A(_9314_), .B(_9643_), .Y(_9644_) );
OAI21X1 OAI21X1_2702 ( .gnd(gnd), .vdd(vdd), .A(_9314_), .B(_9596_), .C(_9644_), .Y(_9645_) );
AOI21X1 AOI21X1_1715 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe36_bF_buf0), .B(_8884_), .C(micro_hash_ucr_3_pipe37_bF_buf3), .Y(_9646_) );
OAI21X1 OAI21X1_2703 ( .gnd(gnd), .vdd(vdd), .A(_9645_), .B(micro_hash_ucr_3_pipe36_bF_buf4), .C(_9646_), .Y(_9647_) );
OAI21X1 OAI21X1_2704 ( .gnd(gnd), .vdd(vdd), .A(_9315_), .B(_9596_), .C(_9647_), .Y(_9648_) );
NAND2X1 NAND2X1_1230 ( .gnd(gnd), .vdd(vdd), .A(_9311__bF_buf2), .B(_9648_), .Y(_9649_) );
OAI21X1 OAI21X1_2705 ( .gnd(gnd), .vdd(vdd), .A(_8884_), .B(_9311__bF_buf1), .C(_9649_), .Y(_9650_) );
AOI21X1 AOI21X1_1716 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe39_bF_buf3), .B(_9596_), .C(micro_hash_ucr_3_pipe40_bF_buf0), .Y(_9651_) );
OAI21X1 OAI21X1_2706 ( .gnd(gnd), .vdd(vdd), .A(_9650_), .B(micro_hash_ucr_3_pipe39_bF_buf2), .C(_9651_), .Y(_9652_) );
OAI21X1 OAI21X1_2707 ( .gnd(gnd), .vdd(vdd), .A(_8884_), .B(_9312__bF_buf1), .C(_9652_), .Y(_9653_) );
AND2X2 AND2X2_680 ( .gnd(gnd), .vdd(vdd), .A(_9653_), .B(_9308_), .Y(_9654_) );
NOR2X1 NOR2X1_1576 ( .gnd(gnd), .vdd(vdd), .A(_9308_), .B(_9596_), .Y(_9655_) );
OAI21X1 OAI21X1_2708 ( .gnd(gnd), .vdd(vdd), .A(_9654_), .B(_9655_), .C(_9310__bF_buf1), .Y(_9656_) );
AOI21X1 AOI21X1_1717 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_2_), .B(micro_hash_ucr_3_pipe42_bF_buf0), .C(micro_hash_ucr_3_pipe43), .Y(_9657_) );
OAI21X1 OAI21X1_2709 ( .gnd(gnd), .vdd(vdd), .A(_9595_), .B(_9309__bF_buf2), .C(_9305__bF_buf3), .Y(_9658_) );
AOI21X1 AOI21X1_1718 ( .gnd(gnd), .vdd(vdd), .A(_9657_), .B(_9656_), .C(_9658_), .Y(_9659_) );
NOR2X1 NOR2X1_1577 ( .gnd(gnd), .vdd(vdd), .A(_8884_), .B(_9305__bF_buf2), .Y(_9660_) );
OAI21X1 OAI21X1_2710 ( .gnd(gnd), .vdd(vdd), .A(_9659_), .B(_9660_), .C(_9307_), .Y(_9661_) );
OAI21X1 OAI21X1_2711 ( .gnd(gnd), .vdd(vdd), .A(_9307_), .B(_9596_), .C(_9661_), .Y(_9662_) );
AND2X2 AND2X2_681 ( .gnd(gnd), .vdd(vdd), .A(_9662_), .B(_9306__bF_buf2), .Y(_9663_) );
OAI21X1 OAI21X1_2712 ( .gnd(gnd), .vdd(vdd), .A(_9663_), .B(_9597_), .C(_9302_), .Y(_9664_) );
OAI21X1 OAI21X1_2713 ( .gnd(gnd), .vdd(vdd), .A(_9302_), .B(_9596_), .C(_9664_), .Y(_9665_) );
AND2X2 AND2X2_682 ( .gnd(gnd), .vdd(vdd), .A(_9665_), .B(_9304__bF_buf0), .Y(_9666_) );
OAI21X1 OAI21X1_2714 ( .gnd(gnd), .vdd(vdd), .A(_8884_), .B(_9304__bF_buf3), .C(_9303_), .Y(_9667_) );
AOI21X1 AOI21X1_1719 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe49_bF_buf0), .B(_9596_), .C(micro_hash_ucr_3_pipe50_bF_buf0), .Y(_9668_) );
OAI21X1 OAI21X1_2715 ( .gnd(gnd), .vdd(vdd), .A(_9666_), .B(_9667_), .C(_9668_), .Y(_9669_) );
NAND2X1 NAND2X1_1231 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_2_), .B(micro_hash_ucr_3_pipe50_bF_buf4), .Y(_9670_) );
AOI21X1 AOI21X1_1720 ( .gnd(gnd), .vdd(vdd), .A(_9670_), .B(_9669_), .C(micro_hash_ucr_3_pipe51), .Y(_9671_) );
NOR2X1 NOR2X1_1578 ( .gnd(gnd), .vdd(vdd), .A(_9301__bF_buf0), .B(_9596_), .Y(_9672_) );
OAI21X1 OAI21X1_2716 ( .gnd(gnd), .vdd(vdd), .A(_9671_), .B(_9672_), .C(_9300__bF_buf0), .Y(_9673_) );
AOI21X1 AOI21X1_1721 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_2_), .B(micro_hash_ucr_3_pipe52_bF_buf1), .C(micro_hash_ucr_3_pipe53), .Y(_9674_) );
OAI21X1 OAI21X1_2717 ( .gnd(gnd), .vdd(vdd), .A(_9595_), .B(_9296_), .C(_9298__bF_buf1), .Y(_9675_) );
AOI21X1 AOI21X1_1722 ( .gnd(gnd), .vdd(vdd), .A(_9674_), .B(_9673_), .C(_9675_), .Y(_9676_) );
NOR2X1 NOR2X1_1579 ( .gnd(gnd), .vdd(vdd), .A(_8884_), .B(_9298__bF_buf0), .Y(_9677_) );
OAI21X1 OAI21X1_2718 ( .gnd(gnd), .vdd(vdd), .A(_9676_), .B(_9677_), .C(_9297_), .Y(_9678_) );
NAND2X1 NAND2X1_1232 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe55), .B(_9595_), .Y(_9679_) );
AOI21X1 AOI21X1_1723 ( .gnd(gnd), .vdd(vdd), .A(_9679_), .B(_9678_), .C(micro_hash_ucr_3_pipe56_bF_buf0), .Y(_9680_) );
OAI21X1 OAI21X1_2719 ( .gnd(gnd), .vdd(vdd), .A(_9680_), .B(_9591_), .C(_9295_), .Y(_9681_) );
NAND2X1 NAND2X1_1233 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe57_bF_buf0), .B(_9595_), .Y(_9682_) );
AOI21X1 AOI21X1_1724 ( .gnd(gnd), .vdd(vdd), .A(_9682_), .B(_9681_), .C(micro_hash_ucr_3_pipe58_bF_buf1), .Y(_9683_) );
OAI21X1 OAI21X1_2720 ( .gnd(gnd), .vdd(vdd), .A(_9683_), .B(_9590_), .C(_9290__bF_buf0), .Y(_9684_) );
NAND2X1 NAND2X1_1234 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe59), .B(_9595_), .Y(_9685_) );
AOI21X1 AOI21X1_1725 ( .gnd(gnd), .vdd(vdd), .A(_9685_), .B(_9684_), .C(micro_hash_ucr_3_pipe60_bF_buf0), .Y(_9686_) );
OAI21X1 OAI21X1_2721 ( .gnd(gnd), .vdd(vdd), .A(_9686_), .B(_9589_), .C(_9291_), .Y(_9687_) );
NAND2X1 NAND2X1_1235 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe61_bF_buf0), .B(_9595_), .Y(_9688_) );
AOI21X1 AOI21X1_1726 ( .gnd(gnd), .vdd(vdd), .A(_9688_), .B(_9687_), .C(micro_hash_ucr_3_pipe62_bF_buf0), .Y(_9689_) );
OAI21X1 OAI21X1_2722 ( .gnd(gnd), .vdd(vdd), .A(_9689_), .B(_9588_), .C(_9289__bF_buf0), .Y(_9690_) );
AOI21X1 AOI21X1_1727 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe63), .B(_9595_), .C(micro_hash_ucr_3_pipe64_bF_buf1), .Y(_9691_) );
OAI21X1 OAI21X1_2723 ( .gnd(gnd), .vdd(vdd), .A(_9288__bF_buf0), .B(micro_hash_ucr_3_a_2_), .C(_9284_), .Y(_9692_) );
AOI21X1 AOI21X1_1728 ( .gnd(gnd), .vdd(vdd), .A(_9691_), .B(_9690_), .C(_9692_), .Y(_9693_) );
OAI21X1 OAI21X1_2724 ( .gnd(gnd), .vdd(vdd), .A(_9596_), .B(_9284_), .C(_9286__bF_buf0), .Y(_9694_) );
OAI22X1 OAI22X1_114 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_2_), .B(_9286__bF_buf3), .C(_9693_), .D(_9694_), .Y(_9695_) );
NOR2X1 NOR2X1_1580 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe67), .B(_9695_), .Y(_9696_) );
NOR2X1 NOR2X1_1581 ( .gnd(gnd), .vdd(vdd), .A(_9285__bF_buf3), .B(_9596_), .Y(_9697_) );
OAI21X1 OAI21X1_2725 ( .gnd(gnd), .vdd(vdd), .A(_9696_), .B(_9697_), .C(_9282__bF_buf1), .Y(_9698_) );
AOI21X1 AOI21X1_1729 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_2_), .B(micro_hash_ucr_3_pipe68_bF_buf0), .C(micro_hash_ucr_3_pipe69), .Y(_9699_) );
OAI21X1 OAI21X1_2726 ( .gnd(gnd), .vdd(vdd), .A(_9595_), .B(_9283__bF_buf3), .C(_8705__bF_buf0), .Y(_9700_) );
AOI21X1 AOI21X1_1730 ( .gnd(gnd), .vdd(vdd), .A(_9699_), .B(_9698_), .C(_9700_), .Y(_8700__2_) );
INVX8 INVX8_269 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_3_bF_buf1_), .Y(_9701_) );
NAND2X1 NAND2X1_1236 ( .gnd(gnd), .vdd(vdd), .A(_9701__bF_buf3), .B(_8794_), .Y(_9702_) );
NAND2X1 NAND2X1_1237 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_3_bF_buf0_), .B(micro_hash_ucr_3_b_3_bF_buf1_), .Y(_9703_) );
NAND2X1 NAND2X1_1238 ( .gnd(gnd), .vdd(vdd), .A(_9703_), .B(_9702_), .Y(_9704_) );
INVX8 INVX8_270 ( .gnd(gnd), .vdd(vdd), .A(_9704_), .Y(_9705_) );
INVX8 INVX8_271 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_3_), .Y(_9706_) );
NAND2X1 NAND2X1_1239 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe58_bF_buf0), .B(_9706__bF_buf3), .Y(_9707_) );
NAND2X1 NAND2X1_1240 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe56_bF_buf4), .B(_9706__bF_buf2), .Y(_9708_) );
NAND2X1 NAND2X1_1241 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe24_bF_buf0), .B(_9706__bF_buf1), .Y(_9709_) );
NAND2X1 NAND2X1_1242 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe22_bF_buf3), .B(_9706__bF_buf0), .Y(_9710_) );
NAND2X1 NAND2X1_1243 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe20_bF_buf0), .B(_9706__bF_buf3), .Y(_9711_) );
NAND2X1 NAND2X1_1244 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe18_bF_buf3), .B(_9706__bF_buf2), .Y(_9712_) );
NAND2X1 NAND2X1_1245 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe17_bF_buf2), .B(_9705__bF_buf3), .Y(_9713_) );
NOR2X1 NOR2X1_1582 ( .gnd(gnd), .vdd(vdd), .A(_9706__bF_buf1), .B(_9336__bF_buf1), .Y(_9714_) );
NAND2X1 NAND2X1_1246 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe15_bF_buf0), .B(_9705__bF_buf2), .Y(_9715_) );
INVX2 INVX2_356 ( .gnd(gnd), .vdd(vdd), .A(_9617_), .Y(_9716_) );
NOR2X1 NOR2X1_1583 ( .gnd(gnd), .vdd(vdd), .A(_9610_), .B(_9716_), .Y(_9717_) );
NOR2X1 NOR2X1_1584 ( .gnd(gnd), .vdd(vdd), .A(H_3_3_), .B(micro_hash_ucr_3_pipe7), .Y(_9718_) );
AOI22X1 AOI22X1_68 ( .gnd(gnd), .vdd(vdd), .A(_9599_), .B(_9704_), .C(_9717_), .D(_9718_), .Y(_9719_) );
AOI21X1 AOI21X1_1731 ( .gnd(gnd), .vdd(vdd), .A(_9706__bF_buf0), .B(_9626_), .C(micro_hash_ucr_3_pipe15_bF_buf3), .Y(_9720_) );
OAI21X1 OAI21X1_2727 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe14_bF_buf3), .B(_9719_), .C(_9720_), .Y(_9721_) );
AOI21X1 AOI21X1_1732 ( .gnd(gnd), .vdd(vdd), .A(_9715_), .B(_9721_), .C(micro_hash_ucr_3_pipe16_bF_buf2), .Y(_9722_) );
OAI21X1 OAI21X1_2728 ( .gnd(gnd), .vdd(vdd), .A(_9722_), .B(_9714_), .C(_9332_), .Y(_9723_) );
NAND3X1 NAND3X1_479 ( .gnd(gnd), .vdd(vdd), .A(_9334__bF_buf0), .B(_9713_), .C(_9723_), .Y(_9724_) );
NAND3X1 NAND3X1_480 ( .gnd(gnd), .vdd(vdd), .A(_9333__bF_buf1), .B(_9712_), .C(_9724_), .Y(_9725_) );
NAND2X1 NAND2X1_1247 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe19), .B(_9705__bF_buf1), .Y(_9726_) );
NAND3X1 NAND3X1_481 ( .gnd(gnd), .vdd(vdd), .A(_9329__bF_buf4), .B(_9726_), .C(_9725_), .Y(_9727_) );
NAND3X1 NAND3X1_482 ( .gnd(gnd), .vdd(vdd), .A(_9331_), .B(_9711_), .C(_9727_), .Y(_9728_) );
NAND2X1 NAND2X1_1248 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe21_bF_buf2), .B(_9705__bF_buf0), .Y(_9729_) );
NAND3X1 NAND3X1_483 ( .gnd(gnd), .vdd(vdd), .A(_9330__bF_buf1), .B(_9729_), .C(_9728_), .Y(_9730_) );
NAND3X1 NAND3X1_484 ( .gnd(gnd), .vdd(vdd), .A(_9326__bF_buf2), .B(_9710_), .C(_9730_), .Y(_9731_) );
NAND2X1 NAND2X1_1249 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe23), .B(_9705__bF_buf3), .Y(_9732_) );
NAND3X1 NAND3X1_485 ( .gnd(gnd), .vdd(vdd), .A(_9328__bF_buf2), .B(_9732_), .C(_9731_), .Y(_9733_) );
NAND3X1 NAND3X1_486 ( .gnd(gnd), .vdd(vdd), .A(_9327_), .B(_9709_), .C(_9733_), .Y(_9734_) );
AOI21X1 AOI21X1_1733 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe25_bF_buf2), .B(_9705__bF_buf2), .C(micro_hash_ucr_3_pipe26_bF_buf4), .Y(_9735_) );
OAI21X1 OAI21X1_2729 ( .gnd(gnd), .vdd(vdd), .A(_9323__bF_buf3), .B(micro_hash_ucr_3_a_3_), .C(_9325__bF_buf2), .Y(_9736_) );
AOI21X1 AOI21X1_1734 ( .gnd(gnd), .vdd(vdd), .A(_9735_), .B(_9734_), .C(_9736_), .Y(_9737_) );
OAI21X1 OAI21X1_2730 ( .gnd(gnd), .vdd(vdd), .A(_9704_), .B(_9325__bF_buf1), .C(_9324__bF_buf1), .Y(_9738_) );
OAI22X1 OAI22X1_115 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_3_), .B(_9324__bF_buf0), .C(_9737_), .D(_9738_), .Y(_9739_) );
NAND2X1 NAND2X1_1250 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe29_bF_buf3), .B(_9705__bF_buf1), .Y(_9740_) );
OAI21X1 OAI21X1_2731 ( .gnd(gnd), .vdd(vdd), .A(_9739_), .B(micro_hash_ucr_3_pipe29_bF_buf2), .C(_9740_), .Y(_9741_) );
NAND2X1 NAND2X1_1251 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe30_bF_buf3), .B(_9706__bF_buf3), .Y(_9742_) );
OAI21X1 OAI21X1_2732 ( .gnd(gnd), .vdd(vdd), .A(_9741_), .B(micro_hash_ucr_3_pipe30_bF_buf2), .C(_9742_), .Y(_9743_) );
NAND2X1 NAND2X1_1252 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe31), .B(_9705__bF_buf0), .Y(_9744_) );
OAI21X1 OAI21X1_2733 ( .gnd(gnd), .vdd(vdd), .A(_9743_), .B(micro_hash_ucr_3_pipe31), .C(_9744_), .Y(_9745_) );
NAND2X1 NAND2X1_1253 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe32_bF_buf0), .B(_9706__bF_buf2), .Y(_9746_) );
OAI21X1 OAI21X1_2734 ( .gnd(gnd), .vdd(vdd), .A(_9745_), .B(micro_hash_ucr_3_pipe32_bF_buf3), .C(_9746_), .Y(_9747_) );
NAND2X1 NAND2X1_1254 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe33_bF_buf3), .B(_9705__bF_buf3), .Y(_9748_) );
OAI21X1 OAI21X1_2735 ( .gnd(gnd), .vdd(vdd), .A(_9747_), .B(micro_hash_ucr_3_pipe33_bF_buf2), .C(_9748_), .Y(_9749_) );
OAI21X1 OAI21X1_2736 ( .gnd(gnd), .vdd(vdd), .A(_9706__bF_buf1), .B(_9318__bF_buf1), .C(_9314_), .Y(_9750_) );
AOI21X1 AOI21X1_1735 ( .gnd(gnd), .vdd(vdd), .A(_9318__bF_buf0), .B(_9749_), .C(_9750_), .Y(_9751_) );
OAI21X1 OAI21X1_2737 ( .gnd(gnd), .vdd(vdd), .A(_9705__bF_buf2), .B(_9314_), .C(_9316__bF_buf1), .Y(_9752_) );
OAI22X1 OAI22X1_116 ( .gnd(gnd), .vdd(vdd), .A(_9706__bF_buf0), .B(_9316__bF_buf0), .C(_9751_), .D(_9752_), .Y(_9753_) );
OAI21X1 OAI21X1_2738 ( .gnd(gnd), .vdd(vdd), .A(_9704_), .B(_9315_), .C(_9311__bF_buf0), .Y(_9754_) );
AOI21X1 AOI21X1_1736 ( .gnd(gnd), .vdd(vdd), .A(_9315_), .B(_9753_), .C(_9754_), .Y(_9755_) );
OAI21X1 OAI21X1_2739 ( .gnd(gnd), .vdd(vdd), .A(_9311__bF_buf4), .B(micro_hash_ucr_3_a_3_), .C(_9313_), .Y(_9756_) );
AOI21X1 AOI21X1_1737 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe39_bF_buf1), .B(_9705__bF_buf1), .C(micro_hash_ucr_3_pipe40_bF_buf4), .Y(_9757_) );
OAI21X1 OAI21X1_2740 ( .gnd(gnd), .vdd(vdd), .A(_9755_), .B(_9756_), .C(_9757_), .Y(_9758_) );
OAI21X1 OAI21X1_2741 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_3_), .B(_9312__bF_buf0), .C(_9758_), .Y(_9759_) );
NAND2X1 NAND2X1_1255 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe41_bF_buf3), .B(_9705__bF_buf0), .Y(_9760_) );
OAI21X1 OAI21X1_2742 ( .gnd(gnd), .vdd(vdd), .A(_9759_), .B(micro_hash_ucr_3_pipe41_bF_buf2), .C(_9760_), .Y(_9761_) );
NAND2X1 NAND2X1_1256 ( .gnd(gnd), .vdd(vdd), .A(_9310__bF_buf0), .B(_9761_), .Y(_9762_) );
OAI21X1 OAI21X1_2743 ( .gnd(gnd), .vdd(vdd), .A(_9706__bF_buf3), .B(_9310__bF_buf4), .C(_9762_), .Y(_9763_) );
OAI21X1 OAI21X1_2744 ( .gnd(gnd), .vdd(vdd), .A(_9704_), .B(_9309__bF_buf1), .C(_9305__bF_buf1), .Y(_9764_) );
AOI21X1 AOI21X1_1738 ( .gnd(gnd), .vdd(vdd), .A(_9309__bF_buf0), .B(_9763_), .C(_9764_), .Y(_9765_) );
NOR2X1 NOR2X1_1585 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_3_), .B(_9305__bF_buf0), .Y(_9766_) );
OAI21X1 OAI21X1_2745 ( .gnd(gnd), .vdd(vdd), .A(_9765_), .B(_9766_), .C(_9307_), .Y(_9767_) );
NAND2X1 NAND2X1_1257 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe45_bF_buf0), .B(_9704_), .Y(_9768_) );
NAND3X1 NAND3X1_487 ( .gnd(gnd), .vdd(vdd), .A(_9306__bF_buf1), .B(_9768_), .C(_9767_), .Y(_9769_) );
AOI21X1 AOI21X1_1739 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_3_), .B(micro_hash_ucr_3_pipe46_bF_buf2), .C(micro_hash_ucr_3_pipe47), .Y(_9770_) );
OAI21X1 OAI21X1_2746 ( .gnd(gnd), .vdd(vdd), .A(_9705__bF_buf3), .B(_9302_), .C(_9304__bF_buf2), .Y(_9771_) );
AOI21X1 AOI21X1_1740 ( .gnd(gnd), .vdd(vdd), .A(_9770_), .B(_9769_), .C(_9771_), .Y(_9772_) );
NOR2X1 NOR2X1_1586 ( .gnd(gnd), .vdd(vdd), .A(_9706__bF_buf2), .B(_9304__bF_buf1), .Y(_9773_) );
OAI21X1 OAI21X1_2747 ( .gnd(gnd), .vdd(vdd), .A(_9772_), .B(_9773_), .C(_9303_), .Y(_9774_) );
AOI21X1 AOI21X1_1741 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe49_bF_buf3), .B(_9705__bF_buf2), .C(micro_hash_ucr_3_pipe50_bF_buf3), .Y(_9775_) );
OAI21X1 OAI21X1_2748 ( .gnd(gnd), .vdd(vdd), .A(_9299__bF_buf1), .B(micro_hash_ucr_3_a_3_), .C(_9301__bF_buf3), .Y(_9776_) );
AOI21X1 AOI21X1_1742 ( .gnd(gnd), .vdd(vdd), .A(_9775_), .B(_9774_), .C(_9776_), .Y(_9777_) );
OAI21X1 OAI21X1_2749 ( .gnd(gnd), .vdd(vdd), .A(_9704_), .B(_9301__bF_buf2), .C(_9300__bF_buf3), .Y(_9778_) );
OAI22X1 OAI22X1_117 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_3_), .B(_9300__bF_buf2), .C(_9777_), .D(_9778_), .Y(_9779_) );
OAI21X1 OAI21X1_2750 ( .gnd(gnd), .vdd(vdd), .A(_9705__bF_buf1), .B(_9296_), .C(_9298__bF_buf4), .Y(_9780_) );
AOI21X1 AOI21X1_1743 ( .gnd(gnd), .vdd(vdd), .A(_9296_), .B(_9779_), .C(_9780_), .Y(_9781_) );
NOR2X1 NOR2X1_1587 ( .gnd(gnd), .vdd(vdd), .A(_9706__bF_buf1), .B(_9298__bF_buf3), .Y(_9782_) );
OAI21X1 OAI21X1_2751 ( .gnd(gnd), .vdd(vdd), .A(_9781_), .B(_9782_), .C(_9297_), .Y(_9783_) );
NAND2X1 NAND2X1_1258 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe55), .B(_9705__bF_buf0), .Y(_9784_) );
NAND3X1 NAND3X1_488 ( .gnd(gnd), .vdd(vdd), .A(_9293__bF_buf0), .B(_9784_), .C(_9783_), .Y(_9785_) );
NAND3X1 NAND3X1_489 ( .gnd(gnd), .vdd(vdd), .A(_9295_), .B(_9708_), .C(_9785_), .Y(_9786_) );
NAND2X1 NAND2X1_1259 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe57_bF_buf3), .B(_9705__bF_buf3), .Y(_9787_) );
NAND3X1 NAND3X1_490 ( .gnd(gnd), .vdd(vdd), .A(_9294__bF_buf4), .B(_9787_), .C(_9786_), .Y(_9788_) );
NAND3X1 NAND3X1_491 ( .gnd(gnd), .vdd(vdd), .A(_9290__bF_buf3), .B(_9707_), .C(_9788_), .Y(_9789_) );
NAND2X1 NAND2X1_1260 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe59), .B(_9705__bF_buf2), .Y(_9790_) );
AOI21X1 AOI21X1_1744 ( .gnd(gnd), .vdd(vdd), .A(_9790_), .B(_9789_), .C(micro_hash_ucr_3_pipe60_bF_buf4), .Y(_9791_) );
OAI21X1 OAI21X1_2752 ( .gnd(gnd), .vdd(vdd), .A(_9706__bF_buf0), .B(_9292__bF_buf0), .C(_9291_), .Y(_9792_) );
OAI22X1 OAI22X1_118 ( .gnd(gnd), .vdd(vdd), .A(_9291_), .B(_9705__bF_buf1), .C(_9791_), .D(_9792_), .Y(_9793_) );
OAI21X1 OAI21X1_2753 ( .gnd(gnd), .vdd(vdd), .A(_9287__bF_buf0), .B(micro_hash_ucr_3_a_3_), .C(_9289__bF_buf3), .Y(_9794_) );
AOI21X1 AOI21X1_1745 ( .gnd(gnd), .vdd(vdd), .A(_9287__bF_buf4), .B(_9793_), .C(_9794_), .Y(_9795_) );
OAI21X1 OAI21X1_2754 ( .gnd(gnd), .vdd(vdd), .A(_9704_), .B(_9289__bF_buf2), .C(_9288__bF_buf3), .Y(_9796_) );
OAI22X1 OAI22X1_119 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_3_), .B(_9288__bF_buf2), .C(_9795_), .D(_9796_), .Y(_9797_) );
NAND2X1 NAND2X1_1261 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe65_bF_buf0), .B(_9705__bF_buf0), .Y(_9798_) );
OAI21X1 OAI21X1_2755 ( .gnd(gnd), .vdd(vdd), .A(_9797_), .B(micro_hash_ucr_3_pipe65_bF_buf3), .C(_9798_), .Y(_9799_) );
NAND2X1 NAND2X1_1262 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe66_bF_buf1), .B(_9706__bF_buf3), .Y(_9800_) );
OAI21X1 OAI21X1_2756 ( .gnd(gnd), .vdd(vdd), .A(_9799_), .B(micro_hash_ucr_3_pipe66_bF_buf0), .C(_9800_), .Y(_9801_) );
NAND2X1 NAND2X1_1263 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe67), .B(_9705__bF_buf3), .Y(_9802_) );
OAI21X1 OAI21X1_2757 ( .gnd(gnd), .vdd(vdd), .A(_9801_), .B(micro_hash_ucr_3_pipe67), .C(_9802_), .Y(_9803_) );
NAND2X1 NAND2X1_1264 ( .gnd(gnd), .vdd(vdd), .A(_9282__bF_buf0), .B(_9803_), .Y(_9804_) );
AOI21X1 AOI21X1_1746 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_3_), .B(micro_hash_ucr_3_pipe68_bF_buf3), .C(micro_hash_ucr_3_pipe69), .Y(_9805_) );
OAI21X1 OAI21X1_2758 ( .gnd(gnd), .vdd(vdd), .A(_9705__bF_buf2), .B(_9283__bF_buf2), .C(_8705__bF_buf13), .Y(_9806_) );
AOI21X1 AOI21X1_1747 ( .gnd(gnd), .vdd(vdd), .A(_9805_), .B(_9804_), .C(_9806_), .Y(_8700__3_) );
NAND2X1 NAND2X1_1265 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_4_), .B(micro_hash_ucr_3_pipe66_bF_buf4), .Y(_9807_) );
NAND2X1 NAND2X1_1266 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_4_), .B(micro_hash_ucr_3_pipe64_bF_buf0), .Y(_9808_) );
NAND2X1 NAND2X1_1267 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_4_), .B(micro_hash_ucr_3_pipe62_bF_buf3), .Y(_9809_) );
NAND2X1 NAND2X1_1268 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_4_), .B(micro_hash_ucr_3_pipe60_bF_buf3), .Y(_9810_) );
NAND2X1 NAND2X1_1269 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_4_), .B(micro_hash_ucr_3_pipe58_bF_buf3), .Y(_9811_) );
NAND2X1 NAND2X1_1270 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_4_), .B(micro_hash_ucr_3_pipe56_bF_buf3), .Y(_9812_) );
NAND2X1 NAND2X1_1271 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_4_), .B(micro_hash_ucr_3_pipe46_bF_buf1), .Y(_9813_) );
NAND2X1 NAND2X1_1272 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe34_bF_buf4), .B(_8903__bF_buf2), .Y(_9814_) );
NAND2X1 NAND2X1_1273 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe32_bF_buf2), .B(_8903__bF_buf1), .Y(_9815_) );
NAND2X1 NAND2X1_1274 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe30_bF_buf1), .B(_8903__bF_buf0), .Y(_9816_) );
NAND2X1 NAND2X1_1275 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe28_bF_buf4), .B(_8903__bF_buf3), .Y(_9817_) );
NAND2X1 NAND2X1_1276 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe26_bF_buf3), .B(_8903__bF_buf2), .Y(_9818_) );
NAND2X1 NAND2X1_1277 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe24_bF_buf4), .B(_8903__bF_buf1), .Y(_9819_) );
NAND2X1 NAND2X1_1278 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe22_bF_buf2), .B(_8903__bF_buf0), .Y(_9820_) );
NAND2X1 NAND2X1_1279 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe20_bF_buf4), .B(_8903__bF_buf3), .Y(_9821_) );
NOR2X1 NOR2X1_1588 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_4_), .B(micro_hash_ucr_3_b_4_bF_buf2_), .Y(_9822_) );
NAND2X1 NAND2X1_1280 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_4_), .B(micro_hash_ucr_3_b_4_bF_buf1_), .Y(_9823_) );
INVX4 INVX4_149 ( .gnd(gnd), .vdd(vdd), .A(_9823_), .Y(_9824_) );
OR2X2 OR2X2_69 ( .gnd(gnd), .vdd(vdd), .A(_9824_), .B(_9822_), .Y(_9825_) );
INVX8 INVX8_272 ( .gnd(gnd), .vdd(vdd), .A(_9825_), .Y(_9826_) );
NAND2X1 NAND2X1_1281 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe19), .B(_9826_), .Y(_9827_) );
NOR2X1 NOR2X1_1589 ( .gnd(gnd), .vdd(vdd), .A(_8903__bF_buf2), .B(_9334__bF_buf3), .Y(_9828_) );
INVX2 INVX2_357 ( .gnd(gnd), .vdd(vdd), .A(_9488_), .Y(_9829_) );
NAND2X1 NAND2X1_1282 ( .gnd(gnd), .vdd(vdd), .A(_9340_), .B(_9343_), .Y(_9830_) );
NOR2X1 NOR2X1_1590 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe7), .B(_9830_), .Y(_9831_) );
NOR2X1 NOR2X1_1591 ( .gnd(gnd), .vdd(vdd), .A(H_3_4_), .B(micro_hash_ucr_3_pipe14_bF_buf2), .Y(_9832_) );
AND2X2 AND2X2_683 ( .gnd(gnd), .vdd(vdd), .A(_9609_), .B(_9832_), .Y(_9833_) );
NAND3X1 NAND3X1_492 ( .gnd(gnd), .vdd(vdd), .A(_9829_), .B(_9833_), .C(_9831_), .Y(_9834_) );
OAI21X1 OAI21X1_2759 ( .gnd(gnd), .vdd(vdd), .A(_9625_), .B(micro_hash_ucr_3_a_4_), .C(_9834_), .Y(_9835_) );
AOI22X1 AOI22X1_69 ( .gnd(gnd), .vdd(vdd), .A(_8903__bF_buf1), .B(micro_hash_ucr_3_pipe14_bF_buf1), .C(_9835_), .D(_9339_), .Y(_9836_) );
AOI21X1 AOI21X1_1748 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe7), .B(_9341_), .C(micro_hash_ucr_3_pipe9), .Y(_9837_) );
OAI21X1 OAI21X1_2760 ( .gnd(gnd), .vdd(vdd), .A(_9837_), .B(micro_hash_ucr_3_pipe10_bF_buf1), .C(_9338_), .Y(_9838_) );
AOI21X1 AOI21X1_1749 ( .gnd(gnd), .vdd(vdd), .A(_9340_), .B(_9838_), .C(micro_hash_ucr_3_pipe13), .Y(_9839_) );
OAI21X1 OAI21X1_2761 ( .gnd(gnd), .vdd(vdd), .A(_9839_), .B(micro_hash_ucr_3_pipe14_bF_buf0), .C(_9337_), .Y(_9840_) );
AOI21X1 AOI21X1_1750 ( .gnd(gnd), .vdd(vdd), .A(_9825_), .B(_9840_), .C(micro_hash_ucr_3_pipe16_bF_buf1), .Y(_9841_) );
OAI21X1 OAI21X1_2762 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe15_bF_buf2), .B(_9836_), .C(_9841_), .Y(_9842_) );
AOI21X1 AOI21X1_1751 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_4_), .B(micro_hash_ucr_3_pipe16_bF_buf0), .C(micro_hash_ucr_3_pipe17_bF_buf1), .Y(_9843_) );
OAI21X1 OAI21X1_2763 ( .gnd(gnd), .vdd(vdd), .A(_9826_), .B(_9332_), .C(_9334__bF_buf2), .Y(_9844_) );
AOI21X1 AOI21X1_1752 ( .gnd(gnd), .vdd(vdd), .A(_9843_), .B(_9842_), .C(_9844_), .Y(_9845_) );
OAI21X1 OAI21X1_2764 ( .gnd(gnd), .vdd(vdd), .A(_9845_), .B(_9828_), .C(_9333__bF_buf0), .Y(_9846_) );
NAND3X1 NAND3X1_493 ( .gnd(gnd), .vdd(vdd), .A(_9329__bF_buf3), .B(_9827_), .C(_9846_), .Y(_9847_) );
NAND3X1 NAND3X1_494 ( .gnd(gnd), .vdd(vdd), .A(_9331_), .B(_9821_), .C(_9847_), .Y(_9848_) );
NAND2X1 NAND2X1_1283 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe21_bF_buf1), .B(_9826_), .Y(_9849_) );
NAND3X1 NAND3X1_495 ( .gnd(gnd), .vdd(vdd), .A(_9330__bF_buf0), .B(_9849_), .C(_9848_), .Y(_9850_) );
NAND3X1 NAND3X1_496 ( .gnd(gnd), .vdd(vdd), .A(_9326__bF_buf1), .B(_9820_), .C(_9850_), .Y(_9851_) );
NAND2X1 NAND2X1_1284 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe23), .B(_9826_), .Y(_9852_) );
NAND3X1 NAND3X1_497 ( .gnd(gnd), .vdd(vdd), .A(_9328__bF_buf1), .B(_9852_), .C(_9851_), .Y(_9853_) );
NAND3X1 NAND3X1_498 ( .gnd(gnd), .vdd(vdd), .A(_9327_), .B(_9819_), .C(_9853_), .Y(_9854_) );
NAND2X1 NAND2X1_1285 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe25_bF_buf1), .B(_9826_), .Y(_9855_) );
NAND3X1 NAND3X1_499 ( .gnd(gnd), .vdd(vdd), .A(_9323__bF_buf2), .B(_9855_), .C(_9854_), .Y(_9856_) );
NAND3X1 NAND3X1_500 ( .gnd(gnd), .vdd(vdd), .A(_9325__bF_buf0), .B(_9818_), .C(_9856_), .Y(_9857_) );
NAND2X1 NAND2X1_1286 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe27), .B(_9826_), .Y(_9858_) );
NAND3X1 NAND3X1_501 ( .gnd(gnd), .vdd(vdd), .A(_9324__bF_buf4), .B(_9858_), .C(_9857_), .Y(_9859_) );
NAND3X1 NAND3X1_502 ( .gnd(gnd), .vdd(vdd), .A(_9320_), .B(_9817_), .C(_9859_), .Y(_9860_) );
NAND2X1 NAND2X1_1287 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe29_bF_buf1), .B(_9826_), .Y(_9861_) );
NAND3X1 NAND3X1_503 ( .gnd(gnd), .vdd(vdd), .A(_9322__bF_buf1), .B(_9861_), .C(_9860_), .Y(_9862_) );
NAND3X1 NAND3X1_504 ( .gnd(gnd), .vdd(vdd), .A(_9321__bF_buf3), .B(_9816_), .C(_9862_), .Y(_9863_) );
NAND2X1 NAND2X1_1288 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe31), .B(_9826_), .Y(_9864_) );
NAND3X1 NAND3X1_505 ( .gnd(gnd), .vdd(vdd), .A(_9317__bF_buf4), .B(_9864_), .C(_9863_), .Y(_9865_) );
NAND3X1 NAND3X1_506 ( .gnd(gnd), .vdd(vdd), .A(_9319_), .B(_9815_), .C(_9865_), .Y(_9866_) );
NAND2X1 NAND2X1_1289 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe33_bF_buf1), .B(_9826_), .Y(_9867_) );
NAND3X1 NAND3X1_507 ( .gnd(gnd), .vdd(vdd), .A(_9318__bF_buf4), .B(_9867_), .C(_9866_), .Y(_9868_) );
NAND3X1 NAND3X1_508 ( .gnd(gnd), .vdd(vdd), .A(_9314_), .B(_9814_), .C(_9868_), .Y(_9869_) );
AOI21X1 AOI21X1_1753 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe35_bF_buf3), .B(_9826_), .C(micro_hash_ucr_3_pipe36_bF_buf3), .Y(_9870_) );
OAI21X1 OAI21X1_2765 ( .gnd(gnd), .vdd(vdd), .A(_9316__bF_buf3), .B(micro_hash_ucr_3_a_4_), .C(_9315_), .Y(_9871_) );
AOI21X1 AOI21X1_1754 ( .gnd(gnd), .vdd(vdd), .A(_9870_), .B(_9869_), .C(_9871_), .Y(_9872_) );
OAI21X1 OAI21X1_2766 ( .gnd(gnd), .vdd(vdd), .A(_9825_), .B(_9315_), .C(_9311__bF_buf3), .Y(_9873_) );
OAI22X1 OAI22X1_120 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_4_), .B(_9311__bF_buf2), .C(_9872_), .D(_9873_), .Y(_9874_) );
NAND2X1 NAND2X1_1290 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe39_bF_buf0), .B(_9826_), .Y(_9875_) );
OAI21X1 OAI21X1_2767 ( .gnd(gnd), .vdd(vdd), .A(_9874_), .B(micro_hash_ucr_3_pipe39_bF_buf3), .C(_9875_), .Y(_9876_) );
NAND2X1 NAND2X1_1291 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe40_bF_buf3), .B(_8903__bF_buf0), .Y(_9877_) );
OAI21X1 OAI21X1_2768 ( .gnd(gnd), .vdd(vdd), .A(_9876_), .B(micro_hash_ucr_3_pipe40_bF_buf2), .C(_9877_), .Y(_9878_) );
NAND2X1 NAND2X1_1292 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe41_bF_buf1), .B(_9826_), .Y(_9879_) );
OAI21X1 OAI21X1_2769 ( .gnd(gnd), .vdd(vdd), .A(_9878_), .B(micro_hash_ucr_3_pipe41_bF_buf0), .C(_9879_), .Y(_9880_) );
OAI21X1 OAI21X1_2770 ( .gnd(gnd), .vdd(vdd), .A(_8903__bF_buf3), .B(_9310__bF_buf3), .C(_9309__bF_buf3), .Y(_9881_) );
AOI21X1 AOI21X1_1755 ( .gnd(gnd), .vdd(vdd), .A(_9310__bF_buf2), .B(_9880_), .C(_9881_), .Y(_9882_) );
OAI21X1 OAI21X1_2771 ( .gnd(gnd), .vdd(vdd), .A(_9826_), .B(_9309__bF_buf2), .C(_9305__bF_buf4), .Y(_9883_) );
OAI22X1 OAI22X1_121 ( .gnd(gnd), .vdd(vdd), .A(_8903__bF_buf2), .B(_9305__bF_buf3), .C(_9882_), .D(_9883_), .Y(_9884_) );
OAI21X1 OAI21X1_2772 ( .gnd(gnd), .vdd(vdd), .A(_9824_), .B(_9822_), .C(micro_hash_ucr_3_pipe45_bF_buf3), .Y(_9885_) );
OAI21X1 OAI21X1_2773 ( .gnd(gnd), .vdd(vdd), .A(_9884_), .B(micro_hash_ucr_3_pipe45_bF_buf2), .C(_9885_), .Y(_9886_) );
OAI21X1 OAI21X1_2774 ( .gnd(gnd), .vdd(vdd), .A(_9886_), .B(micro_hash_ucr_3_pipe46_bF_buf0), .C(_9813_), .Y(_9887_) );
OAI21X1 OAI21X1_2775 ( .gnd(gnd), .vdd(vdd), .A(_9825_), .B(_9302_), .C(_9304__bF_buf0), .Y(_9888_) );
AOI21X1 AOI21X1_1756 ( .gnd(gnd), .vdd(vdd), .A(_9302_), .B(_9887_), .C(_9888_), .Y(_9889_) );
OAI21X1 OAI21X1_2776 ( .gnd(gnd), .vdd(vdd), .A(_9304__bF_buf3), .B(micro_hash_ucr_3_a_4_), .C(_9303_), .Y(_9890_) );
AOI21X1 AOI21X1_1757 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe49_bF_buf2), .B(_9826_), .C(micro_hash_ucr_3_pipe50_bF_buf2), .Y(_9891_) );
OAI21X1 OAI21X1_2777 ( .gnd(gnd), .vdd(vdd), .A(_9889_), .B(_9890_), .C(_9891_), .Y(_9892_) );
NAND2X1 NAND2X1_1293 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe50_bF_buf1), .B(_8903__bF_buf1), .Y(_9893_) );
NAND3X1 NAND3X1_509 ( .gnd(gnd), .vdd(vdd), .A(_9301__bF_buf1), .B(_9893_), .C(_9892_), .Y(_9894_) );
NAND2X1 NAND2X1_1294 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe51), .B(_9826_), .Y(_9895_) );
AOI21X1 AOI21X1_1758 ( .gnd(gnd), .vdd(vdd), .A(_9895_), .B(_9894_), .C(micro_hash_ucr_3_pipe52_bF_buf0), .Y(_9896_) );
OAI21X1 OAI21X1_2778 ( .gnd(gnd), .vdd(vdd), .A(_8903__bF_buf0), .B(_9300__bF_buf1), .C(_9296_), .Y(_9897_) );
AOI21X1 AOI21X1_1759 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe53), .B(_9825_), .C(micro_hash_ucr_3_pipe54_bF_buf0), .Y(_9898_) );
OAI21X1 OAI21X1_2779 ( .gnd(gnd), .vdd(vdd), .A(_9896_), .B(_9897_), .C(_9898_), .Y(_9899_) );
NAND2X1 NAND2X1_1295 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_4_), .B(micro_hash_ucr_3_pipe54_bF_buf3), .Y(_9900_) );
NAND3X1 NAND3X1_510 ( .gnd(gnd), .vdd(vdd), .A(_9297_), .B(_9900_), .C(_9899_), .Y(_9901_) );
OAI21X1 OAI21X1_2780 ( .gnd(gnd), .vdd(vdd), .A(_9824_), .B(_9822_), .C(micro_hash_ucr_3_pipe55), .Y(_9902_) );
NAND3X1 NAND3X1_511 ( .gnd(gnd), .vdd(vdd), .A(_9293__bF_buf3), .B(_9902_), .C(_9901_), .Y(_9903_) );
NAND3X1 NAND3X1_512 ( .gnd(gnd), .vdd(vdd), .A(_9295_), .B(_9812_), .C(_9903_), .Y(_9904_) );
OAI21X1 OAI21X1_2781 ( .gnd(gnd), .vdd(vdd), .A(_9824_), .B(_9822_), .C(micro_hash_ucr_3_pipe57_bF_buf2), .Y(_9905_) );
NAND3X1 NAND3X1_513 ( .gnd(gnd), .vdd(vdd), .A(_9294__bF_buf3), .B(_9905_), .C(_9904_), .Y(_9906_) );
NAND3X1 NAND3X1_514 ( .gnd(gnd), .vdd(vdd), .A(_9290__bF_buf2), .B(_9811_), .C(_9906_), .Y(_9907_) );
OAI21X1 OAI21X1_2782 ( .gnd(gnd), .vdd(vdd), .A(_9824_), .B(_9822_), .C(micro_hash_ucr_3_pipe59), .Y(_9908_) );
NAND3X1 NAND3X1_515 ( .gnd(gnd), .vdd(vdd), .A(_9292__bF_buf3), .B(_9908_), .C(_9907_), .Y(_9909_) );
NAND3X1 NAND3X1_516 ( .gnd(gnd), .vdd(vdd), .A(_9291_), .B(_9810_), .C(_9909_), .Y(_9910_) );
OAI21X1 OAI21X1_2783 ( .gnd(gnd), .vdd(vdd), .A(_9824_), .B(_9822_), .C(micro_hash_ucr_3_pipe61_bF_buf3), .Y(_9911_) );
NAND3X1 NAND3X1_517 ( .gnd(gnd), .vdd(vdd), .A(_9287__bF_buf3), .B(_9911_), .C(_9910_), .Y(_9912_) );
NAND3X1 NAND3X1_518 ( .gnd(gnd), .vdd(vdd), .A(_9289__bF_buf1), .B(_9809_), .C(_9912_), .Y(_9913_) );
OAI21X1 OAI21X1_2784 ( .gnd(gnd), .vdd(vdd), .A(_9824_), .B(_9822_), .C(micro_hash_ucr_3_pipe63), .Y(_9914_) );
NAND3X1 NAND3X1_519 ( .gnd(gnd), .vdd(vdd), .A(_9288__bF_buf1), .B(_9914_), .C(_9913_), .Y(_9915_) );
NAND3X1 NAND3X1_520 ( .gnd(gnd), .vdd(vdd), .A(_9284_), .B(_9808_), .C(_9915_), .Y(_9916_) );
OAI21X1 OAI21X1_2785 ( .gnd(gnd), .vdd(vdd), .A(_9824_), .B(_9822_), .C(micro_hash_ucr_3_pipe65_bF_buf2), .Y(_9917_) );
NAND3X1 NAND3X1_521 ( .gnd(gnd), .vdd(vdd), .A(_9286__bF_buf2), .B(_9917_), .C(_9916_), .Y(_9918_) );
NAND3X1 NAND3X1_522 ( .gnd(gnd), .vdd(vdd), .A(_9285__bF_buf2), .B(_9807_), .C(_9918_), .Y(_9919_) );
OAI21X1 OAI21X1_2786 ( .gnd(gnd), .vdd(vdd), .A(_9824_), .B(_9822_), .C(micro_hash_ucr_3_pipe67), .Y(_9920_) );
NAND3X1 NAND3X1_523 ( .gnd(gnd), .vdd(vdd), .A(_9282__bF_buf4), .B(_9920_), .C(_9919_), .Y(_9921_) );
AOI21X1 AOI21X1_1760 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_4_), .B(micro_hash_ucr_3_pipe68_bF_buf2), .C(micro_hash_ucr_3_pipe69), .Y(_9922_) );
OAI21X1 OAI21X1_2787 ( .gnd(gnd), .vdd(vdd), .A(_9826_), .B(_9283__bF_buf1), .C(_8705__bF_buf12), .Y(_9923_) );
AOI21X1 AOI21X1_1761 ( .gnd(gnd), .vdd(vdd), .A(_9922_), .B(_9921_), .C(_9923_), .Y(_8700__4_) );
NAND2X1 NAND2X1_1296 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_5_bF_buf1_), .B(micro_hash_ucr_3_pipe62_bF_buf2), .Y(_9924_) );
NOR2X1 NOR2X1_1592 ( .gnd(gnd), .vdd(vdd), .A(_8909_), .B(_9293__bF_buf2), .Y(_9925_) );
NOR2X1 NOR2X1_1593 ( .gnd(gnd), .vdd(vdd), .A(_8909_), .B(_9298__bF_buf2), .Y(_9926_) );
NOR2X1 NOR2X1_1594 ( .gnd(gnd), .vdd(vdd), .A(_8909_), .B(_9300__bF_buf0), .Y(_9927_) );
NOR2X1 NOR2X1_1595 ( .gnd(gnd), .vdd(vdd), .A(_8909_), .B(_9299__bF_buf0), .Y(_9928_) );
NAND2X1 NAND2X1_1297 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_5_bF_buf0_), .B(micro_hash_ucr_3_pipe40_bF_buf1), .Y(_9929_) );
NAND2X1 NAND2X1_1298 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_5_bF_buf3_), .B(micro_hash_ucr_3_pipe38_bF_buf3), .Y(_9930_) );
NAND2X1 NAND2X1_1299 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_5_bF_buf2_), .B(micro_hash_ucr_3_pipe36_bF_buf2), .Y(_9931_) );
INVX1 INVX1_626 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_5_), .Y(_9932_) );
NAND2X1 NAND2X1_1300 ( .gnd(gnd), .vdd(vdd), .A(_9932_), .B(_8814__bF_buf2), .Y(_9933_) );
NAND2X1 NAND2X1_1301 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_5_), .B(micro_hash_ucr_3_b_5_bF_buf1_), .Y(_9934_) );
NAND2X1 NAND2X1_1302 ( .gnd(gnd), .vdd(vdd), .A(_9934_), .B(_9933_), .Y(_9935_) );
INVX8 INVX8_273 ( .gnd(gnd), .vdd(vdd), .A(_9935_), .Y(_9936_) );
NOR2X1 NOR2X1_1596 ( .gnd(gnd), .vdd(vdd), .A(_8909_), .B(_9330__bF_buf4), .Y(_9937_) );
NAND2X1 NAND2X1_1303 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe21_bF_buf0), .B(_9936_), .Y(_9938_) );
NOR2X1 NOR2X1_1597 ( .gnd(gnd), .vdd(vdd), .A(_8909_), .B(_9329__bF_buf2), .Y(_9939_) );
NOR2X1 NOR2X1_1598 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_5_bF_buf1_), .B(_9627_), .Y(_9940_) );
INVX1 INVX1_627 ( .gnd(gnd), .vdd(vdd), .A(_9717_), .Y(_9941_) );
NOR2X1 NOR2X1_1599 ( .gnd(gnd), .vdd(vdd), .A(H_3_5_), .B(micro_hash_ucr_3_pipe14_bF_buf3), .Y(_9942_) );
NAND3X1 NAND3X1_524 ( .gnd(gnd), .vdd(vdd), .A(_9344_), .B(_9620_), .C(_9942_), .Y(_9943_) );
NOR2X1 NOR2X1_1600 ( .gnd(gnd), .vdd(vdd), .A(_9943_), .B(_9941_), .Y(_9944_) );
OAI21X1 OAI21X1_2788 ( .gnd(gnd), .vdd(vdd), .A(_9940_), .B(_9944_), .C(_9332_), .Y(_9945_) );
AND2X2 AND2X2_684 ( .gnd(gnd), .vdd(vdd), .A(_9945_), .B(_9334__bF_buf1), .Y(_9946_) );
OAI21X1 OAI21X1_2789 ( .gnd(gnd), .vdd(vdd), .A(_9602_), .B(_9936_), .C(_9946_), .Y(_9947_) );
AOI21X1 AOI21X1_1762 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_5_bF_buf0_), .B(micro_hash_ucr_3_pipe18_bF_buf2), .C(micro_hash_ucr_3_pipe19), .Y(_9948_) );
OAI21X1 OAI21X1_2790 ( .gnd(gnd), .vdd(vdd), .A(_9936_), .B(_9333__bF_buf3), .C(_9329__bF_buf1), .Y(_9949_) );
AOI21X1 AOI21X1_1763 ( .gnd(gnd), .vdd(vdd), .A(_9948_), .B(_9947_), .C(_9949_), .Y(_9950_) );
OAI21X1 OAI21X1_2791 ( .gnd(gnd), .vdd(vdd), .A(_9950_), .B(_9939_), .C(_9331_), .Y(_9951_) );
AOI21X1 AOI21X1_1764 ( .gnd(gnd), .vdd(vdd), .A(_9938_), .B(_9951_), .C(micro_hash_ucr_3_pipe22_bF_buf1), .Y(_9952_) );
OAI21X1 OAI21X1_2792 ( .gnd(gnd), .vdd(vdd), .A(_9952_), .B(_9937_), .C(_9326__bF_buf0), .Y(_9953_) );
AOI21X1 AOI21X1_1765 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe23), .B(_9936_), .C(micro_hash_ucr_3_pipe24_bF_buf3), .Y(_9954_) );
OAI21X1 OAI21X1_2793 ( .gnd(gnd), .vdd(vdd), .A(_9328__bF_buf0), .B(micro_hash_ucr_3_a_5_bF_buf3_), .C(_9327_), .Y(_9955_) );
AOI21X1 AOI21X1_1766 ( .gnd(gnd), .vdd(vdd), .A(_9954_), .B(_9953_), .C(_9955_), .Y(_9956_) );
OAI21X1 OAI21X1_2794 ( .gnd(gnd), .vdd(vdd), .A(_9935_), .B(_9327_), .C(_9323__bF_buf1), .Y(_9957_) );
OAI22X1 OAI22X1_122 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_5_bF_buf2_), .B(_9323__bF_buf0), .C(_9956_), .D(_9957_), .Y(_9958_) );
OAI21X1 OAI21X1_2795 ( .gnd(gnd), .vdd(vdd), .A(_9936_), .B(_9325__bF_buf3), .C(_9324__bF_buf3), .Y(_9959_) );
AOI21X1 AOI21X1_1767 ( .gnd(gnd), .vdd(vdd), .A(_9325__bF_buf2), .B(_9958_), .C(_9959_), .Y(_9960_) );
NOR2X1 NOR2X1_1601 ( .gnd(gnd), .vdd(vdd), .A(_8909_), .B(_9324__bF_buf2), .Y(_9961_) );
OAI21X1 OAI21X1_2796 ( .gnd(gnd), .vdd(vdd), .A(_9960_), .B(_9961_), .C(_9320_), .Y(_9962_) );
AOI21X1 AOI21X1_1768 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe29_bF_buf0), .B(_9936_), .C(micro_hash_ucr_3_pipe30_bF_buf0), .Y(_9963_) );
OAI21X1 OAI21X1_2797 ( .gnd(gnd), .vdd(vdd), .A(_9322__bF_buf0), .B(micro_hash_ucr_3_a_5_bF_buf1_), .C(_9321__bF_buf2), .Y(_9964_) );
AOI21X1 AOI21X1_1769 ( .gnd(gnd), .vdd(vdd), .A(_9963_), .B(_9962_), .C(_9964_), .Y(_9965_) );
OAI21X1 OAI21X1_2798 ( .gnd(gnd), .vdd(vdd), .A(_9935_), .B(_9321__bF_buf1), .C(_9317__bF_buf3), .Y(_9966_) );
OAI22X1 OAI22X1_123 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_5_bF_buf0_), .B(_9317__bF_buf2), .C(_9965_), .D(_9966_), .Y(_9967_) );
NAND2X1 NAND2X1_1304 ( .gnd(gnd), .vdd(vdd), .A(_9319_), .B(_9967_), .Y(_9968_) );
OAI21X1 OAI21X1_2799 ( .gnd(gnd), .vdd(vdd), .A(_9319_), .B(_9936_), .C(_9968_), .Y(_9969_) );
NAND2X1 NAND2X1_1305 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_5_bF_buf3_), .B(micro_hash_ucr_3_pipe34_bF_buf3), .Y(_9970_) );
OAI21X1 OAI21X1_2800 ( .gnd(gnd), .vdd(vdd), .A(_9969_), .B(micro_hash_ucr_3_pipe34_bF_buf2), .C(_9970_), .Y(_9971_) );
NAND2X1 NAND2X1_1306 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe35_bF_buf2), .B(_9935_), .Y(_9972_) );
OAI21X1 OAI21X1_2801 ( .gnd(gnd), .vdd(vdd), .A(_9971_), .B(micro_hash_ucr_3_pipe35_bF_buf1), .C(_9972_), .Y(_9973_) );
OAI21X1 OAI21X1_2802 ( .gnd(gnd), .vdd(vdd), .A(_9973_), .B(micro_hash_ucr_3_pipe36_bF_buf1), .C(_9931_), .Y(_9974_) );
NAND2X1 NAND2X1_1307 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe37_bF_buf2), .B(_9935_), .Y(_9975_) );
OAI21X1 OAI21X1_2803 ( .gnd(gnd), .vdd(vdd), .A(_9974_), .B(micro_hash_ucr_3_pipe37_bF_buf1), .C(_9975_), .Y(_9976_) );
OAI21X1 OAI21X1_2804 ( .gnd(gnd), .vdd(vdd), .A(_9976_), .B(micro_hash_ucr_3_pipe38_bF_buf2), .C(_9930_), .Y(_9977_) );
NAND2X1 NAND2X1_1308 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe39_bF_buf2), .B(_9935_), .Y(_9978_) );
OAI21X1 OAI21X1_2805 ( .gnd(gnd), .vdd(vdd), .A(_9977_), .B(micro_hash_ucr_3_pipe39_bF_buf1), .C(_9978_), .Y(_9979_) );
OAI21X1 OAI21X1_2806 ( .gnd(gnd), .vdd(vdd), .A(_9979_), .B(micro_hash_ucr_3_pipe40_bF_buf0), .C(_9929_), .Y(_9980_) );
NAND2X1 NAND2X1_1309 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe41_bF_buf3), .B(_9935_), .Y(_9981_) );
OAI21X1 OAI21X1_2807 ( .gnd(gnd), .vdd(vdd), .A(_9980_), .B(micro_hash_ucr_3_pipe41_bF_buf2), .C(_9981_), .Y(_9982_) );
NOR2X1 NOR2X1_1602 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe42_bF_buf3), .B(_9982_), .Y(_9983_) );
OAI21X1 OAI21X1_2808 ( .gnd(gnd), .vdd(vdd), .A(_8909_), .B(_9310__bF_buf1), .C(_9309__bF_buf1), .Y(_9984_) );
AOI21X1 AOI21X1_1770 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe43), .B(_9935_), .C(micro_hash_ucr_3_pipe44_bF_buf2), .Y(_9985_) );
OAI21X1 OAI21X1_2809 ( .gnd(gnd), .vdd(vdd), .A(_9983_), .B(_9984_), .C(_9985_), .Y(_9986_) );
NAND2X1 NAND2X1_1310 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_5_bF_buf2_), .B(micro_hash_ucr_3_pipe44_bF_buf1), .Y(_9987_) );
AOI21X1 AOI21X1_1771 ( .gnd(gnd), .vdd(vdd), .A(_9987_), .B(_9986_), .C(micro_hash_ucr_3_pipe45_bF_buf1), .Y(_9988_) );
NOR2X1 NOR2X1_1603 ( .gnd(gnd), .vdd(vdd), .A(_9307_), .B(_9935_), .Y(_9989_) );
OAI21X1 OAI21X1_2810 ( .gnd(gnd), .vdd(vdd), .A(_9988_), .B(_9989_), .C(_9306__bF_buf0), .Y(_9990_) );
AOI21X1 AOI21X1_1772 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_5_bF_buf1_), .B(micro_hash_ucr_3_pipe46_bF_buf4), .C(micro_hash_ucr_3_pipe47), .Y(_9991_) );
OAI21X1 OAI21X1_2811 ( .gnd(gnd), .vdd(vdd), .A(_9936_), .B(_9302_), .C(_9304__bF_buf2), .Y(_9992_) );
AOI21X1 AOI21X1_1773 ( .gnd(gnd), .vdd(vdd), .A(_9991_), .B(_9990_), .C(_9992_), .Y(_9993_) );
NOR2X1 NOR2X1_1604 ( .gnd(gnd), .vdd(vdd), .A(_8909_), .B(_9304__bF_buf1), .Y(_9994_) );
OAI21X1 OAI21X1_2812 ( .gnd(gnd), .vdd(vdd), .A(_9993_), .B(_9994_), .C(_9303_), .Y(_9995_) );
NAND2X1 NAND2X1_1311 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe49_bF_buf1), .B(_9936_), .Y(_9996_) );
AOI21X1 AOI21X1_1774 ( .gnd(gnd), .vdd(vdd), .A(_9996_), .B(_9995_), .C(micro_hash_ucr_3_pipe50_bF_buf0), .Y(_9997_) );
OAI21X1 OAI21X1_2813 ( .gnd(gnd), .vdd(vdd), .A(_9997_), .B(_9928_), .C(_9301__bF_buf0), .Y(_9998_) );
NAND2X1 NAND2X1_1312 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe51), .B(_9936_), .Y(_9999_) );
AOI21X1 AOI21X1_1775 ( .gnd(gnd), .vdd(vdd), .A(_9999_), .B(_9998_), .C(micro_hash_ucr_3_pipe52_bF_buf4), .Y(_10000_) );
OAI21X1 OAI21X1_2814 ( .gnd(gnd), .vdd(vdd), .A(_10000_), .B(_9927_), .C(_9296_), .Y(_10001_) );
NAND2X1 NAND2X1_1313 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe53), .B(_9936_), .Y(_10002_) );
AOI21X1 AOI21X1_1776 ( .gnd(gnd), .vdd(vdd), .A(_10002_), .B(_10001_), .C(micro_hash_ucr_3_pipe54_bF_buf2), .Y(_10003_) );
OAI21X1 OAI21X1_2815 ( .gnd(gnd), .vdd(vdd), .A(_10003_), .B(_9926_), .C(_9297_), .Y(_10004_) );
NAND2X1 NAND2X1_1314 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe55), .B(_9936_), .Y(_10005_) );
AOI21X1 AOI21X1_1777 ( .gnd(gnd), .vdd(vdd), .A(_10005_), .B(_10004_), .C(micro_hash_ucr_3_pipe56_bF_buf2), .Y(_10006_) );
OAI21X1 OAI21X1_2816 ( .gnd(gnd), .vdd(vdd), .A(_10006_), .B(_9925_), .C(_9295_), .Y(_10007_) );
AOI21X1 AOI21X1_1778 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe57_bF_buf1), .B(_9936_), .C(micro_hash_ucr_3_pipe58_bF_buf2), .Y(_10008_) );
OAI21X1 OAI21X1_2817 ( .gnd(gnd), .vdd(vdd), .A(_9294__bF_buf2), .B(micro_hash_ucr_3_a_5_bF_buf0_), .C(_9290__bF_buf1), .Y(_10009_) );
AOI21X1 AOI21X1_1779 ( .gnd(gnd), .vdd(vdd), .A(_10008_), .B(_10007_), .C(_10009_), .Y(_10010_) );
OAI21X1 OAI21X1_2818 ( .gnd(gnd), .vdd(vdd), .A(_9935_), .B(_9290__bF_buf0), .C(_9292__bF_buf2), .Y(_10011_) );
OAI22X1 OAI22X1_124 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_5_bF_buf3_), .B(_9292__bF_buf1), .C(_10010_), .D(_10011_), .Y(_10012_) );
NOR2X1 NOR2X1_1605 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe61_bF_buf2), .B(_10012_), .Y(_10013_) );
NOR2X1 NOR2X1_1606 ( .gnd(gnd), .vdd(vdd), .A(_9291_), .B(_9935_), .Y(_10014_) );
OAI21X1 OAI21X1_2819 ( .gnd(gnd), .vdd(vdd), .A(_10013_), .B(_10014_), .C(_9287__bF_buf2), .Y(_10015_) );
AOI21X1 AOI21X1_1780 ( .gnd(gnd), .vdd(vdd), .A(_9924_), .B(_10015_), .C(micro_hash_ucr_3_pipe63), .Y(_10016_) );
OAI21X1 OAI21X1_2820 ( .gnd(gnd), .vdd(vdd), .A(_9935_), .B(_9289__bF_buf0), .C(_9288__bF_buf0), .Y(_10017_) );
AOI21X1 AOI21X1_1781 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe64_bF_buf4), .B(_8909_), .C(micro_hash_ucr_3_pipe65_bF_buf1), .Y(_10018_) );
OAI21X1 OAI21X1_2821 ( .gnd(gnd), .vdd(vdd), .A(_10016_), .B(_10017_), .C(_10018_), .Y(_10019_) );
AOI21X1 AOI21X1_1782 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe65_bF_buf0), .B(_9936_), .C(micro_hash_ucr_3_pipe66_bF_buf3), .Y(_10020_) );
AOI22X1 AOI22X1_70 ( .gnd(gnd), .vdd(vdd), .A(_8909_), .B(micro_hash_ucr_3_pipe66_bF_buf2), .C(_10019_), .D(_10020_), .Y(_10021_) );
AOI21X1 AOI21X1_1783 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe67), .B(_9935_), .C(micro_hash_ucr_3_pipe68_bF_buf1), .Y(_10022_) );
OAI21X1 OAI21X1_2822 ( .gnd(gnd), .vdd(vdd), .A(_10021_), .B(micro_hash_ucr_3_pipe67), .C(_10022_), .Y(_10023_) );
AOI21X1 AOI21X1_1784 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_5_bF_buf2_), .B(micro_hash_ucr_3_pipe68_bF_buf0), .C(micro_hash_ucr_3_pipe69), .Y(_10024_) );
OAI21X1 OAI21X1_2823 ( .gnd(gnd), .vdd(vdd), .A(_9936_), .B(_9283__bF_buf0), .C(_8705__bF_buf11), .Y(_10025_) );
AOI21X1 AOI21X1_1785 ( .gnd(gnd), .vdd(vdd), .A(_10024_), .B(_10023_), .C(_10025_), .Y(_8700__5_) );
NAND2X1 NAND2X1_1315 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_6_bF_buf1_), .B(micro_hash_ucr_3_pipe54_bF_buf1), .Y(_10026_) );
NAND2X1 NAND2X1_1316 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_6_bF_buf0_), .B(micro_hash_ucr_3_pipe52_bF_buf3), .Y(_10027_) );
NAND2X1 NAND2X1_1317 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_6_bF_buf3_), .B(micro_hash_ucr_3_pipe50_bF_buf4), .Y(_10028_) );
NAND2X1 NAND2X1_1318 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_6_bF_buf2_), .B(micro_hash_ucr_3_pipe48_bF_buf1), .Y(_10029_) );
NAND2X1 NAND2X1_1319 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_6_bF_buf1_), .B(micro_hash_ucr_3_pipe46_bF_buf3), .Y(_10030_) );
NAND2X1 NAND2X1_1320 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_6_bF_buf0_), .B(micro_hash_ucr_3_pipe44_bF_buf0), .Y(_10031_) );
NAND2X1 NAND2X1_1321 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_6_bF_buf3_), .B(micro_hash_ucr_3_pipe42_bF_buf2), .Y(_10032_) );
NAND2X1 NAND2X1_1322 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_6_bF_buf2_), .B(micro_hash_ucr_3_pipe40_bF_buf4), .Y(_10033_) );
NAND2X1 NAND2X1_1323 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_6_bF_buf1_), .B(micro_hash_ucr_3_pipe38_bF_buf1), .Y(_10034_) );
NOR2X1 NOR2X1_1607 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_6_), .B(micro_hash_ucr_3_b_6_bF_buf1_), .Y(_10035_) );
NOR2X1 NOR2X1_1608 ( .gnd(gnd), .vdd(vdd), .A(_12893_), .B(_8828_), .Y(_10036_) );
NOR2X1 NOR2X1_1609 ( .gnd(gnd), .vdd(vdd), .A(_10035_), .B(_10036_), .Y(_10037_) );
INVX4 INVX4_150 ( .gnd(gnd), .vdd(vdd), .A(_10037_), .Y(_10038_) );
NAND2X1 NAND2X1_1324 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe26_bF_buf2), .B(_8923_), .Y(_10039_) );
OAI21X1 OAI21X1_2824 ( .gnd(gnd), .vdd(vdd), .A(_10038_), .B(_9339_), .C(_9335__bF_buf2), .Y(_10040_) );
OR2X2 OR2X2_70 ( .gnd(gnd), .vdd(vdd), .A(_9625_), .B(micro_hash_ucr_3_a_6_bF_buf0_), .Y(_10041_) );
NOR2X1 NOR2X1_1610 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe11), .B(micro_hash_ucr_3_pipe7), .Y(_10042_) );
NAND2X1 NAND2X1_1325 ( .gnd(gnd), .vdd(vdd), .A(_8920_), .B(_10042_), .Y(_10043_) );
NOR2X1 NOR2X1_1611 ( .gnd(gnd), .vdd(vdd), .A(_10043_), .B(_9716_), .Y(_10044_) );
AOI21X1 AOI21X1_1786 ( .gnd(gnd), .vdd(vdd), .A(_9366_), .B(_9837_), .C(_10037_), .Y(_10045_) );
OAI21X1 OAI21X1_2825 ( .gnd(gnd), .vdd(vdd), .A(_10037_), .B(_9366_), .C(micro_hash_ucr_3_pipe10_bF_buf0), .Y(_10046_) );
AND2X2 AND2X2_685 ( .gnd(gnd), .vdd(vdd), .A(_10046_), .B(_9379_), .Y(_10047_) );
OAI21X1 OAI21X1_2826 ( .gnd(gnd), .vdd(vdd), .A(_10044_), .B(_10045_), .C(_10047_), .Y(_10048_) );
AOI21X1 AOI21X1_1787 ( .gnd(gnd), .vdd(vdd), .A(_10041_), .B(_10048_), .C(_10040_), .Y(_10049_) );
OAI21X1 OAI21X1_2827 ( .gnd(gnd), .vdd(vdd), .A(_9335__bF_buf1), .B(micro_hash_ucr_3_a_6_bF_buf3_), .C(_9337_), .Y(_10050_) );
OAI22X1 OAI22X1_125 ( .gnd(gnd), .vdd(vdd), .A(_9337_), .B(_10038_), .C(_10049_), .D(_10050_), .Y(_10051_) );
NAND2X1 NAND2X1_1326 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe16_bF_buf4), .B(_8923_), .Y(_10052_) );
OAI21X1 OAI21X1_2828 ( .gnd(gnd), .vdd(vdd), .A(_10051_), .B(micro_hash_ucr_3_pipe16_bF_buf3), .C(_10052_), .Y(_10053_) );
NAND2X1 NAND2X1_1327 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe17_bF_buf0), .B(_10037_), .Y(_10054_) );
OAI21X1 OAI21X1_2829 ( .gnd(gnd), .vdd(vdd), .A(_10053_), .B(micro_hash_ucr_3_pipe17_bF_buf3), .C(_10054_), .Y(_10055_) );
OAI21X1 OAI21X1_2830 ( .gnd(gnd), .vdd(vdd), .A(_8923_), .B(_9334__bF_buf0), .C(_9333__bF_buf2), .Y(_10056_) );
AOI21X1 AOI21X1_1788 ( .gnd(gnd), .vdd(vdd), .A(_9334__bF_buf3), .B(_10055_), .C(_10056_), .Y(_10057_) );
OAI21X1 OAI21X1_2831 ( .gnd(gnd), .vdd(vdd), .A(_10037_), .B(_9333__bF_buf1), .C(_9329__bF_buf0), .Y(_10058_) );
OAI22X1 OAI22X1_126 ( .gnd(gnd), .vdd(vdd), .A(_8923_), .B(_9329__bF_buf4), .C(_10057_), .D(_10058_), .Y(_10059_) );
OAI21X1 OAI21X1_2832 ( .gnd(gnd), .vdd(vdd), .A(_10038_), .B(_9331_), .C(_9330__bF_buf3), .Y(_10060_) );
AOI21X1 AOI21X1_1789 ( .gnd(gnd), .vdd(vdd), .A(_9331_), .B(_10059_), .C(_10060_), .Y(_10061_) );
OAI21X1 OAI21X1_2833 ( .gnd(gnd), .vdd(vdd), .A(_9330__bF_buf2), .B(micro_hash_ucr_3_a_6_bF_buf2_), .C(_9326__bF_buf3), .Y(_10062_) );
AOI21X1 AOI21X1_1790 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe23), .B(_10037_), .C(micro_hash_ucr_3_pipe24_bF_buf2), .Y(_10063_) );
OAI21X1 OAI21X1_2834 ( .gnd(gnd), .vdd(vdd), .A(_10061_), .B(_10062_), .C(_10063_), .Y(_10064_) );
NAND2X1 NAND2X1_1328 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe24_bF_buf1), .B(_8923_), .Y(_10065_) );
AOI21X1 AOI21X1_1791 ( .gnd(gnd), .vdd(vdd), .A(_10065_), .B(_10064_), .C(micro_hash_ucr_3_pipe25_bF_buf0), .Y(_10066_) );
NOR2X1 NOR2X1_1612 ( .gnd(gnd), .vdd(vdd), .A(_9327_), .B(_10037_), .Y(_10067_) );
OAI21X1 OAI21X1_2835 ( .gnd(gnd), .vdd(vdd), .A(_10066_), .B(_10067_), .C(_9323__bF_buf3), .Y(_10068_) );
NAND3X1 NAND3X1_525 ( .gnd(gnd), .vdd(vdd), .A(_9325__bF_buf1), .B(_10039_), .C(_10068_), .Y(_10069_) );
NAND2X1 NAND2X1_1329 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe27), .B(_10037_), .Y(_10070_) );
AOI21X1 AOI21X1_1792 ( .gnd(gnd), .vdd(vdd), .A(_10070_), .B(_10069_), .C(micro_hash_ucr_3_pipe28_bF_buf3), .Y(_10071_) );
OAI21X1 OAI21X1_2836 ( .gnd(gnd), .vdd(vdd), .A(_8923_), .B(_9324__bF_buf1), .C(_9320_), .Y(_10072_) );
AOI21X1 AOI21X1_1793 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe29_bF_buf3), .B(_10038_), .C(micro_hash_ucr_3_pipe30_bF_buf4), .Y(_10073_) );
OAI21X1 OAI21X1_2837 ( .gnd(gnd), .vdd(vdd), .A(_10071_), .B(_10072_), .C(_10073_), .Y(_10074_) );
NAND2X1 NAND2X1_1330 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_6_bF_buf1_), .B(micro_hash_ucr_3_pipe30_bF_buf3), .Y(_10075_) );
AOI21X1 AOI21X1_1794 ( .gnd(gnd), .vdd(vdd), .A(_10075_), .B(_10074_), .C(micro_hash_ucr_3_pipe31), .Y(_10076_) );
OAI21X1 OAI21X1_2838 ( .gnd(gnd), .vdd(vdd), .A(_10038_), .B(_9321__bF_buf0), .C(_9317__bF_buf1), .Y(_10077_) );
AOI21X1 AOI21X1_1795 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe32_bF_buf1), .B(_8923_), .C(micro_hash_ucr_3_pipe33_bF_buf0), .Y(_10078_) );
OAI21X1 OAI21X1_2839 ( .gnd(gnd), .vdd(vdd), .A(_10076_), .B(_10077_), .C(_10078_), .Y(_10079_) );
OAI21X1 OAI21X1_2840 ( .gnd(gnd), .vdd(vdd), .A(_9319_), .B(_10038_), .C(_10079_), .Y(_10080_) );
NAND2X1 NAND2X1_1331 ( .gnd(gnd), .vdd(vdd), .A(_9318__bF_buf3), .B(_10080_), .Y(_10081_) );
OAI21X1 OAI21X1_2841 ( .gnd(gnd), .vdd(vdd), .A(_8923_), .B(_9318__bF_buf2), .C(_10081_), .Y(_10082_) );
AOI21X1 AOI21X1_1796 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe35_bF_buf0), .B(_10038_), .C(micro_hash_ucr_3_pipe36_bF_buf0), .Y(_10083_) );
OAI21X1 OAI21X1_2842 ( .gnd(gnd), .vdd(vdd), .A(_10082_), .B(micro_hash_ucr_3_pipe35_bF_buf3), .C(_10083_), .Y(_10084_) );
NAND2X1 NAND2X1_1332 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_6_bF_buf0_), .B(micro_hash_ucr_3_pipe36_bF_buf4), .Y(_10085_) );
NAND3X1 NAND3X1_526 ( .gnd(gnd), .vdd(vdd), .A(_9315_), .B(_10085_), .C(_10084_), .Y(_10086_) );
OAI21X1 OAI21X1_2843 ( .gnd(gnd), .vdd(vdd), .A(_10036_), .B(_10035_), .C(micro_hash_ucr_3_pipe37_bF_buf0), .Y(_10087_) );
NAND3X1 NAND3X1_527 ( .gnd(gnd), .vdd(vdd), .A(_9311__bF_buf1), .B(_10087_), .C(_10086_), .Y(_10088_) );
NAND3X1 NAND3X1_528 ( .gnd(gnd), .vdd(vdd), .A(_9313_), .B(_10034_), .C(_10088_), .Y(_10089_) );
OAI21X1 OAI21X1_2844 ( .gnd(gnd), .vdd(vdd), .A(_10036_), .B(_10035_), .C(micro_hash_ucr_3_pipe39_bF_buf0), .Y(_10090_) );
NAND3X1 NAND3X1_529 ( .gnd(gnd), .vdd(vdd), .A(_9312__bF_buf3), .B(_10090_), .C(_10089_), .Y(_10091_) );
NAND3X1 NAND3X1_530 ( .gnd(gnd), .vdd(vdd), .A(_9308_), .B(_10033_), .C(_10091_), .Y(_10092_) );
OAI21X1 OAI21X1_2845 ( .gnd(gnd), .vdd(vdd), .A(_10036_), .B(_10035_), .C(micro_hash_ucr_3_pipe41_bF_buf1), .Y(_10093_) );
NAND3X1 NAND3X1_531 ( .gnd(gnd), .vdd(vdd), .A(_9310__bF_buf0), .B(_10093_), .C(_10092_), .Y(_10094_) );
NAND3X1 NAND3X1_532 ( .gnd(gnd), .vdd(vdd), .A(_9309__bF_buf0), .B(_10032_), .C(_10094_), .Y(_10095_) );
OAI21X1 OAI21X1_2846 ( .gnd(gnd), .vdd(vdd), .A(_10036_), .B(_10035_), .C(micro_hash_ucr_3_pipe43), .Y(_10096_) );
NAND3X1 NAND3X1_533 ( .gnd(gnd), .vdd(vdd), .A(_9305__bF_buf2), .B(_10096_), .C(_10095_), .Y(_10097_) );
NAND3X1 NAND3X1_534 ( .gnd(gnd), .vdd(vdd), .A(_9307_), .B(_10031_), .C(_10097_), .Y(_10098_) );
OAI21X1 OAI21X1_2847 ( .gnd(gnd), .vdd(vdd), .A(_10036_), .B(_10035_), .C(micro_hash_ucr_3_pipe45_bF_buf0), .Y(_10099_) );
NAND3X1 NAND3X1_535 ( .gnd(gnd), .vdd(vdd), .A(_9306__bF_buf3), .B(_10099_), .C(_10098_), .Y(_10100_) );
NAND3X1 NAND3X1_536 ( .gnd(gnd), .vdd(vdd), .A(_9302_), .B(_10030_), .C(_10100_), .Y(_10101_) );
OAI21X1 OAI21X1_2848 ( .gnd(gnd), .vdd(vdd), .A(_10036_), .B(_10035_), .C(micro_hash_ucr_3_pipe47), .Y(_10102_) );
NAND3X1 NAND3X1_537 ( .gnd(gnd), .vdd(vdd), .A(_9304__bF_buf0), .B(_10102_), .C(_10101_), .Y(_10103_) );
NAND3X1 NAND3X1_538 ( .gnd(gnd), .vdd(vdd), .A(_9303_), .B(_10029_), .C(_10103_), .Y(_10104_) );
OAI21X1 OAI21X1_2849 ( .gnd(gnd), .vdd(vdd), .A(_10036_), .B(_10035_), .C(micro_hash_ucr_3_pipe49_bF_buf0), .Y(_10105_) );
NAND3X1 NAND3X1_539 ( .gnd(gnd), .vdd(vdd), .A(_9299__bF_buf3), .B(_10105_), .C(_10104_), .Y(_10106_) );
NAND3X1 NAND3X1_540 ( .gnd(gnd), .vdd(vdd), .A(_9301__bF_buf3), .B(_10028_), .C(_10106_), .Y(_10107_) );
OAI21X1 OAI21X1_2850 ( .gnd(gnd), .vdd(vdd), .A(_10036_), .B(_10035_), .C(micro_hash_ucr_3_pipe51), .Y(_10108_) );
NAND3X1 NAND3X1_541 ( .gnd(gnd), .vdd(vdd), .A(_9300__bF_buf3), .B(_10108_), .C(_10107_), .Y(_10109_) );
NAND3X1 NAND3X1_542 ( .gnd(gnd), .vdd(vdd), .A(_9296_), .B(_10027_), .C(_10109_), .Y(_10110_) );
OAI21X1 OAI21X1_2851 ( .gnd(gnd), .vdd(vdd), .A(_10036_), .B(_10035_), .C(micro_hash_ucr_3_pipe53), .Y(_10111_) );
NAND3X1 NAND3X1_543 ( .gnd(gnd), .vdd(vdd), .A(_9298__bF_buf1), .B(_10111_), .C(_10110_), .Y(_10112_) );
AOI21X1 AOI21X1_1797 ( .gnd(gnd), .vdd(vdd), .A(_10026_), .B(_10112_), .C(micro_hash_ucr_3_pipe55), .Y(_10113_) );
OAI21X1 OAI21X1_2852 ( .gnd(gnd), .vdd(vdd), .A(_10038_), .B(_9297_), .C(_9293__bF_buf1), .Y(_10114_) );
AOI21X1 AOI21X1_1798 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe56_bF_buf1), .B(_8923_), .C(micro_hash_ucr_3_pipe57_bF_buf0), .Y(_10115_) );
OAI21X1 OAI21X1_2853 ( .gnd(gnd), .vdd(vdd), .A(_10113_), .B(_10114_), .C(_10115_), .Y(_10116_) );
AOI21X1 AOI21X1_1799 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe57_bF_buf3), .B(_10037_), .C(micro_hash_ucr_3_pipe58_bF_buf1), .Y(_10117_) );
AOI22X1 AOI22X1_71 ( .gnd(gnd), .vdd(vdd), .A(_8923_), .B(micro_hash_ucr_3_pipe58_bF_buf0), .C(_10116_), .D(_10117_), .Y(_10118_) );
OAI21X1 OAI21X1_2854 ( .gnd(gnd), .vdd(vdd), .A(_10036_), .B(_10035_), .C(micro_hash_ucr_3_pipe59), .Y(_10119_) );
OAI21X1 OAI21X1_2855 ( .gnd(gnd), .vdd(vdd), .A(_10118_), .B(micro_hash_ucr_3_pipe59), .C(_10119_), .Y(_10120_) );
AOI21X1 AOI21X1_1800 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_6_bF_buf3_), .B(micro_hash_ucr_3_pipe60_bF_buf2), .C(micro_hash_ucr_3_pipe61_bF_buf1), .Y(_10121_) );
OAI21X1 OAI21X1_2856 ( .gnd(gnd), .vdd(vdd), .A(_10120_), .B(micro_hash_ucr_3_pipe60_bF_buf1), .C(_10121_), .Y(_10122_) );
OAI21X1 OAI21X1_2857 ( .gnd(gnd), .vdd(vdd), .A(_10036_), .B(_10035_), .C(micro_hash_ucr_3_pipe61_bF_buf0), .Y(_10123_) );
AOI21X1 AOI21X1_1801 ( .gnd(gnd), .vdd(vdd), .A(_10123_), .B(_10122_), .C(micro_hash_ucr_3_pipe62_bF_buf1), .Y(_10124_) );
OAI21X1 OAI21X1_2858 ( .gnd(gnd), .vdd(vdd), .A(_9287__bF_buf1), .B(micro_hash_ucr_3_a_6_bF_buf2_), .C(_9289__bF_buf3), .Y(_10125_) );
AOI21X1 AOI21X1_1802 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe63), .B(_10037_), .C(micro_hash_ucr_3_pipe64_bF_buf3), .Y(_10126_) );
OAI21X1 OAI21X1_2859 ( .gnd(gnd), .vdd(vdd), .A(_10124_), .B(_10125_), .C(_10126_), .Y(_10127_) );
NAND2X1 NAND2X1_1333 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe64_bF_buf2), .B(_8923_), .Y(_10128_) );
NAND3X1 NAND3X1_544 ( .gnd(gnd), .vdd(vdd), .A(_9284_), .B(_10128_), .C(_10127_), .Y(_10129_) );
NAND2X1 NAND2X1_1334 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe65_bF_buf3), .B(_10037_), .Y(_10130_) );
AOI21X1 AOI21X1_1803 ( .gnd(gnd), .vdd(vdd), .A(_10130_), .B(_10129_), .C(micro_hash_ucr_3_pipe66_bF_buf1), .Y(_10131_) );
OAI21X1 OAI21X1_2860 ( .gnd(gnd), .vdd(vdd), .A(_8923_), .B(_9286__bF_buf1), .C(_9285__bF_buf1), .Y(_10132_) );
AOI21X1 AOI21X1_1804 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe67), .B(_10038_), .C(micro_hash_ucr_3_pipe68_bF_buf3), .Y(_10133_) );
OAI21X1 OAI21X1_2861 ( .gnd(gnd), .vdd(vdd), .A(_10131_), .B(_10132_), .C(_10133_), .Y(_10134_) );
AOI21X1 AOI21X1_1805 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_6_bF_buf1_), .B(micro_hash_ucr_3_pipe68_bF_buf2), .C(micro_hash_ucr_3_pipe69), .Y(_10135_) );
OAI21X1 OAI21X1_2862 ( .gnd(gnd), .vdd(vdd), .A(_10037_), .B(_9283__bF_buf3), .C(_8705__bF_buf10), .Y(_10136_) );
AOI21X1 AOI21X1_1806 ( .gnd(gnd), .vdd(vdd), .A(_10135_), .B(_10134_), .C(_10136_), .Y(_8700__6_) );
NAND2X1 NAND2X1_1335 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_7_bF_buf2_), .B(micro_hash_ucr_3_pipe60_bF_buf0), .Y(_10137_) );
NAND2X1 NAND2X1_1336 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_7_bF_buf1_), .B(micro_hash_ucr_3_pipe58_bF_buf3), .Y(_10138_) );
NAND2X1 NAND2X1_1337 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_7_bF_buf0_), .B(micro_hash_ucr_3_pipe56_bF_buf0), .Y(_10139_) );
NAND2X1 NAND2X1_1338 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_7_bF_buf3_), .B(micro_hash_ucr_3_pipe54_bF_buf0), .Y(_10140_) );
NAND2X1 NAND2X1_1339 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_7_bF_buf2_), .B(micro_hash_ucr_3_pipe52_bF_buf2), .Y(_10141_) );
NAND2X1 NAND2X1_1340 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_7_bF_buf1_), .B(micro_hash_ucr_3_pipe50_bF_buf3), .Y(_10142_) );
NAND2X1 NAND2X1_1341 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_7_bF_buf0_), .B(micro_hash_ucr_3_pipe48_bF_buf0), .Y(_10143_) );
INVX8 INVX8_274 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_7_bF_buf3_), .Y(_10144_) );
NAND2X1 NAND2X1_1342 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe42_bF_buf1), .B(_10144_), .Y(_10145_) );
NOR2X1 NOR2X1_1613 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_7_), .B(micro_hash_ucr_3_b_7_bF_buf2_), .Y(_10146_) );
NAND2X1 NAND2X1_1343 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_7_), .B(micro_hash_ucr_3_b_7_bF_buf1_), .Y(_10147_) );
INVX4 INVX4_151 ( .gnd(gnd), .vdd(vdd), .A(_10147_), .Y(_10148_) );
OR2X2 OR2X2_71 ( .gnd(gnd), .vdd(vdd), .A(_10148_), .B(_10146_), .Y(_10149_) );
INVX8 INVX8_275 ( .gnd(gnd), .vdd(vdd), .A(_10149_), .Y(_10150_) );
NAND2X1 NAND2X1_1344 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe17_bF_buf2), .B(_10150_), .Y(_10151_) );
NAND2X1 NAND2X1_1345 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe15_bF_buf1), .B(_10150_), .Y(_10152_) );
NOR2X1 NOR2X1_1614 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_7_bF_buf2_), .B(_9340_), .Y(_10153_) );
NAND2X1 NAND2X1_1346 ( .gnd(gnd), .vdd(vdd), .A(_10144_), .B(_9371_), .Y(_10154_) );
NOR2X1 NOR2X1_1615 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe10_bF_buf3), .B(_9372_), .Y(_10155_) );
NOR2X1 NOR2X1_1616 ( .gnd(gnd), .vdd(vdd), .A(H_3_7_), .B(micro_hash_ucr_3_pipe12), .Y(_10156_) );
NAND3X1 NAND3X1_545 ( .gnd(gnd), .vdd(vdd), .A(_9829_), .B(_10156_), .C(_10155_), .Y(_10157_) );
AOI21X1 AOI21X1_1807 ( .gnd(gnd), .vdd(vdd), .A(_10154_), .B(_10157_), .C(micro_hash_ucr_3_pipe11), .Y(_10158_) );
OAI21X1 OAI21X1_2863 ( .gnd(gnd), .vdd(vdd), .A(_10158_), .B(_10153_), .C(_9339_), .Y(_10159_) );
AOI21X1 AOI21X1_1808 ( .gnd(gnd), .vdd(vdd), .A(_10149_), .B(_9599_), .C(micro_hash_ucr_3_pipe14_bF_buf2), .Y(_10160_) );
AOI22X1 AOI22X1_72 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_7_bF_buf1_), .B(micro_hash_ucr_3_pipe14_bF_buf1), .C(_10159_), .D(_10160_), .Y(_10161_) );
OAI21X1 OAI21X1_2864 ( .gnd(gnd), .vdd(vdd), .A(_10161_), .B(micro_hash_ucr_3_pipe15_bF_buf0), .C(_10152_), .Y(_10162_) );
NAND2X1 NAND2X1_1347 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe16_bF_buf2), .B(_10144_), .Y(_10163_) );
OAI21X1 OAI21X1_2865 ( .gnd(gnd), .vdd(vdd), .A(_10162_), .B(micro_hash_ucr_3_pipe16_bF_buf1), .C(_10163_), .Y(_10164_) );
OAI21X1 OAI21X1_2866 ( .gnd(gnd), .vdd(vdd), .A(_10164_), .B(micro_hash_ucr_3_pipe17_bF_buf1), .C(_10151_), .Y(_10165_) );
OAI21X1 OAI21X1_2867 ( .gnd(gnd), .vdd(vdd), .A(_10144_), .B(_9334__bF_buf2), .C(_9333__bF_buf0), .Y(_10166_) );
AOI21X1 AOI21X1_1809 ( .gnd(gnd), .vdd(vdd), .A(_9334__bF_buf1), .B(_10165_), .C(_10166_), .Y(_10167_) );
OAI21X1 OAI21X1_2868 ( .gnd(gnd), .vdd(vdd), .A(_10150_), .B(_9333__bF_buf3), .C(_9329__bF_buf3), .Y(_10168_) );
OAI22X1 OAI22X1_127 ( .gnd(gnd), .vdd(vdd), .A(_10144_), .B(_9329__bF_buf2), .C(_10167_), .D(_10168_), .Y(_10169_) );
OAI21X1 OAI21X1_2869 ( .gnd(gnd), .vdd(vdd), .A(_10148_), .B(_10146_), .C(micro_hash_ucr_3_pipe21_bF_buf3), .Y(_10170_) );
OAI21X1 OAI21X1_2870 ( .gnd(gnd), .vdd(vdd), .A(_10169_), .B(micro_hash_ucr_3_pipe21_bF_buf2), .C(_10170_), .Y(_10171_) );
AOI21X1 AOI21X1_1810 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_7_bF_buf0_), .B(micro_hash_ucr_3_pipe22_bF_buf0), .C(micro_hash_ucr_3_pipe23), .Y(_10172_) );
OAI21X1 OAI21X1_2871 ( .gnd(gnd), .vdd(vdd), .A(_10171_), .B(micro_hash_ucr_3_pipe22_bF_buf4), .C(_10172_), .Y(_10173_) );
OAI21X1 OAI21X1_2872 ( .gnd(gnd), .vdd(vdd), .A(_9326__bF_buf2), .B(_10150_), .C(_10173_), .Y(_10174_) );
NAND2X1 NAND2X1_1348 ( .gnd(gnd), .vdd(vdd), .A(_9328__bF_buf3), .B(_10174_), .Y(_10175_) );
OAI21X1 OAI21X1_2873 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_7_bF_buf3_), .B(_9328__bF_buf2), .C(_10175_), .Y(_10176_) );
NAND2X1 NAND2X1_1349 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe25_bF_buf3), .B(_10150_), .Y(_10177_) );
OAI21X1 OAI21X1_2874 ( .gnd(gnd), .vdd(vdd), .A(_10176_), .B(micro_hash_ucr_3_pipe25_bF_buf2), .C(_10177_), .Y(_10178_) );
NAND2X1 NAND2X1_1350 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe26_bF_buf1), .B(_10144_), .Y(_10179_) );
OAI21X1 OAI21X1_2875 ( .gnd(gnd), .vdd(vdd), .A(_10178_), .B(micro_hash_ucr_3_pipe26_bF_buf0), .C(_10179_), .Y(_10180_) );
NAND2X1 NAND2X1_1351 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe27), .B(_10150_), .Y(_10181_) );
OAI21X1 OAI21X1_2876 ( .gnd(gnd), .vdd(vdd), .A(_10180_), .B(micro_hash_ucr_3_pipe27), .C(_10181_), .Y(_10182_) );
OAI21X1 OAI21X1_2877 ( .gnd(gnd), .vdd(vdd), .A(_10144_), .B(_9324__bF_buf0), .C(_9320_), .Y(_10183_) );
AOI21X1 AOI21X1_1811 ( .gnd(gnd), .vdd(vdd), .A(_9324__bF_buf4), .B(_10182_), .C(_10183_), .Y(_10184_) );
NOR2X1 NOR2X1_1617 ( .gnd(gnd), .vdd(vdd), .A(_9320_), .B(_10150_), .Y(_10185_) );
OAI21X1 OAI21X1_2878 ( .gnd(gnd), .vdd(vdd), .A(_10184_), .B(_10185_), .C(_9322__bF_buf3), .Y(_10186_) );
AOI21X1 AOI21X1_1812 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe30_bF_buf2), .B(_10144_), .C(micro_hash_ucr_3_pipe31), .Y(_10187_) );
OAI21X1 OAI21X1_2879 ( .gnd(gnd), .vdd(vdd), .A(_10149_), .B(_9321__bF_buf3), .C(_9317__bF_buf0), .Y(_10188_) );
AOI21X1 AOI21X1_1813 ( .gnd(gnd), .vdd(vdd), .A(_10187_), .B(_10186_), .C(_10188_), .Y(_10189_) );
NOR2X1 NOR2X1_1618 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_7_bF_buf2_), .B(_9317__bF_buf4), .Y(_10190_) );
NOR3X1 NOR3X1_8 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe33_bF_buf3), .B(_10190_), .C(_10189_), .Y(_10191_) );
OAI21X1 OAI21X1_2880 ( .gnd(gnd), .vdd(vdd), .A(_10149_), .B(_9319_), .C(_9318__bF_buf1), .Y(_10192_) );
AOI21X1 AOI21X1_1814 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe34_bF_buf1), .B(_10144_), .C(micro_hash_ucr_3_pipe35_bF_buf2), .Y(_10193_) );
OAI21X1 OAI21X1_2881 ( .gnd(gnd), .vdd(vdd), .A(_10191_), .B(_10192_), .C(_10193_), .Y(_10194_) );
AOI21X1 AOI21X1_1815 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe35_bF_buf1), .B(_10150_), .C(micro_hash_ucr_3_pipe36_bF_buf3), .Y(_10195_) );
AOI22X1 AOI22X1_73 ( .gnd(gnd), .vdd(vdd), .A(_10144_), .B(micro_hash_ucr_3_pipe36_bF_buf2), .C(_10194_), .D(_10195_), .Y(_10196_) );
OAI21X1 OAI21X1_2882 ( .gnd(gnd), .vdd(vdd), .A(_10149_), .B(_9315_), .C(_9311__bF_buf0), .Y(_10197_) );
AOI21X1 AOI21X1_1816 ( .gnd(gnd), .vdd(vdd), .A(_9315_), .B(_10196_), .C(_10197_), .Y(_10198_) );
OAI21X1 OAI21X1_2883 ( .gnd(gnd), .vdd(vdd), .A(_9311__bF_buf4), .B(micro_hash_ucr_3_a_7_bF_buf1_), .C(_9313_), .Y(_10199_) );
AOI21X1 AOI21X1_1817 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe39_bF_buf3), .B(_10150_), .C(micro_hash_ucr_3_pipe40_bF_buf3), .Y(_10200_) );
OAI21X1 OAI21X1_2884 ( .gnd(gnd), .vdd(vdd), .A(_10198_), .B(_10199_), .C(_10200_), .Y(_10201_) );
NAND2X1 NAND2X1_1352 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe40_bF_buf2), .B(_10144_), .Y(_10202_) );
NAND3X1 NAND3X1_546 ( .gnd(gnd), .vdd(vdd), .A(_9308_), .B(_10202_), .C(_10201_), .Y(_10203_) );
NAND2X1 NAND2X1_1353 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe41_bF_buf0), .B(_10150_), .Y(_10204_) );
NAND3X1 NAND3X1_547 ( .gnd(gnd), .vdd(vdd), .A(_9310__bF_buf4), .B(_10204_), .C(_10203_), .Y(_10205_) );
NAND3X1 NAND3X1_548 ( .gnd(gnd), .vdd(vdd), .A(_9309__bF_buf3), .B(_10145_), .C(_10205_), .Y(_10206_) );
NAND2X1 NAND2X1_1354 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe43), .B(_10150_), .Y(_10207_) );
AOI21X1 AOI21X1_1818 ( .gnd(gnd), .vdd(vdd), .A(_10207_), .B(_10206_), .C(micro_hash_ucr_3_pipe44_bF_buf3), .Y(_10208_) );
OAI21X1 OAI21X1_2885 ( .gnd(gnd), .vdd(vdd), .A(_10144_), .B(_9305__bF_buf1), .C(_9307_), .Y(_10209_) );
AOI21X1 AOI21X1_1819 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe45_bF_buf3), .B(_10149_), .C(micro_hash_ucr_3_pipe46_bF_buf2), .Y(_10210_) );
OAI21X1 OAI21X1_2886 ( .gnd(gnd), .vdd(vdd), .A(_10208_), .B(_10209_), .C(_10210_), .Y(_10211_) );
NAND2X1 NAND2X1_1355 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_7_bF_buf0_), .B(micro_hash_ucr_3_pipe46_bF_buf1), .Y(_10212_) );
NAND3X1 NAND3X1_549 ( .gnd(gnd), .vdd(vdd), .A(_9302_), .B(_10212_), .C(_10211_), .Y(_10213_) );
OAI21X1 OAI21X1_2887 ( .gnd(gnd), .vdd(vdd), .A(_10148_), .B(_10146_), .C(micro_hash_ucr_3_pipe47), .Y(_10214_) );
NAND3X1 NAND3X1_550 ( .gnd(gnd), .vdd(vdd), .A(_9304__bF_buf3), .B(_10214_), .C(_10213_), .Y(_10215_) );
NAND3X1 NAND3X1_551 ( .gnd(gnd), .vdd(vdd), .A(_9303_), .B(_10143_), .C(_10215_), .Y(_10216_) );
OAI21X1 OAI21X1_2888 ( .gnd(gnd), .vdd(vdd), .A(_10148_), .B(_10146_), .C(micro_hash_ucr_3_pipe49_bF_buf3), .Y(_10217_) );
NAND3X1 NAND3X1_552 ( .gnd(gnd), .vdd(vdd), .A(_9299__bF_buf2), .B(_10217_), .C(_10216_), .Y(_10218_) );
NAND3X1 NAND3X1_553 ( .gnd(gnd), .vdd(vdd), .A(_9301__bF_buf2), .B(_10142_), .C(_10218_), .Y(_10219_) );
OAI21X1 OAI21X1_2889 ( .gnd(gnd), .vdd(vdd), .A(_10148_), .B(_10146_), .C(micro_hash_ucr_3_pipe51), .Y(_10220_) );
NAND3X1 NAND3X1_554 ( .gnd(gnd), .vdd(vdd), .A(_9300__bF_buf2), .B(_10220_), .C(_10219_), .Y(_10221_) );
NAND3X1 NAND3X1_555 ( .gnd(gnd), .vdd(vdd), .A(_9296_), .B(_10141_), .C(_10221_), .Y(_10222_) );
OAI21X1 OAI21X1_2890 ( .gnd(gnd), .vdd(vdd), .A(_10148_), .B(_10146_), .C(micro_hash_ucr_3_pipe53), .Y(_10223_) );
NAND3X1 NAND3X1_556 ( .gnd(gnd), .vdd(vdd), .A(_9298__bF_buf0), .B(_10223_), .C(_10222_), .Y(_10224_) );
NAND3X1 NAND3X1_557 ( .gnd(gnd), .vdd(vdd), .A(_9297_), .B(_10140_), .C(_10224_), .Y(_10225_) );
OAI21X1 OAI21X1_2891 ( .gnd(gnd), .vdd(vdd), .A(_10148_), .B(_10146_), .C(micro_hash_ucr_3_pipe55), .Y(_10226_) );
NAND3X1 NAND3X1_558 ( .gnd(gnd), .vdd(vdd), .A(_9293__bF_buf0), .B(_10226_), .C(_10225_), .Y(_10227_) );
NAND3X1 NAND3X1_559 ( .gnd(gnd), .vdd(vdd), .A(_9295_), .B(_10139_), .C(_10227_), .Y(_10228_) );
OAI21X1 OAI21X1_2892 ( .gnd(gnd), .vdd(vdd), .A(_10148_), .B(_10146_), .C(micro_hash_ucr_3_pipe57_bF_buf2), .Y(_10229_) );
NAND3X1 NAND3X1_560 ( .gnd(gnd), .vdd(vdd), .A(_9294__bF_buf1), .B(_10229_), .C(_10228_), .Y(_10230_) );
NAND3X1 NAND3X1_561 ( .gnd(gnd), .vdd(vdd), .A(_9290__bF_buf3), .B(_10138_), .C(_10230_), .Y(_10231_) );
OAI21X1 OAI21X1_2893 ( .gnd(gnd), .vdd(vdd), .A(_10148_), .B(_10146_), .C(micro_hash_ucr_3_pipe59), .Y(_10232_) );
NAND3X1 NAND3X1_562 ( .gnd(gnd), .vdd(vdd), .A(_9292__bF_buf0), .B(_10232_), .C(_10231_), .Y(_10233_) );
AOI21X1 AOI21X1_1820 ( .gnd(gnd), .vdd(vdd), .A(_10137_), .B(_10233_), .C(micro_hash_ucr_3_pipe61_bF_buf3), .Y(_10234_) );
OAI21X1 OAI21X1_2894 ( .gnd(gnd), .vdd(vdd), .A(_10149_), .B(_9291_), .C(_9287__bF_buf0), .Y(_10235_) );
AOI21X1 AOI21X1_1821 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe62_bF_buf0), .B(_10144_), .C(micro_hash_ucr_3_pipe63), .Y(_10236_) );
OAI21X1 OAI21X1_2895 ( .gnd(gnd), .vdd(vdd), .A(_10234_), .B(_10235_), .C(_10236_), .Y(_10237_) );
AOI21X1 AOI21X1_1822 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe63), .B(_10150_), .C(micro_hash_ucr_3_pipe64_bF_buf1), .Y(_10238_) );
NAND2X1 NAND2X1_1356 ( .gnd(gnd), .vdd(vdd), .A(_10238_), .B(_10237_), .Y(_10239_) );
NAND2X1 NAND2X1_1357 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe64_bF_buf0), .B(_10144_), .Y(_10240_) );
NAND3X1 NAND3X1_563 ( .gnd(gnd), .vdd(vdd), .A(_9284_), .B(_10240_), .C(_10239_), .Y(_10241_) );
NAND2X1 NAND2X1_1358 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe65_bF_buf2), .B(_10150_), .Y(_10242_) );
AOI21X1 AOI21X1_1823 ( .gnd(gnd), .vdd(vdd), .A(_10242_), .B(_10241_), .C(micro_hash_ucr_3_pipe66_bF_buf0), .Y(_10243_) );
OAI21X1 OAI21X1_2896 ( .gnd(gnd), .vdd(vdd), .A(_10144_), .B(_9286__bF_buf0), .C(_9285__bF_buf0), .Y(_10244_) );
AOI21X1 AOI21X1_1824 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe67), .B(_10149_), .C(micro_hash_ucr_3_pipe68_bF_buf1), .Y(_10245_) );
OAI21X1 OAI21X1_2897 ( .gnd(gnd), .vdd(vdd), .A(_10243_), .B(_10244_), .C(_10245_), .Y(_10246_) );
AOI21X1 AOI21X1_1825 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_a_7_bF_buf3_), .B(micro_hash_ucr_3_pipe68_bF_buf0), .C(micro_hash_ucr_3_pipe69), .Y(_10247_) );
OAI21X1 OAI21X1_2898 ( .gnd(gnd), .vdd(vdd), .A(_10150_), .B(_9283__bF_buf2), .C(_8705__bF_buf9), .Y(_10248_) );
AOI21X1 AOI21X1_1826 ( .gnd(gnd), .vdd(vdd), .A(_10247_), .B(_10246_), .C(_10248_), .Y(_8700__7_) );
INVX1 INVX1_628 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_k_0_), .Y(_10249_) );
NOR2X1 NOR2X1_1619 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe40_bF_buf1), .B(micro_hash_ucr_3_pipe7), .Y(_10250_) );
AOI21X1 AOI21X1_1827 ( .gnd(gnd), .vdd(vdd), .A(_10249_), .B(_10250_), .C(_8800__bF_buf3), .Y(_8704__0_) );
NAND2X1 NAND2X1_1359 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_k_1_), .B(_10250_), .Y(_10251_) );
NOR2X1 NOR2X1_1620 ( .gnd(gnd), .vdd(vdd), .A(_10251_), .B(_8800__bF_buf2), .Y(_8704__1_) );
NAND2X1 NAND2X1_1360 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_k_2_), .B(_10250_), .Y(_10252_) );
NOR2X1 NOR2X1_1621 ( .gnd(gnd), .vdd(vdd), .A(_10252_), .B(_8800__bF_buf1), .Y(_8704__2_) );
OAI21X1 OAI21X1_2899 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe7), .B(micro_hash_ucr_3_k_3_), .C(_9312__bF_buf2), .Y(_10253_) );
NOR2X1 NOR2X1_1622 ( .gnd(gnd), .vdd(vdd), .A(_10253_), .B(_8800__bF_buf0), .Y(_8704__3_) );
OAI21X1 OAI21X1_2900 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe7), .B(micro_hash_ucr_3_k_4_), .C(_9312__bF_buf1), .Y(_10254_) );
NOR2X1 NOR2X1_1623 ( .gnd(gnd), .vdd(vdd), .A(_10254_), .B(_8800__bF_buf12), .Y(_8704__4_) );
INVX2 INVX2_358 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_k_5_), .Y(_10255_) );
OAI21X1 OAI21X1_2901 ( .gnd(gnd), .vdd(vdd), .A(_10255_), .B(micro_hash_ucr_3_pipe7), .C(_9312__bF_buf0), .Y(_10256_) );
AND2X2 AND2X2_686 ( .gnd(gnd), .vdd(vdd), .A(_8705__bF_buf8), .B(_10256_), .Y(_8704__5_) );
NAND2X1 NAND2X1_1361 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_k_6_), .B(_10250_), .Y(_10257_) );
NOR2X1 NOR2X1_1624 ( .gnd(gnd), .vdd(vdd), .A(_10257_), .B(_8800__bF_buf11), .Y(_8704__6_) );
INVX1 INVX1_629 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_k_7_), .Y(_10258_) );
AOI21X1 AOI21X1_1828 ( .gnd(gnd), .vdd(vdd), .A(_10258_), .B(_10250_), .C(_8800__bF_buf10), .Y(_8704__7_) );
NAND2X1 NAND2X1_1362 ( .gnd(gnd), .vdd(vdd), .A(_12902_), .B(_8862__bF_buf2), .Y(_10259_) );
NOR2X1 NOR2X1_1625 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe39_bF_buf2), .B(micro_hash_ucr_3_pipe37_bF_buf3), .Y(_10260_) );
NAND3X1 NAND3X1_564 ( .gnd(gnd), .vdd(vdd), .A(_9314_), .B(_9319_), .C(_10260_), .Y(_10261_) );
NOR2X1 NOR2X1_1626 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe31), .B(_10261_), .Y(_10262_) );
INVX1 INVX1_630 ( .gnd(gnd), .vdd(vdd), .A(_10262_), .Y(_10263_) );
NOR2X1 NOR2X1_1627 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe29_bF_buf2), .B(_10263_), .Y(_10264_) );
NOR2X1 NOR2X1_1628 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe23), .B(micro_hash_ucr_3_pipe21_bF_buf1), .Y(_10265_) );
INVX1 INVX1_631 ( .gnd(gnd), .vdd(vdd), .A(_10265_), .Y(_10266_) );
NOR2X1 NOR2X1_1629 ( .gnd(gnd), .vdd(vdd), .A(_9372_), .B(_10266_), .Y(_10267_) );
NAND3X1 NAND3X1_565 ( .gnd(gnd), .vdd(vdd), .A(_9332_), .B(_9333__bF_buf2), .C(_9366_), .Y(_10268_) );
NOR2X1 NOR2X1_1630 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe27), .B(micro_hash_ucr_3_pipe25_bF_buf1), .Y(_10269_) );
NAND2X1 NAND2X1_1363 ( .gnd(gnd), .vdd(vdd), .A(_9337_), .B(_10269_), .Y(_10270_) );
NOR2X1 NOR2X1_1631 ( .gnd(gnd), .vdd(vdd), .A(_10270_), .B(_10268_), .Y(_10271_) );
AND2X2 AND2X2_687 ( .gnd(gnd), .vdd(vdd), .A(_10271_), .B(_10267_), .Y(_10272_) );
NAND2X1 NAND2X1_1364 ( .gnd(gnd), .vdd(vdd), .A(_10272_), .B(_10264_), .Y(_10273_) );
INVX2 INVX2_359 ( .gnd(gnd), .vdd(vdd), .A(_10273_), .Y(_10274_) );
AOI21X1 AOI21X1_1829 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_0_bF_buf0_), .B(micro_hash_ucr_3_a_0_bF_buf3_), .C(_10274_), .Y(_10275_) );
NOR2X1 NOR2X1_1632 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe47), .B(micro_hash_ucr_3_pipe45_bF_buf2), .Y(_10276_) );
NOR2X1 NOR2X1_1633 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe41_bF_buf3), .B(micro_hash_ucr_3_pipe43), .Y(_10277_) );
NAND2X1 NAND2X1_1365 ( .gnd(gnd), .vdd(vdd), .A(_10276_), .B(_10277_), .Y(_10278_) );
INVX2 INVX2_360 ( .gnd(gnd), .vdd(vdd), .A(_10278_), .Y(_10279_) );
NOR2X1 NOR2X1_1634 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe51), .B(micro_hash_ucr_3_pipe49_bF_buf2), .Y(_10280_) );
INVX1 INVX1_632 ( .gnd(gnd), .vdd(vdd), .A(_10280_), .Y(_10281_) );
NOR2X1 NOR2X1_1635 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe59), .B(micro_hash_ucr_3_pipe57_bF_buf1), .Y(_10282_) );
INVX1 INVX1_633 ( .gnd(gnd), .vdd(vdd), .A(_10282_), .Y(_10283_) );
NOR2X1 NOR2X1_1636 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe65_bF_buf1), .B(micro_hash_ucr_3_pipe67), .Y(_10284_) );
NAND3X1 NAND3X1_566 ( .gnd(gnd), .vdd(vdd), .A(_9289__bF_buf2), .B(_9291_), .C(_10284_), .Y(_10285_) );
NOR2X1 NOR2X1_1637 ( .gnd(gnd), .vdd(vdd), .A(_10283_), .B(_10285_), .Y(_10286_) );
NOR2X1 NOR2X1_1638 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe53), .B(micro_hash_ucr_3_pipe55), .Y(_10287_) );
NAND2X1 NAND2X1_1366 ( .gnd(gnd), .vdd(vdd), .A(_10287_), .B(_10286_), .Y(_10288_) );
NOR2X1 NOR2X1_1639 ( .gnd(gnd), .vdd(vdd), .A(_10281_), .B(_10288_), .Y(_10289_) );
NAND2X1 NAND2X1_1367 ( .gnd(gnd), .vdd(vdd), .A(_10279_), .B(_10289_), .Y(_10290_) );
OAI21X1 OAI21X1_2902 ( .gnd(gnd), .vdd(vdd), .A(_10275_), .B(_10290_), .C(_10259_), .Y(_10291_) );
INVX2 INVX2_361 ( .gnd(gnd), .vdd(vdd), .A(_10290_), .Y(_10292_) );
INVX1 INVX1_634 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_x_0_), .Y(_10293_) );
NOR2X1 NOR2X1_1640 ( .gnd(gnd), .vdd(vdd), .A(_10293_), .B(_10273_), .Y(_10294_) );
AOI21X1 AOI21X1_1830 ( .gnd(gnd), .vdd(vdd), .A(_10292_), .B(_10294_), .C(micro_hash_ucr_3_pipe69), .Y(_10295_) );
OAI21X1 OAI21X1_2903 ( .gnd(gnd), .vdd(vdd), .A(_9283__bF_buf1), .B(_10259_), .C(_8705__bF_buf7), .Y(_10296_) );
AOI21X1 AOI21X1_1831 ( .gnd(gnd), .vdd(vdd), .A(_10295_), .B(_10291_), .C(_10296_), .Y(_8778__0_) );
NAND2X1 NAND2X1_1368 ( .gnd(gnd), .vdd(vdd), .A(_12908__bF_buf1), .B(_8868__bF_buf3), .Y(_10297_) );
OAI21X1 OAI21X1_2904 ( .gnd(gnd), .vdd(vdd), .A(_12908__bF_buf0), .B(_8868__bF_buf2), .C(_10273_), .Y(_10298_) );
NAND2X1 NAND2X1_1369 ( .gnd(gnd), .vdd(vdd), .A(_10292_), .B(_10298_), .Y(_10299_) );
NAND2X1 NAND2X1_1370 ( .gnd(gnd), .vdd(vdd), .A(_10269_), .B(_10265_), .Y(_10300_) );
NOR2X1 NOR2X1_1641 ( .gnd(gnd), .vdd(vdd), .A(_10300_), .B(_10278_), .Y(_10301_) );
NAND2X1 NAND2X1_1371 ( .gnd(gnd), .vdd(vdd), .A(_10280_), .B(_10287_), .Y(_10302_) );
NOR2X1 NOR2X1_1642 ( .gnd(gnd), .vdd(vdd), .A(_10302_), .B(_10261_), .Y(_10303_) );
NAND2X1 NAND2X1_1372 ( .gnd(gnd), .vdd(vdd), .A(_10301_), .B(_10303_), .Y(_10304_) );
NOR2X1 NOR2X1_1643 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe15_bF_buf3), .B(_9372_), .Y(_10305_) );
AND2X2 AND2X2_688 ( .gnd(gnd), .vdd(vdd), .A(_10305_), .B(_9332_), .Y(_10306_) );
NOR2X1 NOR2X1_1644 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe29_bF_buf1), .B(micro_hash_ucr_3_pipe31), .Y(_10307_) );
INVX1 INVX1_635 ( .gnd(gnd), .vdd(vdd), .A(_10307_), .Y(_10308_) );
NAND3X1 NAND3X1_567 ( .gnd(gnd), .vdd(vdd), .A(_9333__bF_buf1), .B(micro_hash_ucr_3_x_1_), .C(_9366_), .Y(_10309_) );
NOR2X1 NOR2X1_1645 ( .gnd(gnd), .vdd(vdd), .A(_10308_), .B(_10309_), .Y(_10310_) );
NAND3X1 NAND3X1_568 ( .gnd(gnd), .vdd(vdd), .A(_10286_), .B(_10310_), .C(_10306_), .Y(_10311_) );
OAI21X1 OAI21X1_2905 ( .gnd(gnd), .vdd(vdd), .A(_10311_), .B(_10304_), .C(_9283__bF_buf0), .Y(_10312_) );
AOI21X1 AOI21X1_1832 ( .gnd(gnd), .vdd(vdd), .A(_10297_), .B(_10299_), .C(_10312_), .Y(_10313_) );
OAI21X1 OAI21X1_2906 ( .gnd(gnd), .vdd(vdd), .A(_9283__bF_buf3), .B(_10297_), .C(_8705__bF_buf6), .Y(_10314_) );
NOR2X1 NOR2X1_1646 ( .gnd(gnd), .vdd(vdd), .A(_10314_), .B(_10313_), .Y(_8778__1_) );
NAND2X1 NAND2X1_1373 ( .gnd(gnd), .vdd(vdd), .A(_8789__bF_buf1), .B(_8884_), .Y(_10315_) );
OAI21X1 OAI21X1_2907 ( .gnd(gnd), .vdd(vdd), .A(_8789__bF_buf0), .B(_8884_), .C(_10273_), .Y(_10316_) );
NAND2X1 NAND2X1_1374 ( .gnd(gnd), .vdd(vdd), .A(_10292_), .B(_10316_), .Y(_10317_) );
INVX1 INVX1_636 ( .gnd(gnd), .vdd(vdd), .A(_10272_), .Y(_10318_) );
NAND2X1 NAND2X1_1375 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_x_2_), .B(_10279_), .Y(_10319_) );
NOR2X1 NOR2X1_1647 ( .gnd(gnd), .vdd(vdd), .A(_10302_), .B(_10319_), .Y(_10320_) );
NAND3X1 NAND3X1_569 ( .gnd(gnd), .vdd(vdd), .A(_10286_), .B(_10320_), .C(_10264_), .Y(_10321_) );
OAI21X1 OAI21X1_2908 ( .gnd(gnd), .vdd(vdd), .A(_10321_), .B(_10318_), .C(_9283__bF_buf2), .Y(_10322_) );
AOI21X1 AOI21X1_1833 ( .gnd(gnd), .vdd(vdd), .A(_10315_), .B(_10317_), .C(_10322_), .Y(_10323_) );
OAI21X1 OAI21X1_2909 ( .gnd(gnd), .vdd(vdd), .A(_9283__bF_buf1), .B(_10315_), .C(_8705__bF_buf5), .Y(_10324_) );
NOR2X1 NOR2X1_1648 ( .gnd(gnd), .vdd(vdd), .A(_10324_), .B(_10323_), .Y(_8778__2_) );
NAND2X1 NAND2X1_1376 ( .gnd(gnd), .vdd(vdd), .A(_8794_), .B(_9706__bF_buf2), .Y(_10325_) );
AOI21X1 AOI21X1_1834 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_3_bF_buf0_), .B(micro_hash_ucr_3_a_3_), .C(_10274_), .Y(_10326_) );
OAI21X1 OAI21X1_2910 ( .gnd(gnd), .vdd(vdd), .A(_10326_), .B(_10290_), .C(_10325_), .Y(_10327_) );
NAND3X1 NAND3X1_570 ( .gnd(gnd), .vdd(vdd), .A(_9320_), .B(micro_hash_ucr_3_x_3_), .C(_10279_), .Y(_10328_) );
NOR2X1 NOR2X1_1649 ( .gnd(gnd), .vdd(vdd), .A(_10328_), .B(_10263_), .Y(_10329_) );
AND2X2 AND2X2_689 ( .gnd(gnd), .vdd(vdd), .A(_10329_), .B(_10272_), .Y(_10330_) );
AOI21X1 AOI21X1_1835 ( .gnd(gnd), .vdd(vdd), .A(_10289_), .B(_10330_), .C(micro_hash_ucr_3_pipe69), .Y(_10331_) );
OAI21X1 OAI21X1_2911 ( .gnd(gnd), .vdd(vdd), .A(_9283__bF_buf0), .B(_10325_), .C(_8705__bF_buf4), .Y(_10332_) );
AOI21X1 AOI21X1_1836 ( .gnd(gnd), .vdd(vdd), .A(_10331_), .B(_10327_), .C(_10332_), .Y(_8778__3_) );
INVX4 INVX4_152 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_4_bF_buf0_), .Y(_10333_) );
NAND2X1 NAND2X1_1377 ( .gnd(gnd), .vdd(vdd), .A(_10333_), .B(_8903__bF_buf3), .Y(_10334_) );
OAI21X1 OAI21X1_2912 ( .gnd(gnd), .vdd(vdd), .A(_10333_), .B(_8903__bF_buf2), .C(_10273_), .Y(_10335_) );
NAND2X1 NAND2X1_1378 ( .gnd(gnd), .vdd(vdd), .A(_10292_), .B(_10335_), .Y(_10336_) );
NOR2X1 NOR2X1_1650 ( .gnd(gnd), .vdd(vdd), .A(_10268_), .B(_10261_), .Y(_10337_) );
NOR2X1 NOR2X1_1651 ( .gnd(gnd), .vdd(vdd), .A(_10308_), .B(_10266_), .Y(_10338_) );
NAND2X1 NAND2X1_1379 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_x_4_), .B(_9373_), .Y(_10339_) );
NOR2X1 NOR2X1_1652 ( .gnd(gnd), .vdd(vdd), .A(_10270_), .B(_10339_), .Y(_10340_) );
NAND3X1 NAND3X1_571 ( .gnd(gnd), .vdd(vdd), .A(_10337_), .B(_10338_), .C(_10340_), .Y(_10341_) );
OAI21X1 OAI21X1_2913 ( .gnd(gnd), .vdd(vdd), .A(_10290_), .B(_10341_), .C(_9283__bF_buf3), .Y(_10342_) );
AOI21X1 AOI21X1_1837 ( .gnd(gnd), .vdd(vdd), .A(_10334_), .B(_10336_), .C(_10342_), .Y(_10343_) );
OAI21X1 OAI21X1_2914 ( .gnd(gnd), .vdd(vdd), .A(_9283__bF_buf2), .B(_10334_), .C(_8705__bF_buf3), .Y(_10344_) );
NOR2X1 NOR2X1_1653 ( .gnd(gnd), .vdd(vdd), .A(_10344_), .B(_10343_), .Y(_8778__4_) );
INVX1 INVX1_637 ( .gnd(gnd), .vdd(vdd), .A(_10260_), .Y(_10345_) );
NAND2X1 NAND2X1_1380 ( .gnd(gnd), .vdd(vdd), .A(_9319_), .B(_9321__bF_buf2), .Y(_10346_) );
NOR2X1 NOR2X1_1654 ( .gnd(gnd), .vdd(vdd), .A(_10346_), .B(_10345_), .Y(_10347_) );
NOR2X1 NOR2X1_1655 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe19), .B(micro_hash_ucr_3_x_5_), .Y(_10348_) );
AND2X2 AND2X2_690 ( .gnd(gnd), .vdd(vdd), .A(_9366_), .B(_10348_), .Y(_10349_) );
NAND3X1 NAND3X1_572 ( .gnd(gnd), .vdd(vdd), .A(_10347_), .B(_10349_), .C(_10306_), .Y(_10350_) );
NOR2X1 NOR2X1_1656 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_5_bF_buf0_), .B(micro_hash_ucr_3_a_5_bF_buf1_), .Y(_10351_) );
NOR2X1 NOR2X1_1657 ( .gnd(gnd), .vdd(vdd), .A(_8814__bF_buf1), .B(_8909_), .Y(_10352_) );
NOR2X1 NOR2X1_1658 ( .gnd(gnd), .vdd(vdd), .A(_10351_), .B(_10352_), .Y(_10353_) );
NAND3X1 NAND3X1_573 ( .gnd(gnd), .vdd(vdd), .A(_9283__bF_buf1), .B(_10280_), .C(_10279_), .Y(_10354_) );
NOR2X1 NOR2X1_1659 ( .gnd(gnd), .vdd(vdd), .A(_10354_), .B(_10288_), .Y(_10355_) );
INVX2 INVX2_362 ( .gnd(gnd), .vdd(vdd), .A(_10355_), .Y(_10356_) );
NOR2X1 NOR2X1_1660 ( .gnd(gnd), .vdd(vdd), .A(_10273_), .B(_10356_), .Y(_10357_) );
OAI21X1 OAI21X1_2915 ( .gnd(gnd), .vdd(vdd), .A(_10357_), .B(_10353_), .C(_10350_), .Y(_10358_) );
NAND2X1 NAND2X1_1381 ( .gnd(gnd), .vdd(vdd), .A(_9314_), .B(_9320_), .Y(_10359_) );
NOR2X1 NOR2X1_1661 ( .gnd(gnd), .vdd(vdd), .A(_10359_), .B(_10300_), .Y(_10360_) );
OAI21X1 OAI21X1_2916 ( .gnd(gnd), .vdd(vdd), .A(_10360_), .B(_10352_), .C(_10355_), .Y(_10361_) );
OAI21X1 OAI21X1_2917 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_5_bF_buf3_), .B(micro_hash_ucr_3_a_5_bF_buf0_), .C(_10361_), .Y(_10362_) );
AOI21X1 AOI21X1_1838 ( .gnd(gnd), .vdd(vdd), .A(_10362_), .B(_10358_), .C(_8800__bF_buf9), .Y(_8778__5_) );
AOI21X1 AOI21X1_1839 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_6_bF_buf0_), .B(micro_hash_ucr_3_a_6_bF_buf0_), .C(_10274_), .Y(_10363_) );
OAI22X1 OAI22X1_128 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_6_bF_buf3_), .B(micro_hash_ucr_3_a_6_bF_buf3_), .C(_10363_), .D(_10356_), .Y(_10364_) );
NAND2X1 NAND2X1_1382 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_x_6_), .B(_10357_), .Y(_10365_) );
AOI21X1 AOI21X1_1840 ( .gnd(gnd), .vdd(vdd), .A(_10365_), .B(_10364_), .C(_8800__bF_buf8), .Y(_8778__6_) );
AOI21X1 AOI21X1_1841 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_7_bF_buf0_), .B(micro_hash_ucr_3_a_7_bF_buf2_), .C(_10274_), .Y(_10366_) );
OAI22X1 OAI22X1_129 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_7_bF_buf3_), .B(micro_hash_ucr_3_a_7_bF_buf1_), .C(_10366_), .D(_10356_), .Y(_10367_) );
NAND3X1 NAND3X1_574 ( .gnd(gnd), .vdd(vdd), .A(_9326__bF_buf1), .B(_9332_), .C(_9338_), .Y(_10368_) );
NAND3X1 NAND3X1_575 ( .gnd(gnd), .vdd(vdd), .A(_10260_), .B(_10269_), .C(_9373_), .Y(_10369_) );
NOR2X1 NOR2X1_1662 ( .gnd(gnd), .vdd(vdd), .A(_10368_), .B(_10369_), .Y(_10370_) );
INVX1 INVX1_638 ( .gnd(gnd), .vdd(vdd), .A(_10286_), .Y(_10371_) );
NOR2X1 NOR2X1_1663 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe35_bF_buf0), .B(_10346_), .Y(_10372_) );
NAND3X1 NAND3X1_576 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_x_7_), .B(_10287_), .C(_10372_), .Y(_10373_) );
NOR2X1 NOR2X1_1664 ( .gnd(gnd), .vdd(vdd), .A(_10373_), .B(_10371_), .Y(_10374_) );
NOR2X1 NOR2X1_1665 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe15_bF_buf2), .B(micro_hash_ucr_3_pipe13), .Y(_10375_) );
NOR2X1 NOR2X1_1666 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe29_bF_buf0), .B(micro_hash_ucr_3_pipe21_bF_buf0), .Y(_10376_) );
NAND3X1 NAND3X1_577 ( .gnd(gnd), .vdd(vdd), .A(_9333__bF_buf0), .B(_10375_), .C(_10376_), .Y(_10377_) );
NOR2X1 NOR2X1_1667 ( .gnd(gnd), .vdd(vdd), .A(_10377_), .B(_10354_), .Y(_10378_) );
NAND3X1 NAND3X1_578 ( .gnd(gnd), .vdd(vdd), .A(_10370_), .B(_10378_), .C(_10374_), .Y(_10379_) );
AOI21X1 AOI21X1_1842 ( .gnd(gnd), .vdd(vdd), .A(_10379_), .B(_10367_), .C(_8800__bF_buf7), .Y(_8778__7_) );
NOR2X1 NOR2X1_1668 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe69), .B(_8800__bF_buf6), .Y(_10380_) );
INVX8 INVX8_276 ( .gnd(gnd), .vdd(vdd), .A(_10380_), .Y(_10381_) );
INVX1 INVX1_639 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_232_), .Y(_10382_) );
NOR2X1 NOR2X1_1669 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_k_0_), .B(micro_hash_ucr_3_x_0_), .Y(_10383_) );
NOR2X1 NOR2X1_1670 ( .gnd(gnd), .vdd(vdd), .A(_10249_), .B(_10293_), .Y(_10384_) );
OAI21X1 OAI21X1_2918 ( .gnd(gnd), .vdd(vdd), .A(_10384_), .B(_10383_), .C(_10382_), .Y(_10385_) );
NOR2X1 NOR2X1_1671 ( .gnd(gnd), .vdd(vdd), .A(_10383_), .B(_10384_), .Y(_10386_) );
INVX8 INVX8_277 ( .gnd(gnd), .vdd(vdd), .A(_10386__bF_buf5), .Y(_10387_) );
NOR2X1 NOR2X1_1672 ( .gnd(gnd), .vdd(vdd), .A(_10382_), .B(_10387__bF_buf3), .Y(_10388_) );
INVX1 INVX1_640 ( .gnd(gnd), .vdd(vdd), .A(_10388_), .Y(_10389_) );
NAND2X1 NAND2X1_1383 ( .gnd(gnd), .vdd(vdd), .A(_10385_), .B(_10389_), .Y(_10390_) );
XNOR2X1 XNOR2X1_391 ( .gnd(gnd), .vdd(vdd), .A(_10386__bF_buf4), .B(micro_hash_ucr_3_Wx_168_), .Y(_10391_) );
NOR2X1 NOR2X1_1673 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_8_), .B(_10386__bF_buf3), .Y(_10392_) );
NAND2X1 NAND2X1_1384 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_8_), .B(_10386__bF_buf2), .Y(_10393_) );
INVX1 INVX1_641 ( .gnd(gnd), .vdd(vdd), .A(_10393_), .Y(_10394_) );
OAI21X1 OAI21X1_2919 ( .gnd(gnd), .vdd(vdd), .A(_10394_), .B(_10392_), .C(micro_hash_ucr_3_pipe10_bF_buf2), .Y(_10395_) );
NAND2X1 NAND2X1_1385 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_0_), .B(_10386__bF_buf1), .Y(_10396_) );
INVX2 INVX2_363 ( .gnd(gnd), .vdd(vdd), .A(_10396_), .Y(_10397_) );
NOR2X1 NOR2X1_1674 ( .gnd(gnd), .vdd(vdd), .A(_9341_), .B(_10397_), .Y(_10398_) );
OAI21X1 OAI21X1_2920 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_0_), .B(_10386__bF_buf0), .C(_10398_), .Y(_10399_) );
NAND2X1 NAND2X1_1386 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe6_bF_buf3), .B(_12847_), .Y(_10400_) );
OAI21X1 OAI21X1_2921 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_0_), .B(micro_hash_ucr_3_pipe6_bF_buf2), .C(_10400_), .Y(_10401_) );
OAI21X1 OAI21X1_2922 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe8), .B(_10401_), .C(_10399_), .Y(_10402_) );
OAI21X1 OAI21X1_2923 ( .gnd(gnd), .vdd(vdd), .A(_10402_), .B(micro_hash_ucr_3_pipe10_bF_buf1), .C(_10395_), .Y(_10403_) );
XNOR2X1 XNOR2X1_392 ( .gnd(gnd), .vdd(vdd), .A(_10386__bF_buf5), .B(micro_hash_ucr_3_Wx_16_), .Y(_10404_) );
MUX2X1 MUX2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_10403_), .B(_10404_), .S(_9340_), .Y(_10405_) );
XOR2X1 XOR2X1_165 ( .gnd(gnd), .vdd(vdd), .A(_10386__bF_buf4), .B(micro_hash_ucr_3_Wx_24_), .Y(_10406_) );
MUX2X1 MUX2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_10405_), .B(_10406_), .S(_9335__bF_buf0), .Y(_10407_) );
INVX1 INVX1_642 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_32_), .Y(_10408_) );
NOR2X1 NOR2X1_1675 ( .gnd(gnd), .vdd(vdd), .A(_10408_), .B(_10387__bF_buf2), .Y(_10409_) );
NOR2X1 NOR2X1_1676 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_32_), .B(_10386__bF_buf3), .Y(_10410_) );
NOR2X1 NOR2X1_1677 ( .gnd(gnd), .vdd(vdd), .A(_10410_), .B(_10409_), .Y(_10411_) );
AOI21X1 AOI21X1_1843 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe16_bF_buf0), .B(_10411_), .C(micro_hash_ucr_3_pipe18_bF_buf1), .Y(_10412_) );
OAI21X1 OAI21X1_2924 ( .gnd(gnd), .vdd(vdd), .A(_10407_), .B(micro_hash_ucr_3_pipe16_bF_buf4), .C(_10412_), .Y(_10413_) );
NOR2X1 NOR2X1_1678 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_40_), .B(_10386__bF_buf2), .Y(_10414_) );
INVX1 INVX1_643 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_40_), .Y(_10415_) );
NOR2X1 NOR2X1_1679 ( .gnd(gnd), .vdd(vdd), .A(_10415_), .B(_10387__bF_buf1), .Y(_10416_) );
OAI21X1 OAI21X1_2925 ( .gnd(gnd), .vdd(vdd), .A(_10416_), .B(_10414_), .C(micro_hash_ucr_3_pipe18_bF_buf0), .Y(_10417_) );
NAND3X1 NAND3X1_579 ( .gnd(gnd), .vdd(vdd), .A(_9329__bF_buf1), .B(_10417_), .C(_10413_), .Y(_10418_) );
INVX1 INVX1_644 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_48_), .Y(_10419_) );
NOR2X1 NOR2X1_1680 ( .gnd(gnd), .vdd(vdd), .A(_10419_), .B(_10387__bF_buf0), .Y(_10420_) );
OAI21X1 OAI21X1_2926 ( .gnd(gnd), .vdd(vdd), .A(_10386__bF_buf1), .B(micro_hash_ucr_3_Wx_48_), .C(micro_hash_ucr_3_pipe20_bF_buf3), .Y(_10421_) );
OAI21X1 OAI21X1_2927 ( .gnd(gnd), .vdd(vdd), .A(_10420_), .B(_10421_), .C(_10418_), .Y(_10422_) );
NOR2X1 NOR2X1_1681 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_56_), .B(_10386__bF_buf0), .Y(_10423_) );
NOR2X1 NOR2X1_1682 ( .gnd(gnd), .vdd(vdd), .A(_9260_), .B(_10387__bF_buf3), .Y(_10424_) );
OAI21X1 OAI21X1_2928 ( .gnd(gnd), .vdd(vdd), .A(_10424_), .B(_10423_), .C(micro_hash_ucr_3_pipe22_bF_buf3), .Y(_10425_) );
OAI21X1 OAI21X1_2929 ( .gnd(gnd), .vdd(vdd), .A(_10422_), .B(micro_hash_ucr_3_pipe22_bF_buf2), .C(_10425_), .Y(_10426_) );
NOR2X1 NOR2X1_1683 ( .gnd(gnd), .vdd(vdd), .A(_9237_), .B(_10387__bF_buf2), .Y(_10427_) );
OAI21X1 OAI21X1_2930 ( .gnd(gnd), .vdd(vdd), .A(_10386__bF_buf5), .B(micro_hash_ucr_3_Wx_64_), .C(micro_hash_ucr_3_pipe24_bF_buf0), .Y(_10428_) );
OAI22X1 OAI22X1_130 ( .gnd(gnd), .vdd(vdd), .A(_10427_), .B(_10428_), .C(_10426_), .D(micro_hash_ucr_3_pipe24_bF_buf4), .Y(_10429_) );
OAI21X1 OAI21X1_2931 ( .gnd(gnd), .vdd(vdd), .A(_10384_), .B(_10383_), .C(_9159_), .Y(_10430_) );
NOR2X1 NOR2X1_1684 ( .gnd(gnd), .vdd(vdd), .A(_9159_), .B(_10387__bF_buf1), .Y(_10431_) );
INVX1 INVX1_645 ( .gnd(gnd), .vdd(vdd), .A(_10431_), .Y(_10432_) );
NAND2X1 NAND2X1_1387 ( .gnd(gnd), .vdd(vdd), .A(_10430_), .B(_10432_), .Y(_10433_) );
AOI21X1 AOI21X1_1844 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe26_bF_buf4), .B(_10433_), .C(micro_hash_ucr_3_pipe28_bF_buf2), .Y(_10434_) );
OAI21X1 OAI21X1_2932 ( .gnd(gnd), .vdd(vdd), .A(_10429_), .B(micro_hash_ucr_3_pipe26_bF_buf3), .C(_10434_), .Y(_10435_) );
NOR2X1 NOR2X1_1685 ( .gnd(gnd), .vdd(vdd), .A(_9214_), .B(_10387__bF_buf0), .Y(_10436_) );
OAI21X1 OAI21X1_2933 ( .gnd(gnd), .vdd(vdd), .A(_10386__bF_buf4), .B(micro_hash_ucr_3_Wx_80_), .C(micro_hash_ucr_3_pipe28_bF_buf1), .Y(_10437_) );
OAI21X1 OAI21X1_2934 ( .gnd(gnd), .vdd(vdd), .A(_10436_), .B(_10437_), .C(_10435_), .Y(_10438_) );
NOR2X1 NOR2X1_1686 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_88_), .B(_10386__bF_buf3), .Y(_10439_) );
NOR2X1 NOR2X1_1687 ( .gnd(gnd), .vdd(vdd), .A(_9182_), .B(_10387__bF_buf3), .Y(_10440_) );
OAI21X1 OAI21X1_2935 ( .gnd(gnd), .vdd(vdd), .A(_10440_), .B(_10439_), .C(micro_hash_ucr_3_pipe30_bF_buf1), .Y(_10441_) );
OAI21X1 OAI21X1_2936 ( .gnd(gnd), .vdd(vdd), .A(_10438_), .B(micro_hash_ucr_3_pipe30_bF_buf0), .C(_10441_), .Y(_10442_) );
NOR2X1 NOR2X1_1688 ( .gnd(gnd), .vdd(vdd), .A(_9040_), .B(_10387__bF_buf2), .Y(_10443_) );
OAI21X1 OAI21X1_2937 ( .gnd(gnd), .vdd(vdd), .A(_10386__bF_buf2), .B(micro_hash_ucr_3_Wx_96_), .C(micro_hash_ucr_3_pipe32_bF_buf0), .Y(_10444_) );
OAI22X1 OAI22X1_131 ( .gnd(gnd), .vdd(vdd), .A(_10443_), .B(_10444_), .C(_10442_), .D(micro_hash_ucr_3_pipe32_bF_buf3), .Y(_10445_) );
XNOR2X1 XNOR2X1_393 ( .gnd(gnd), .vdd(vdd), .A(_10386__bF_buf1), .B(micro_hash_ucr_3_Wx_104_), .Y(_10446_) );
AOI21X1 AOI21X1_1845 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe34_bF_buf0), .B(_10446_), .C(micro_hash_ucr_3_pipe36_bF_buf1), .Y(_10447_) );
OAI21X1 OAI21X1_2938 ( .gnd(gnd), .vdd(vdd), .A(_10445_), .B(micro_hash_ucr_3_pipe34_bF_buf4), .C(_10447_), .Y(_10448_) );
NOR2X1 NOR2X1_1689 ( .gnd(gnd), .vdd(vdd), .A(_9114_), .B(_10387__bF_buf1), .Y(_10449_) );
OAI21X1 OAI21X1_2939 ( .gnd(gnd), .vdd(vdd), .A(_10386__bF_buf0), .B(micro_hash_ucr_3_Wx_112_), .C(micro_hash_ucr_3_pipe36_bF_buf0), .Y(_10450_) );
OAI21X1 OAI21X1_2940 ( .gnd(gnd), .vdd(vdd), .A(_10449_), .B(_10450_), .C(_10448_), .Y(_10451_) );
NOR2X1 NOR2X1_1690 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_120_), .B(_10386__bF_buf5), .Y(_10452_) );
NOR2X1 NOR2X1_1691 ( .gnd(gnd), .vdd(vdd), .A(_9018_), .B(_10387__bF_buf0), .Y(_10453_) );
OAI21X1 OAI21X1_2941 ( .gnd(gnd), .vdd(vdd), .A(_10453_), .B(_10452_), .C(micro_hash_ucr_3_pipe38_bF_buf0), .Y(_10454_) );
OAI21X1 OAI21X1_2942 ( .gnd(gnd), .vdd(vdd), .A(_10451_), .B(micro_hash_ucr_3_pipe38_bF_buf3), .C(_10454_), .Y(_10455_) );
NOR2X1 NOR2X1_1692 ( .gnd(gnd), .vdd(vdd), .A(_9068_), .B(_10387__bF_buf3), .Y(_10456_) );
NOR2X1 NOR2X1_1693 ( .gnd(gnd), .vdd(vdd), .A(_9312__bF_buf3), .B(_10456_), .Y(_10457_) );
OAI21X1 OAI21X1_2943 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_128_), .B(_10386__bF_buf4), .C(_10457_), .Y(_10458_) );
OAI21X1 OAI21X1_2944 ( .gnd(gnd), .vdd(vdd), .A(_10455_), .B(micro_hash_ucr_3_pipe40_bF_buf0), .C(_10458_), .Y(_10459_) );
NOR2X1 NOR2X1_1694 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_136_), .B(_10386__bF_buf3), .Y(_10460_) );
NOR2X1 NOR2X1_1695 ( .gnd(gnd), .vdd(vdd), .A(_9183_), .B(_10387__bF_buf2), .Y(_10461_) );
OAI21X1 OAI21X1_2945 ( .gnd(gnd), .vdd(vdd), .A(_10461_), .B(_10460_), .C(micro_hash_ucr_3_pipe42_bF_buf0), .Y(_10462_) );
AND2X2 AND2X2_691 ( .gnd(gnd), .vdd(vdd), .A(_10462_), .B(_9305__bF_buf0), .Y(_10463_) );
OAI21X1 OAI21X1_2946 ( .gnd(gnd), .vdd(vdd), .A(_10459_), .B(micro_hash_ucr_3_pipe42_bF_buf3), .C(_10463_), .Y(_10464_) );
NOR2X1 NOR2X1_1696 ( .gnd(gnd), .vdd(vdd), .A(_8932_), .B(_10387__bF_buf1), .Y(_10465_) );
OAI21X1 OAI21X1_2947 ( .gnd(gnd), .vdd(vdd), .A(_10386__bF_buf2), .B(micro_hash_ucr_3_Wx_144_), .C(micro_hash_ucr_3_pipe44_bF_buf2), .Y(_10466_) );
OAI21X1 OAI21X1_2948 ( .gnd(gnd), .vdd(vdd), .A(_10465_), .B(_10466_), .C(_10464_), .Y(_10467_) );
NOR2X1 NOR2X1_1697 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_152_), .B(_10386__bF_buf1), .Y(_10468_) );
NOR2X1 NOR2X1_1698 ( .gnd(gnd), .vdd(vdd), .A(_8991_), .B(_10387__bF_buf0), .Y(_10469_) );
OAI21X1 OAI21X1_2949 ( .gnd(gnd), .vdd(vdd), .A(_10469_), .B(_10468_), .C(micro_hash_ucr_3_pipe46_bF_buf0), .Y(_10470_) );
OAI21X1 OAI21X1_2950 ( .gnd(gnd), .vdd(vdd), .A(_10467_), .B(micro_hash_ucr_3_pipe46_bF_buf4), .C(_10470_), .Y(_10471_) );
NOR2X1 NOR2X1_1699 ( .gnd(gnd), .vdd(vdd), .A(_8962_), .B(_10387__bF_buf3), .Y(_10472_) );
OAI21X1 OAI21X1_2951 ( .gnd(gnd), .vdd(vdd), .A(_10386__bF_buf0), .B(micro_hash_ucr_3_Wx_160_), .C(micro_hash_ucr_3_pipe48_bF_buf4), .Y(_10473_) );
OAI22X1 OAI22X1_132 ( .gnd(gnd), .vdd(vdd), .A(_10472_), .B(_10473_), .C(_10471_), .D(micro_hash_ucr_3_pipe48_bF_buf3), .Y(_10474_) );
NAND2X1 NAND2X1_1388 ( .gnd(gnd), .vdd(vdd), .A(_9299__bF_buf1), .B(_10474_), .Y(_10475_) );
OAI21X1 OAI21X1_2952 ( .gnd(gnd), .vdd(vdd), .A(_9299__bF_buf0), .B(_10391_), .C(_10475_), .Y(_10476_) );
NOR2X1 NOR2X1_1700 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_176_), .B(_10386__bF_buf5), .Y(_10477_) );
NOR2X1 NOR2X1_1701 ( .gnd(gnd), .vdd(vdd), .A(_9069_), .B(_10387__bF_buf2), .Y(_10478_) );
OAI21X1 OAI21X1_2953 ( .gnd(gnd), .vdd(vdd), .A(_10478_), .B(_10477_), .C(micro_hash_ucr_3_pipe52_bF_buf1), .Y(_10479_) );
OAI21X1 OAI21X1_2954 ( .gnd(gnd), .vdd(vdd), .A(_10476_), .B(micro_hash_ucr_3_pipe52_bF_buf0), .C(_10479_), .Y(_10480_) );
NOR2X1 NOR2X1_1702 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_184_), .B(_10386__bF_buf4), .Y(_10481_) );
AND2X2 AND2X2_692 ( .gnd(gnd), .vdd(vdd), .A(_10386__bF_buf3), .B(micro_hash_ucr_3_Wx_184_), .Y(_10482_) );
OAI21X1 OAI21X1_2955 ( .gnd(gnd), .vdd(vdd), .A(_10482_), .B(_10481_), .C(micro_hash_ucr_3_pipe54_bF_buf3), .Y(_10483_) );
NAND2X1 NAND2X1_1389 ( .gnd(gnd), .vdd(vdd), .A(_9293__bF_buf3), .B(_10483_), .Y(_10484_) );
AOI21X1 AOI21X1_1846 ( .gnd(gnd), .vdd(vdd), .A(_9298__bF_buf4), .B(_10480_), .C(_10484_), .Y(_10485_) );
NOR2X1 NOR2X1_1703 ( .gnd(gnd), .vdd(vdd), .A(_8933_), .B(_10387__bF_buf1), .Y(_10486_) );
OAI21X1 OAI21X1_2956 ( .gnd(gnd), .vdd(vdd), .A(_10386__bF_buf2), .B(micro_hash_ucr_3_Wx_192_), .C(micro_hash_ucr_3_pipe56_bF_buf4), .Y(_10487_) );
OAI21X1 OAI21X1_2957 ( .gnd(gnd), .vdd(vdd), .A(_10486_), .B(_10487_), .C(_9294__bF_buf0), .Y(_10488_) );
XOR2X1 XOR2X1_166 ( .gnd(gnd), .vdd(vdd), .A(_10386__bF_buf1), .B(micro_hash_ucr_3_Wx_200_), .Y(_10489_) );
OAI22X1 OAI22X1_133 ( .gnd(gnd), .vdd(vdd), .A(_9294__bF_buf4), .B(_10489_), .C(_10485_), .D(_10488_), .Y(_10490_) );
NOR2X1 NOR2X1_1704 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe60_bF_buf4), .B(_10490_), .Y(_10491_) );
NOR2X1 NOR2X1_1705 ( .gnd(gnd), .vdd(vdd), .A(_8963_), .B(_10387__bF_buf0), .Y(_10492_) );
OAI21X1 OAI21X1_2958 ( .gnd(gnd), .vdd(vdd), .A(_10386__bF_buf0), .B(micro_hash_ucr_3_Wx_208_), .C(micro_hash_ucr_3_pipe60_bF_buf3), .Y(_10493_) );
OAI21X1 OAI21X1_2959 ( .gnd(gnd), .vdd(vdd), .A(_10492_), .B(_10493_), .C(_9287__bF_buf4), .Y(_10494_) );
NOR2X1 NOR2X1_1706 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_216_), .B(_10386__bF_buf5), .Y(_10495_) );
NOR2X1 NOR2X1_1707 ( .gnd(gnd), .vdd(vdd), .A(_8834_), .B(_10387__bF_buf3), .Y(_10496_) );
OAI21X1 OAI21X1_2960 ( .gnd(gnd), .vdd(vdd), .A(_10496_), .B(_10495_), .C(micro_hash_ucr_3_pipe62_bF_buf3), .Y(_10497_) );
AND2X2 AND2X2_693 ( .gnd(gnd), .vdd(vdd), .A(_10497_), .B(_9288__bF_buf3), .Y(_10498_) );
OAI21X1 OAI21X1_2961 ( .gnd(gnd), .vdd(vdd), .A(_10491_), .B(_10494_), .C(_10498_), .Y(_10499_) );
AND2X2 AND2X2_694 ( .gnd(gnd), .vdd(vdd), .A(_10386__bF_buf4), .B(micro_hash_ucr_3_Wx_224_), .Y(_10500_) );
OAI21X1 OAI21X1_2962 ( .gnd(gnd), .vdd(vdd), .A(_10386__bF_buf3), .B(micro_hash_ucr_3_Wx_224_), .C(micro_hash_ucr_3_pipe64_bF_buf4), .Y(_10501_) );
OAI21X1 OAI21X1_2963 ( .gnd(gnd), .vdd(vdd), .A(_10500_), .B(_10501_), .C(_10499_), .Y(_10502_) );
NAND2X1 NAND2X1_1390 ( .gnd(gnd), .vdd(vdd), .A(_9286__bF_buf3), .B(_10502_), .Y(_10503_) );
OAI21X1 OAI21X1_2964 ( .gnd(gnd), .vdd(vdd), .A(_9286__bF_buf2), .B(_10390_), .C(_10503_), .Y(_10504_) );
NOR2X1 NOR2X1_1708 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_240_), .B(_10386__bF_buf2), .Y(_10505_) );
AND2X2 AND2X2_695 ( .gnd(gnd), .vdd(vdd), .A(_10386__bF_buf1), .B(micro_hash_ucr_3_Wx_240_), .Y(_10506_) );
OAI21X1 OAI21X1_2965 ( .gnd(gnd), .vdd(vdd), .A(_10506_), .B(_10505_), .C(micro_hash_ucr_3_pipe68_bF_buf3), .Y(_10507_) );
OAI21X1 OAI21X1_2966 ( .gnd(gnd), .vdd(vdd), .A(_10504_), .B(micro_hash_ucr_3_pipe68_bF_buf2), .C(_10507_), .Y(_10508_) );
INVX2 INVX2_364 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_248_), .Y(_10509_) );
AOI21X1 AOI21X1_1847 ( .gnd(gnd), .vdd(vdd), .A(_10509_), .B(_10387__bF_buf2), .C(_8800__bF_buf5), .Y(_10510_) );
OAI21X1 OAI21X1_2967 ( .gnd(gnd), .vdd(vdd), .A(_10509_), .B(_10387__bF_buf1), .C(_10510_), .Y(_10511_) );
AOI22X1 AOI22X1_74 ( .gnd(gnd), .vdd(vdd), .A(_10381_), .B(_10511_), .C(_10508_), .D(_9283__bF_buf0), .Y(_8702__0_) );
NOR2X1 NOR2X1_1709 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_k_1_), .B(micro_hash_ucr_3_x_1_), .Y(_10512_) );
INVX1 INVX1_646 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_k_1_), .Y(_10513_) );
INVX1 INVX1_647 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_x_1_), .Y(_10514_) );
NOR2X1 NOR2X1_1710 ( .gnd(gnd), .vdd(vdd), .A(_10513_), .B(_10514_), .Y(_10515_) );
NOR2X1 NOR2X1_1711 ( .gnd(gnd), .vdd(vdd), .A(_10512_), .B(_10515_), .Y(_10516_) );
NAND2X1 NAND2X1_1391 ( .gnd(gnd), .vdd(vdd), .A(_10384_), .B(_10516_), .Y(_10517_) );
OR2X2 OR2X2_72 ( .gnd(gnd), .vdd(vdd), .A(_10516_), .B(_10384_), .Y(_10518_) );
NAND2X1 NAND2X1_1392 ( .gnd(gnd), .vdd(vdd), .A(_10517_), .B(_10518_), .Y(_10519_) );
XNOR2X1 XNOR2X1_394 ( .gnd(gnd), .vdd(vdd), .A(_10519__bF_buf5), .B(micro_hash_ucr_3_Wx_217_), .Y(_10520_) );
XNOR2X1 XNOR2X1_395 ( .gnd(gnd), .vdd(vdd), .A(_10520_), .B(_10496_), .Y(_10521_) );
INVX8 INVX8_278 ( .gnd(gnd), .vdd(vdd), .A(_10519__bF_buf4), .Y(_10522_) );
NOR2X1 NOR2X1_1712 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_153_), .B(_10522__bF_buf4), .Y(_10523_) );
NOR2X1 NOR2X1_1713 ( .gnd(gnd), .vdd(vdd), .A(_8994_), .B(_10519__bF_buf3), .Y(_10524_) );
NOR2X1 NOR2X1_1714 ( .gnd(gnd), .vdd(vdd), .A(_10524_), .B(_10523_), .Y(_10525_) );
XNOR2X1 XNOR2X1_396 ( .gnd(gnd), .vdd(vdd), .A(_10525_), .B(_10469_), .Y(_10526_) );
NOR2X1 NOR2X1_1715 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_121_), .B(_10522__bF_buf3), .Y(_10527_) );
NOR2X1 NOR2X1_1716 ( .gnd(gnd), .vdd(vdd), .A(_9021_), .B(_10519__bF_buf2), .Y(_10528_) );
NOR2X1 NOR2X1_1717 ( .gnd(gnd), .vdd(vdd), .A(_10528_), .B(_10527_), .Y(_10529_) );
XNOR2X1 XNOR2X1_397 ( .gnd(gnd), .vdd(vdd), .A(_10529_), .B(_10453_), .Y(_10530_) );
INVX2 INVX2_365 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_9_), .Y(_10531_) );
XNOR2X1 XNOR2X1_398 ( .gnd(gnd), .vdd(vdd), .A(_10519__bF_buf1), .B(_10531_), .Y(_10532_) );
OR2X2 OR2X2_73 ( .gnd(gnd), .vdd(vdd), .A(_10532_), .B(_10393_), .Y(_10533_) );
AOI21X1 AOI21X1_1848 ( .gnd(gnd), .vdd(vdd), .A(_10393_), .B(_10532_), .C(_9342_), .Y(_10534_) );
XNOR2X1 XNOR2X1_399 ( .gnd(gnd), .vdd(vdd), .A(_10519__bF_buf0), .B(micro_hash_ucr_3_Wx_1_), .Y(_10535_) );
NOR2X1 NOR2X1_1718 ( .gnd(gnd), .vdd(vdd), .A(_10397_), .B(_10535_), .Y(_10536_) );
AND2X2 AND2X2_696 ( .gnd(gnd), .vdd(vdd), .A(_10535_), .B(_10397_), .Y(_10537_) );
OAI21X1 OAI21X1_2968 ( .gnd(gnd), .vdd(vdd), .A(_10537_), .B(_10536_), .C(micro_hash_ucr_3_pipe8), .Y(_10538_) );
NAND2X1 NAND2X1_1393 ( .gnd(gnd), .vdd(vdd), .A(_9483_), .B(_9345_), .Y(_10539_) );
OAI21X1 OAI21X1_2969 ( .gnd(gnd), .vdd(vdd), .A(H_3_17_), .B(_9345_), .C(_10539_), .Y(_10540_) );
AOI21X1 AOI21X1_1849 ( .gnd(gnd), .vdd(vdd), .A(_9341_), .B(_10540_), .C(micro_hash_ucr_3_pipe10_bF_buf0), .Y(_10541_) );
AOI22X1 AOI22X1_75 ( .gnd(gnd), .vdd(vdd), .A(_10533_), .B(_10534_), .C(_10538_), .D(_10541_), .Y(_10542_) );
AND2X2 AND2X2_697 ( .gnd(gnd), .vdd(vdd), .A(_10386__bF_buf0), .B(micro_hash_ucr_3_Wx_16_), .Y(_10543_) );
XNOR2X1 XNOR2X1_400 ( .gnd(gnd), .vdd(vdd), .A(_10519__bF_buf5), .B(micro_hash_ucr_3_Wx_17_), .Y(_10544_) );
XNOR2X1 XNOR2X1_401 ( .gnd(gnd), .vdd(vdd), .A(_10544_), .B(_10543_), .Y(_10545_) );
MUX2X1 MUX2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_10542_), .B(_10545_), .S(_9340_), .Y(_10546_) );
NAND2X1 NAND2X1_1394 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_24_), .B(_10386__bF_buf5), .Y(_10547_) );
XOR2X1 XOR2X1_167 ( .gnd(gnd), .vdd(vdd), .A(_10519__bF_buf4), .B(micro_hash_ucr_3_Wx_25_), .Y(_10548_) );
AND2X2 AND2X2_698 ( .gnd(gnd), .vdd(vdd), .A(_10548_), .B(_10547_), .Y(_10549_) );
NOR2X1 NOR2X1_1719 ( .gnd(gnd), .vdd(vdd), .A(_10547_), .B(_10548_), .Y(_10550_) );
OAI21X1 OAI21X1_2970 ( .gnd(gnd), .vdd(vdd), .A(_10549_), .B(_10550_), .C(micro_hash_ucr_3_pipe14_bF_buf0), .Y(_10551_) );
OAI21X1 OAI21X1_2971 ( .gnd(gnd), .vdd(vdd), .A(_10546_), .B(micro_hash_ucr_3_pipe14_bF_buf3), .C(_10551_), .Y(_10552_) );
INVX2 INVX2_366 ( .gnd(gnd), .vdd(vdd), .A(_10409_), .Y(_10553_) );
NOR2X1 NOR2X1_1720 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_33_), .B(_10522__bF_buf2), .Y(_10554_) );
NAND2X1 NAND2X1_1395 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_33_), .B(_10522__bF_buf1), .Y(_10555_) );
INVX1 INVX1_648 ( .gnd(gnd), .vdd(vdd), .A(_10555_), .Y(_10556_) );
NOR2X1 NOR2X1_1721 ( .gnd(gnd), .vdd(vdd), .A(_10554_), .B(_10556_), .Y(_10557_) );
XNOR2X1 XNOR2X1_402 ( .gnd(gnd), .vdd(vdd), .A(_10557_), .B(_10553_), .Y(_10558_) );
AOI21X1 AOI21X1_1850 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe16_bF_buf3), .B(_10558_), .C(micro_hash_ucr_3_pipe18_bF_buf4), .Y(_10559_) );
OAI21X1 OAI21X1_2972 ( .gnd(gnd), .vdd(vdd), .A(_10552_), .B(micro_hash_ucr_3_pipe16_bF_buf2), .C(_10559_), .Y(_10560_) );
INVX2 INVX2_367 ( .gnd(gnd), .vdd(vdd), .A(_10420_), .Y(_10561_) );
NOR2X1 NOR2X1_1722 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_49_), .B(_10522__bF_buf0), .Y(_10562_) );
NAND2X1 NAND2X1_1396 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_49_), .B(_10522__bF_buf4), .Y(_10563_) );
INVX1 INVX1_649 ( .gnd(gnd), .vdd(vdd), .A(_10563_), .Y(_10564_) );
NOR2X1 NOR2X1_1723 ( .gnd(gnd), .vdd(vdd), .A(_10562_), .B(_10564_), .Y(_10565_) );
XNOR2X1 XNOR2X1_403 ( .gnd(gnd), .vdd(vdd), .A(_10565_), .B(_10561_), .Y(_10566_) );
NOR2X1 NOR2X1_1724 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_41_), .B(_10522__bF_buf3), .Y(_10567_) );
NAND2X1 NAND2X1_1397 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_41_), .B(_10522__bF_buf2), .Y(_10568_) );
INVX1 INVX1_650 ( .gnd(gnd), .vdd(vdd), .A(_10568_), .Y(_10569_) );
NOR2X1 NOR2X1_1725 ( .gnd(gnd), .vdd(vdd), .A(_10567_), .B(_10569_), .Y(_10570_) );
XNOR2X1 XNOR2X1_404 ( .gnd(gnd), .vdd(vdd), .A(_10570_), .B(_10416_), .Y(_10571_) );
AOI21X1 AOI21X1_1851 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe18_bF_buf3), .B(_10571_), .C(micro_hash_ucr_3_pipe20_bF_buf2), .Y(_10572_) );
AOI22X1 AOI22X1_76 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe20_bF_buf1), .B(_10566_), .C(_10560_), .D(_10572_), .Y(_10573_) );
NAND2X1 NAND2X1_1398 ( .gnd(gnd), .vdd(vdd), .A(_9330__bF_buf1), .B(_10573_), .Y(_10574_) );
NOR2X1 NOR2X1_1726 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_57_), .B(_10522__bF_buf1), .Y(_10575_) );
NOR2X1 NOR2X1_1727 ( .gnd(gnd), .vdd(vdd), .A(_9263_), .B(_10519__bF_buf3), .Y(_10576_) );
NOR2X1 NOR2X1_1728 ( .gnd(gnd), .vdd(vdd), .A(_10576_), .B(_10575_), .Y(_10577_) );
XOR2X1 XOR2X1_168 ( .gnd(gnd), .vdd(vdd), .A(_10577_), .B(_10424_), .Y(_10578_) );
OAI21X1 OAI21X1_2973 ( .gnd(gnd), .vdd(vdd), .A(_9330__bF_buf0), .B(_10578_), .C(_10574_), .Y(_10579_) );
XNOR2X1 XNOR2X1_405 ( .gnd(gnd), .vdd(vdd), .A(_10519__bF_buf2), .B(micro_hash_ucr_3_Wx_65_), .Y(_10580_) );
XOR2X1 XOR2X1_169 ( .gnd(gnd), .vdd(vdd), .A(_10580_), .B(_10427_), .Y(_10581_) );
AOI21X1 AOI21X1_1852 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe24_bF_buf3), .B(_10581_), .C(micro_hash_ucr_3_pipe26_bF_buf2), .Y(_10582_) );
OAI21X1 OAI21X1_2974 ( .gnd(gnd), .vdd(vdd), .A(_10579_), .B(micro_hash_ucr_3_pipe24_bF_buf2), .C(_10582_), .Y(_10583_) );
NOR2X1 NOR2X1_1729 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_73_), .B(_10522__bF_buf0), .Y(_10584_) );
NOR2X1 NOR2X1_1730 ( .gnd(gnd), .vdd(vdd), .A(_9162_), .B(_10519__bF_buf1), .Y(_10585_) );
NOR2X1 NOR2X1_1731 ( .gnd(gnd), .vdd(vdd), .A(_10585_), .B(_10584_), .Y(_10586_) );
NAND2X1 NAND2X1_1399 ( .gnd(gnd), .vdd(vdd), .A(_10431_), .B(_10586_), .Y(_10587_) );
OAI21X1 OAI21X1_2975 ( .gnd(gnd), .vdd(vdd), .A(_10584_), .B(_10585_), .C(_10432_), .Y(_10588_) );
NAND2X1 NAND2X1_1400 ( .gnd(gnd), .vdd(vdd), .A(_10588_), .B(_10587_), .Y(_10589_) );
AOI21X1 AOI21X1_1853 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe26_bF_buf1), .B(_10589_), .C(micro_hash_ucr_3_pipe28_bF_buf0), .Y(_10590_) );
XNOR2X1 XNOR2X1_406 ( .gnd(gnd), .vdd(vdd), .A(_10519__bF_buf0), .B(micro_hash_ucr_3_Wx_81_), .Y(_10591_) );
NAND2X1 NAND2X1_1401 ( .gnd(gnd), .vdd(vdd), .A(_10436_), .B(_10591_), .Y(_10592_) );
NOR2X1 NOR2X1_1732 ( .gnd(gnd), .vdd(vdd), .A(_10436_), .B(_10591_), .Y(_10593_) );
NOR2X1 NOR2X1_1733 ( .gnd(gnd), .vdd(vdd), .A(_9324__bF_buf3), .B(_10593_), .Y(_10594_) );
AOI22X1 AOI22X1_77 ( .gnd(gnd), .vdd(vdd), .A(_10592_), .B(_10594_), .C(_10583_), .D(_10590_), .Y(_10595_) );
NOR2X1 NOR2X1_1734 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_89_), .B(_10522__bF_buf4), .Y(_10596_) );
NOR2X1 NOR2X1_1735 ( .gnd(gnd), .vdd(vdd), .A(_9186_), .B(_10519__bF_buf5), .Y(_10597_) );
NOR2X1 NOR2X1_1736 ( .gnd(gnd), .vdd(vdd), .A(_10597_), .B(_10596_), .Y(_10598_) );
AND2X2 AND2X2_699 ( .gnd(gnd), .vdd(vdd), .A(_10598_), .B(_10440_), .Y(_10599_) );
OAI21X1 OAI21X1_2976 ( .gnd(gnd), .vdd(vdd), .A(_10598_), .B(_10440_), .C(micro_hash_ucr_3_pipe30_bF_buf4), .Y(_10600_) );
OAI22X1 OAI22X1_134 ( .gnd(gnd), .vdd(vdd), .A(_10599_), .B(_10600_), .C(_10595_), .D(micro_hash_ucr_3_pipe30_bF_buf3), .Y(_10601_) );
XNOR2X1 XNOR2X1_407 ( .gnd(gnd), .vdd(vdd), .A(_10519__bF_buf4), .B(micro_hash_ucr_3_Wx_97_), .Y(_10602_) );
NOR2X1 NOR2X1_1737 ( .gnd(gnd), .vdd(vdd), .A(_10443_), .B(_10602_), .Y(_10603_) );
NAND2X1 NAND2X1_1402 ( .gnd(gnd), .vdd(vdd), .A(_10443_), .B(_10602_), .Y(_10604_) );
NAND2X1 NAND2X1_1403 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe32_bF_buf2), .B(_10604_), .Y(_10605_) );
OAI21X1 OAI21X1_2977 ( .gnd(gnd), .vdd(vdd), .A(_10605_), .B(_10603_), .C(_9318__bF_buf0), .Y(_10606_) );
AOI21X1 AOI21X1_1854 ( .gnd(gnd), .vdd(vdd), .A(_9317__bF_buf3), .B(_10601_), .C(_10606_), .Y(_10607_) );
AND2X2 AND2X2_700 ( .gnd(gnd), .vdd(vdd), .A(_10386__bF_buf4), .B(micro_hash_ucr_3_Wx_104_), .Y(_10608_) );
NOR2X1 NOR2X1_1738 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_105_), .B(_10522__bF_buf3), .Y(_10609_) );
NOR2X1 NOR2X1_1739 ( .gnd(gnd), .vdd(vdd), .A(_9139_), .B(_10519__bF_buf3), .Y(_10610_) );
NOR2X1 NOR2X1_1740 ( .gnd(gnd), .vdd(vdd), .A(_10610_), .B(_10609_), .Y(_10611_) );
AND2X2 AND2X2_701 ( .gnd(gnd), .vdd(vdd), .A(_10611_), .B(_10608_), .Y(_10612_) );
NOR2X1 NOR2X1_1741 ( .gnd(gnd), .vdd(vdd), .A(_10608_), .B(_10611_), .Y(_10613_) );
OAI21X1 OAI21X1_2978 ( .gnd(gnd), .vdd(vdd), .A(_10612_), .B(_10613_), .C(micro_hash_ucr_3_pipe34_bF_buf3), .Y(_10614_) );
NAND2X1 NAND2X1_1404 ( .gnd(gnd), .vdd(vdd), .A(_9316__bF_buf2), .B(_10614_), .Y(_10615_) );
NOR2X1 NOR2X1_1742 ( .gnd(gnd), .vdd(vdd), .A(_10615_), .B(_10607_), .Y(_10616_) );
XNOR2X1 XNOR2X1_408 ( .gnd(gnd), .vdd(vdd), .A(_10519__bF_buf2), .B(micro_hash_ucr_3_Wx_113_), .Y(_10617_) );
NOR2X1 NOR2X1_1743 ( .gnd(gnd), .vdd(vdd), .A(_10449_), .B(_10617_), .Y(_10618_) );
NAND2X1 NAND2X1_1405 ( .gnd(gnd), .vdd(vdd), .A(_10449_), .B(_10617_), .Y(_10619_) );
NAND2X1 NAND2X1_1406 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe36_bF_buf4), .B(_10619_), .Y(_10620_) );
NOR2X1 NOR2X1_1744 ( .gnd(gnd), .vdd(vdd), .A(_10618_), .B(_10620_), .Y(_10621_) );
OAI21X1 OAI21X1_2979 ( .gnd(gnd), .vdd(vdd), .A(_10616_), .B(_10621_), .C(_9311__bF_buf3), .Y(_10622_) );
OAI21X1 OAI21X1_2980 ( .gnd(gnd), .vdd(vdd), .A(_9311__bF_buf2), .B(_10530_), .C(_10622_), .Y(_10623_) );
XNOR2X1 XNOR2X1_409 ( .gnd(gnd), .vdd(vdd), .A(_10519__bF_buf1), .B(micro_hash_ucr_3_Wx_129_), .Y(_10624_) );
NOR2X1 NOR2X1_1745 ( .gnd(gnd), .vdd(vdd), .A(_10456_), .B(_10624_), .Y(_10625_) );
NAND2X1 NAND2X1_1407 ( .gnd(gnd), .vdd(vdd), .A(_10456_), .B(_10624_), .Y(_10626_) );
NAND2X1 NAND2X1_1408 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe40_bF_buf4), .B(_10626_), .Y(_10627_) );
OAI21X1 OAI21X1_2981 ( .gnd(gnd), .vdd(vdd), .A(_10627_), .B(_10625_), .C(_9310__bF_buf3), .Y(_10628_) );
AOI21X1 AOI21X1_1855 ( .gnd(gnd), .vdd(vdd), .A(_9312__bF_buf2), .B(_10623_), .C(_10628_), .Y(_10629_) );
NOR2X1 NOR2X1_1746 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_137_), .B(_10522__bF_buf2), .Y(_10630_) );
NOR2X1 NOR2X1_1747 ( .gnd(gnd), .vdd(vdd), .A(_9187_), .B(_10519__bF_buf0), .Y(_10631_) );
NOR2X1 NOR2X1_1748 ( .gnd(gnd), .vdd(vdd), .A(_10631_), .B(_10630_), .Y(_10632_) );
AND2X2 AND2X2_702 ( .gnd(gnd), .vdd(vdd), .A(_10632_), .B(_10461_), .Y(_10633_) );
NOR2X1 NOR2X1_1749 ( .gnd(gnd), .vdd(vdd), .A(_10461_), .B(_10632_), .Y(_10634_) );
OAI21X1 OAI21X1_2982 ( .gnd(gnd), .vdd(vdd), .A(_10633_), .B(_10634_), .C(micro_hash_ucr_3_pipe42_bF_buf2), .Y(_10635_) );
NAND2X1 NAND2X1_1409 ( .gnd(gnd), .vdd(vdd), .A(_9305__bF_buf4), .B(_10635_), .Y(_10636_) );
NOR2X1 NOR2X1_1750 ( .gnd(gnd), .vdd(vdd), .A(_10636_), .B(_10629_), .Y(_10637_) );
XNOR2X1 XNOR2X1_410 ( .gnd(gnd), .vdd(vdd), .A(_10519__bF_buf5), .B(micro_hash_ucr_3_Wx_145_), .Y(_10638_) );
NOR2X1 NOR2X1_1751 ( .gnd(gnd), .vdd(vdd), .A(_10465_), .B(_10638_), .Y(_10639_) );
NAND2X1 NAND2X1_1410 ( .gnd(gnd), .vdd(vdd), .A(_10465_), .B(_10638_), .Y(_10640_) );
NAND2X1 NAND2X1_1411 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe44_bF_buf1), .B(_10640_), .Y(_10641_) );
NOR2X1 NOR2X1_1752 ( .gnd(gnd), .vdd(vdd), .A(_10639_), .B(_10641_), .Y(_10642_) );
OAI21X1 OAI21X1_2983 ( .gnd(gnd), .vdd(vdd), .A(_10637_), .B(_10642_), .C(_9306__bF_buf2), .Y(_10643_) );
OAI21X1 OAI21X1_2984 ( .gnd(gnd), .vdd(vdd), .A(_9306__bF_buf1), .B(_10526_), .C(_10643_), .Y(_10644_) );
NOR2X1 NOR2X1_1753 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_161_), .B(_10522__bF_buf1), .Y(_10645_) );
NOR2X1 NOR2X1_1754 ( .gnd(gnd), .vdd(vdd), .A(_8966_), .B(_10519__bF_buf4), .Y(_10646_) );
NOR2X1 NOR2X1_1755 ( .gnd(gnd), .vdd(vdd), .A(_10646_), .B(_10645_), .Y(_10647_) );
NOR2X1 NOR2X1_1756 ( .gnd(gnd), .vdd(vdd), .A(_10472_), .B(_10647_), .Y(_10648_) );
NAND2X1 NAND2X1_1412 ( .gnd(gnd), .vdd(vdd), .A(_10472_), .B(_10647_), .Y(_10649_) );
INVX1 INVX1_651 ( .gnd(gnd), .vdd(vdd), .A(_10649_), .Y(_10650_) );
OAI21X1 OAI21X1_2985 ( .gnd(gnd), .vdd(vdd), .A(_10650_), .B(_10648_), .C(micro_hash_ucr_3_pipe48_bF_buf2), .Y(_10651_) );
OAI21X1 OAI21X1_2986 ( .gnd(gnd), .vdd(vdd), .A(_10644_), .B(micro_hash_ucr_3_pipe48_bF_buf1), .C(_10651_), .Y(_10652_) );
AND2X2 AND2X2_703 ( .gnd(gnd), .vdd(vdd), .A(_10386__bF_buf3), .B(micro_hash_ucr_3_Wx_168_), .Y(_10653_) );
NOR2X1 NOR2X1_1757 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_169_), .B(_10522__bF_buf0), .Y(_10654_) );
NOR2X1 NOR2X1_1758 ( .gnd(gnd), .vdd(vdd), .A(_8836_), .B(_10519__bF_buf3), .Y(_10655_) );
NOR2X1 NOR2X1_1759 ( .gnd(gnd), .vdd(vdd), .A(_10655_), .B(_10654_), .Y(_10656_) );
AND2X2 AND2X2_704 ( .gnd(gnd), .vdd(vdd), .A(_10656_), .B(_10653_), .Y(_10657_) );
NOR2X1 NOR2X1_1760 ( .gnd(gnd), .vdd(vdd), .A(_10653_), .B(_10656_), .Y(_10658_) );
OAI21X1 OAI21X1_2987 ( .gnd(gnd), .vdd(vdd), .A(_10657_), .B(_10658_), .C(micro_hash_ucr_3_pipe50_bF_buf2), .Y(_10659_) );
NAND2X1 NAND2X1_1413 ( .gnd(gnd), .vdd(vdd), .A(_9300__bF_buf1), .B(_10659_), .Y(_10660_) );
AOI21X1 AOI21X1_1856 ( .gnd(gnd), .vdd(vdd), .A(_9299__bF_buf3), .B(_10652_), .C(_10660_), .Y(_10661_) );
XNOR2X1 XNOR2X1_411 ( .gnd(gnd), .vdd(vdd), .A(_10519__bF_buf2), .B(micro_hash_ucr_3_Wx_177_), .Y(_10662_) );
NOR2X1 NOR2X1_1761 ( .gnd(gnd), .vdd(vdd), .A(_10478_), .B(_10662_), .Y(_10663_) );
NAND2X1 NAND2X1_1414 ( .gnd(gnd), .vdd(vdd), .A(_10478_), .B(_10662_), .Y(_10664_) );
NAND2X1 NAND2X1_1415 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe52_bF_buf4), .B(_10664_), .Y(_10665_) );
OAI21X1 OAI21X1_2988 ( .gnd(gnd), .vdd(vdd), .A(_10665_), .B(_10663_), .C(_9298__bF_buf3), .Y(_10666_) );
XNOR2X1 XNOR2X1_412 ( .gnd(gnd), .vdd(vdd), .A(_10519__bF_buf1), .B(micro_hash_ucr_3_Wx_185_), .Y(_10667_) );
XOR2X1 XOR2X1_170 ( .gnd(gnd), .vdd(vdd), .A(_10667_), .B(_10482_), .Y(_10668_) );
OAI22X1 OAI22X1_135 ( .gnd(gnd), .vdd(vdd), .A(_9298__bF_buf2), .B(_10668_), .C(_10661_), .D(_10666_), .Y(_10669_) );
NOR2X1 NOR2X1_1762 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_193_), .B(_10522__bF_buf4), .Y(_10670_) );
NOR2X1 NOR2X1_1763 ( .gnd(gnd), .vdd(vdd), .A(_8937_), .B(_10519__bF_buf0), .Y(_10671_) );
NOR2X1 NOR2X1_1764 ( .gnd(gnd), .vdd(vdd), .A(_10671_), .B(_10670_), .Y(_10672_) );
NOR2X1 NOR2X1_1765 ( .gnd(gnd), .vdd(vdd), .A(_10486_), .B(_10672_), .Y(_10673_) );
NAND2X1 NAND2X1_1416 ( .gnd(gnd), .vdd(vdd), .A(_10486_), .B(_10672_), .Y(_10674_) );
INVX1 INVX1_652 ( .gnd(gnd), .vdd(vdd), .A(_10674_), .Y(_10675_) );
NOR2X1 NOR2X1_1766 ( .gnd(gnd), .vdd(vdd), .A(_10673_), .B(_10675_), .Y(_10676_) );
AOI21X1 AOI21X1_1857 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe56_bF_buf3), .B(_10676_), .C(micro_hash_ucr_3_pipe58_bF_buf2), .Y(_10677_) );
OAI21X1 OAI21X1_2989 ( .gnd(gnd), .vdd(vdd), .A(_10669_), .B(micro_hash_ucr_3_pipe56_bF_buf2), .C(_10677_), .Y(_10678_) );
NAND2X1 NAND2X1_1417 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_200_), .B(_10386__bF_buf2), .Y(_10679_) );
NOR2X1 NOR2X1_1767 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_201_), .B(_10522__bF_buf3), .Y(_10680_) );
NAND2X1 NAND2X1_1418 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_201_), .B(_10522__bF_buf2), .Y(_10681_) );
INVX1 INVX1_653 ( .gnd(gnd), .vdd(vdd), .A(_10681_), .Y(_10682_) );
NOR2X1 NOR2X1_1768 ( .gnd(gnd), .vdd(vdd), .A(_10680_), .B(_10682_), .Y(_10683_) );
INVX1 INVX1_654 ( .gnd(gnd), .vdd(vdd), .A(_10683_), .Y(_10684_) );
NOR2X1 NOR2X1_1769 ( .gnd(gnd), .vdd(vdd), .A(_10679_), .B(_10684_), .Y(_10685_) );
AOI21X1 AOI21X1_1858 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_200_), .B(_10386__bF_buf1), .C(_10683_), .Y(_10686_) );
OAI21X1 OAI21X1_2990 ( .gnd(gnd), .vdd(vdd), .A(_10685_), .B(_10686_), .C(micro_hash_ucr_3_pipe58_bF_buf1), .Y(_10687_) );
NAND3X1 NAND3X1_580 ( .gnd(gnd), .vdd(vdd), .A(_9292__bF_buf3), .B(_10687_), .C(_10678_), .Y(_10688_) );
NOR2X1 NOR2X1_1770 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_209_), .B(_10522__bF_buf1), .Y(_10689_) );
NOR2X1 NOR2X1_1771 ( .gnd(gnd), .vdd(vdd), .A(_8967_), .B(_10519__bF_buf5), .Y(_10690_) );
NOR2X1 NOR2X1_1772 ( .gnd(gnd), .vdd(vdd), .A(_10690_), .B(_10689_), .Y(_10691_) );
NAND2X1 NAND2X1_1419 ( .gnd(gnd), .vdd(vdd), .A(_10492_), .B(_10691_), .Y(_10692_) );
INVX1 INVX1_655 ( .gnd(gnd), .vdd(vdd), .A(_10692_), .Y(_10693_) );
OAI21X1 OAI21X1_2991 ( .gnd(gnd), .vdd(vdd), .A(_10691_), .B(_10492_), .C(micro_hash_ucr_3_pipe60_bF_buf2), .Y(_10694_) );
OAI21X1 OAI21X1_2992 ( .gnd(gnd), .vdd(vdd), .A(_10693_), .B(_10694_), .C(_10688_), .Y(_10695_) );
NAND2X1 NAND2X1_1420 ( .gnd(gnd), .vdd(vdd), .A(_9287__bF_buf3), .B(_10695_), .Y(_10696_) );
OAI21X1 OAI21X1_2993 ( .gnd(gnd), .vdd(vdd), .A(_9287__bF_buf2), .B(_10521_), .C(_10696_), .Y(_10697_) );
NOR2X1 NOR2X1_1773 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_225_), .B(_10522__bF_buf0), .Y(_10698_) );
INVX2 INVX2_368 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_225_), .Y(_10699_) );
NOR2X1 NOR2X1_1774 ( .gnd(gnd), .vdd(vdd), .A(_10699_), .B(_10519__bF_buf4), .Y(_10700_) );
NOR2X1 NOR2X1_1775 ( .gnd(gnd), .vdd(vdd), .A(_10700_), .B(_10698_), .Y(_10701_) );
NAND2X1 NAND2X1_1421 ( .gnd(gnd), .vdd(vdd), .A(_10500_), .B(_10701_), .Y(_10702_) );
INVX1 INVX1_656 ( .gnd(gnd), .vdd(vdd), .A(_10702_), .Y(_10703_) );
NOR2X1 NOR2X1_1776 ( .gnd(gnd), .vdd(vdd), .A(_10500_), .B(_10701_), .Y(_10704_) );
OAI21X1 OAI21X1_2994 ( .gnd(gnd), .vdd(vdd), .A(_10703_), .B(_10704_), .C(micro_hash_ucr_3_pipe64_bF_buf3), .Y(_10705_) );
OAI21X1 OAI21X1_2995 ( .gnd(gnd), .vdd(vdd), .A(_10697_), .B(micro_hash_ucr_3_pipe64_bF_buf2), .C(_10705_), .Y(_10706_) );
NOR2X1 NOR2X1_1777 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_233_), .B(_10522__bF_buf4), .Y(_10707_) );
AND2X2 AND2X2_705 ( .gnd(gnd), .vdd(vdd), .A(_10522__bF_buf3), .B(micro_hash_ucr_3_Wx_233_), .Y(_10708_) );
NOR2X1 NOR2X1_1778 ( .gnd(gnd), .vdd(vdd), .A(_10707_), .B(_10708_), .Y(_10709_) );
AND2X2 AND2X2_706 ( .gnd(gnd), .vdd(vdd), .A(_10709_), .B(_10388_), .Y(_10710_) );
OAI21X1 OAI21X1_2996 ( .gnd(gnd), .vdd(vdd), .A(_10709_), .B(_10388_), .C(micro_hash_ucr_3_pipe66_bF_buf4), .Y(_10711_) );
OAI22X1 OAI22X1_136 ( .gnd(gnd), .vdd(vdd), .A(_10710_), .B(_10711_), .C(_10706_), .D(micro_hash_ucr_3_pipe66_bF_buf3), .Y(_10712_) );
XNOR2X1 XNOR2X1_413 ( .gnd(gnd), .vdd(vdd), .A(_10519__bF_buf3), .B(micro_hash_ucr_3_Wx_241_), .Y(_10713_) );
NOR2X1 NOR2X1_1779 ( .gnd(gnd), .vdd(vdd), .A(_10506_), .B(_10713_), .Y(_10714_) );
NAND2X1 NAND2X1_1422 ( .gnd(gnd), .vdd(vdd), .A(_10506_), .B(_10713_), .Y(_10715_) );
NAND2X1 NAND2X1_1423 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe68_bF_buf1), .B(_10715_), .Y(_10716_) );
OAI21X1 OAI21X1_2997 ( .gnd(gnd), .vdd(vdd), .A(_10716_), .B(_10714_), .C(_9283__bF_buf3), .Y(_10717_) );
AOI21X1 AOI21X1_1859 ( .gnd(gnd), .vdd(vdd), .A(_9282__bF_buf3), .B(_10712_), .C(_10717_), .Y(_10718_) );
NOR2X1 NOR2X1_1780 ( .gnd(gnd), .vdd(vdd), .A(_10509_), .B(_10387__bF_buf0), .Y(_10719_) );
NOR2X1 NOR2X1_1781 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_249_), .B(_10522__bF_buf2), .Y(_10720_) );
INVX1 INVX1_657 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_249_), .Y(_10721_) );
NOR2X1 NOR2X1_1782 ( .gnd(gnd), .vdd(vdd), .A(_10721_), .B(_10519__bF_buf2), .Y(_10722_) );
NOR2X1 NOR2X1_1783 ( .gnd(gnd), .vdd(vdd), .A(_10722_), .B(_10720_), .Y(_10723_) );
AOI21X1 AOI21X1_1860 ( .gnd(gnd), .vdd(vdd), .A(_10719_), .B(_10723_), .C(_8800__bF_buf4), .Y(_10724_) );
OAI21X1 OAI21X1_2998 ( .gnd(gnd), .vdd(vdd), .A(_10719_), .B(_10723_), .C(_10724_), .Y(_10725_) );
AOI21X1 AOI21X1_1861 ( .gnd(gnd), .vdd(vdd), .A(_10381_), .B(_10725_), .C(_10718_), .Y(_8702__1_) );
INVX1 INVX1_658 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_17_), .Y(_10726_) );
NAND2X1 NAND2X1_1424 ( .gnd(gnd), .vdd(vdd), .A(_10543_), .B(_10544_), .Y(_10727_) );
OAI21X1 OAI21X1_2999 ( .gnd(gnd), .vdd(vdd), .A(_10726_), .B(_10519__bF_buf1), .C(_10727_), .Y(_10728_) );
OAI21X1 OAI21X1_3000 ( .gnd(gnd), .vdd(vdd), .A(_10513_), .B(_10514_), .C(_10517_), .Y(_10729_) );
INVX1 INVX1_659 ( .gnd(gnd), .vdd(vdd), .A(_10729_), .Y(_10730_) );
INVX1 INVX1_660 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_k_2_), .Y(_10731_) );
INVX1 INVX1_661 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_x_2_), .Y(_10732_) );
NAND2X1 NAND2X1_1425 ( .gnd(gnd), .vdd(vdd), .A(_10731_), .B(_10732_), .Y(_10733_) );
NOR2X1 NOR2X1_1784 ( .gnd(gnd), .vdd(vdd), .A(_10731_), .B(_10732_), .Y(_10734_) );
INVX2 INVX2_369 ( .gnd(gnd), .vdd(vdd), .A(_10734_), .Y(_10735_) );
NAND2X1 NAND2X1_1426 ( .gnd(gnd), .vdd(vdd), .A(_10733_), .B(_10735_), .Y(_10736_) );
NOR2X1 NOR2X1_1785 ( .gnd(gnd), .vdd(vdd), .A(_10736_), .B(_10730_), .Y(_10737_) );
AOI21X1 AOI21X1_1862 ( .gnd(gnd), .vdd(vdd), .A(_10733_), .B(_10735_), .C(_10729_), .Y(_10738_) );
NOR2X1 NOR2X1_1786 ( .gnd(gnd), .vdd(vdd), .A(_10738__bF_buf3), .B(_10737__bF_buf3), .Y(_10739_) );
NOR2X1 NOR2X1_1787 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_18_), .B(_10739__bF_buf3), .Y(_10740_) );
AND2X2 AND2X2_707 ( .gnd(gnd), .vdd(vdd), .A(_10739__bF_buf2), .B(micro_hash_ucr_3_Wx_18_), .Y(_10741_) );
NOR2X1 NOR2X1_1788 ( .gnd(gnd), .vdd(vdd), .A(_10740_), .B(_10741_), .Y(_10742_) );
XNOR2X1 XNOR2X1_414 ( .gnd(gnd), .vdd(vdd), .A(_10742_), .B(_10728_), .Y(_10743_) );
OAI21X1 OAI21X1_3001 ( .gnd(gnd), .vdd(vdd), .A(_10531_), .B(_10519__bF_buf0), .C(_10533_), .Y(_10744_) );
INVX2 INVX2_370 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_10_), .Y(_10745_) );
XNOR2X1 XNOR2X1_415 ( .gnd(gnd), .vdd(vdd), .A(_10739__bF_buf1), .B(_10745_), .Y(_10746_) );
NAND2X1 NAND2X1_1427 ( .gnd(gnd), .vdd(vdd), .A(_10744_), .B(_10746_), .Y(_10747_) );
INVX1 INVX1_662 ( .gnd(gnd), .vdd(vdd), .A(_10747_), .Y(_10748_) );
OAI21X1 OAI21X1_3002 ( .gnd(gnd), .vdd(vdd), .A(_10746_), .B(_10744_), .C(micro_hash_ucr_3_pipe10_bF_buf3), .Y(_10749_) );
AOI21X1 AOI21X1_1863 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_1_), .B(_10522__bF_buf1), .C(_10537_), .Y(_10750_) );
XNOR2X1 XNOR2X1_416 ( .gnd(gnd), .vdd(vdd), .A(_10739__bF_buf0), .B(micro_hash_ucr_3_Wx_2_), .Y(_10751_) );
NAND2X1 NAND2X1_1428 ( .gnd(gnd), .vdd(vdd), .A(_10750_), .B(_10751_), .Y(_10752_) );
NOR2X1 NOR2X1_1789 ( .gnd(gnd), .vdd(vdd), .A(_10750_), .B(_10751_), .Y(_10753_) );
INVX1 INVX1_663 ( .gnd(gnd), .vdd(vdd), .A(_10753_), .Y(_10754_) );
AOI21X1 AOI21X1_1864 ( .gnd(gnd), .vdd(vdd), .A(_10752_), .B(_10754_), .C(_9341_), .Y(_10755_) );
NAND2X1 NAND2X1_1429 ( .gnd(gnd), .vdd(vdd), .A(H_3_18_), .B(micro_hash_ucr_3_pipe6_bF_buf1), .Y(_10756_) );
OAI21X1 OAI21X1_3003 ( .gnd(gnd), .vdd(vdd), .A(_9593__bF_buf2), .B(micro_hash_ucr_3_pipe6_bF_buf0), .C(_10756_), .Y(_10757_) );
OAI21X1 OAI21X1_3004 ( .gnd(gnd), .vdd(vdd), .A(_10757_), .B(micro_hash_ucr_3_pipe8), .C(_9342_), .Y(_10758_) );
OAI22X1 OAI22X1_137 ( .gnd(gnd), .vdd(vdd), .A(_10748_), .B(_10749_), .C(_10755_), .D(_10758_), .Y(_10759_) );
NAND2X1 NAND2X1_1430 ( .gnd(gnd), .vdd(vdd), .A(_9340_), .B(_10759_), .Y(_10760_) );
OAI21X1 OAI21X1_3005 ( .gnd(gnd), .vdd(vdd), .A(_9340_), .B(_10743_), .C(_10760_), .Y(_10761_) );
NAND2X1 NAND2X1_1431 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_25_), .B(_10522__bF_buf0), .Y(_10762_) );
OAI21X1 OAI21X1_3006 ( .gnd(gnd), .vdd(vdd), .A(_10548_), .B(_10547_), .C(_10762_), .Y(_10763_) );
INVX2 INVX2_371 ( .gnd(gnd), .vdd(vdd), .A(_10763_), .Y(_10764_) );
XNOR2X1 XNOR2X1_417 ( .gnd(gnd), .vdd(vdd), .A(_10739__bF_buf3), .B(micro_hash_ucr_3_Wx_26_), .Y(_10765_) );
NOR2X1 NOR2X1_1790 ( .gnd(gnd), .vdd(vdd), .A(_10764_), .B(_10765_), .Y(_10766_) );
AND2X2 AND2X2_708 ( .gnd(gnd), .vdd(vdd), .A(_10764_), .B(_10765_), .Y(_10767_) );
OAI21X1 OAI21X1_3007 ( .gnd(gnd), .vdd(vdd), .A(_10766_), .B(_10767_), .C(micro_hash_ucr_3_pipe14_bF_buf2), .Y(_10768_) );
OAI21X1 OAI21X1_3008 ( .gnd(gnd), .vdd(vdd), .A(_10761_), .B(micro_hash_ucr_3_pipe14_bF_buf1), .C(_10768_), .Y(_10769_) );
OAI21X1 OAI21X1_3009 ( .gnd(gnd), .vdd(vdd), .A(_10554_), .B(_10553_), .C(_10555_), .Y(_10770_) );
INVX2 INVX2_372 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_34_), .Y(_10771_) );
XNOR2X1 XNOR2X1_418 ( .gnd(gnd), .vdd(vdd), .A(_10739__bF_buf2), .B(_10771_), .Y(_10772_) );
NOR2X1 NOR2X1_1791 ( .gnd(gnd), .vdd(vdd), .A(_10770_), .B(_10772_), .Y(_10773_) );
NAND2X1 NAND2X1_1432 ( .gnd(gnd), .vdd(vdd), .A(_10770_), .B(_10772_), .Y(_10774_) );
NAND2X1 NAND2X1_1433 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe16_bF_buf1), .B(_10774_), .Y(_10775_) );
OAI22X1 OAI22X1_138 ( .gnd(gnd), .vdd(vdd), .A(_10773_), .B(_10775_), .C(_10769_), .D(micro_hash_ucr_3_pipe16_bF_buf0), .Y(_10776_) );
INVX1 INVX1_664 ( .gnd(gnd), .vdd(vdd), .A(_10416_), .Y(_10777_) );
OAI21X1 OAI21X1_3010 ( .gnd(gnd), .vdd(vdd), .A(_10567_), .B(_10777_), .C(_10568_), .Y(_10778_) );
INVX2 INVX2_373 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_42_), .Y(_10779_) );
XNOR2X1 XNOR2X1_419 ( .gnd(gnd), .vdd(vdd), .A(_10739__bF_buf1), .B(_10779_), .Y(_10780_) );
NOR2X1 NOR2X1_1792 ( .gnd(gnd), .vdd(vdd), .A(_10778_), .B(_10780_), .Y(_10781_) );
NAND2X1 NAND2X1_1434 ( .gnd(gnd), .vdd(vdd), .A(_10778_), .B(_10780_), .Y(_10782_) );
INVX1 INVX1_665 ( .gnd(gnd), .vdd(vdd), .A(_10782_), .Y(_10783_) );
OAI21X1 OAI21X1_3011 ( .gnd(gnd), .vdd(vdd), .A(_10783_), .B(_10781_), .C(micro_hash_ucr_3_pipe18_bF_buf2), .Y(_10784_) );
OAI21X1 OAI21X1_3012 ( .gnd(gnd), .vdd(vdd), .A(_10776_), .B(micro_hash_ucr_3_pipe18_bF_buf1), .C(_10784_), .Y(_10785_) );
OAI21X1 OAI21X1_3013 ( .gnd(gnd), .vdd(vdd), .A(_10562_), .B(_10561_), .C(_10563_), .Y(_10786_) );
INVX2 INVX2_374 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_50_), .Y(_10787_) );
XNOR2X1 XNOR2X1_420 ( .gnd(gnd), .vdd(vdd), .A(_10739__bF_buf0), .B(_10787_), .Y(_10788_) );
NOR2X1 NOR2X1_1793 ( .gnd(gnd), .vdd(vdd), .A(_10786_), .B(_10788_), .Y(_10789_) );
NAND2X1 NAND2X1_1435 ( .gnd(gnd), .vdd(vdd), .A(_10786_), .B(_10788_), .Y(_10790_) );
INVX1 INVX1_666 ( .gnd(gnd), .vdd(vdd), .A(_10790_), .Y(_10791_) );
OAI21X1 OAI21X1_3014 ( .gnd(gnd), .vdd(vdd), .A(_10791_), .B(_10789_), .C(micro_hash_ucr_3_pipe20_bF_buf0), .Y(_10792_) );
NAND2X1 NAND2X1_1436 ( .gnd(gnd), .vdd(vdd), .A(_9330__bF_buf4), .B(_10792_), .Y(_10793_) );
AOI21X1 AOI21X1_1865 ( .gnd(gnd), .vdd(vdd), .A(_9329__bF_buf0), .B(_10785_), .C(_10793_), .Y(_10794_) );
AOI21X1 AOI21X1_1866 ( .gnd(gnd), .vdd(vdd), .A(_10424_), .B(_10577_), .C(_10576_), .Y(_10795_) );
OAI21X1 OAI21X1_3015 ( .gnd(gnd), .vdd(vdd), .A(_10737__bF_buf2), .B(_10738__bF_buf2), .C(_9266_), .Y(_10796_) );
INVX1 INVX1_667 ( .gnd(gnd), .vdd(vdd), .A(_10796_), .Y(_10797_) );
INVX8 INVX8_279 ( .gnd(gnd), .vdd(vdd), .A(_10739__bF_buf3), .Y(_10798_) );
NOR2X1 NOR2X1_1794 ( .gnd(gnd), .vdd(vdd), .A(_9266_), .B(_10798__bF_buf5), .Y(_10799_) );
NOR3X1 NOR3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_10799_), .B(_10797_), .C(_10795_), .Y(_10800_) );
OAI21X1 OAI21X1_3016 ( .gnd(gnd), .vdd(vdd), .A(_10799_), .B(_10797_), .C(_10795_), .Y(_10801_) );
NAND2X1 NAND2X1_1437 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe22_bF_buf1), .B(_10801_), .Y(_10802_) );
OAI21X1 OAI21X1_3017 ( .gnd(gnd), .vdd(vdd), .A(_10802_), .B(_10800_), .C(_9328__bF_buf1), .Y(_10803_) );
NAND2X1 NAND2X1_1438 ( .gnd(gnd), .vdd(vdd), .A(_10427_), .B(_10580_), .Y(_10804_) );
OAI21X1 OAI21X1_3018 ( .gnd(gnd), .vdd(vdd), .A(_9240_), .B(_10519__bF_buf5), .C(_10804_), .Y(_10805_) );
OAI21X1 OAI21X1_3019 ( .gnd(gnd), .vdd(vdd), .A(_10737__bF_buf1), .B(_10738__bF_buf1), .C(_9243_), .Y(_10806_) );
NOR2X1 NOR2X1_1795 ( .gnd(gnd), .vdd(vdd), .A(_9243_), .B(_10798__bF_buf4), .Y(_10807_) );
INVX1 INVX1_668 ( .gnd(gnd), .vdd(vdd), .A(_10807_), .Y(_10808_) );
NAND2X1 NAND2X1_1439 ( .gnd(gnd), .vdd(vdd), .A(_10806_), .B(_10808_), .Y(_10809_) );
XOR2X1 XOR2X1_171 ( .gnd(gnd), .vdd(vdd), .A(_10809_), .B(_10805_), .Y(_10810_) );
AOI21X1 AOI21X1_1867 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe24_bF_buf1), .B(_10810_), .C(micro_hash_ucr_3_pipe26_bF_buf0), .Y(_10811_) );
OAI21X1 OAI21X1_3020 ( .gnd(gnd), .vdd(vdd), .A(_10794_), .B(_10803_), .C(_10811_), .Y(_10812_) );
OAI21X1 OAI21X1_3021 ( .gnd(gnd), .vdd(vdd), .A(_9162_), .B(_10519__bF_buf4), .C(_10587_), .Y(_10813_) );
XNOR2X1 XNOR2X1_421 ( .gnd(gnd), .vdd(vdd), .A(_10739__bF_buf2), .B(_9165_), .Y(_10814_) );
NAND2X1 NAND2X1_1440 ( .gnd(gnd), .vdd(vdd), .A(_10814_), .B(_10813_), .Y(_10815_) );
INVX1 INVX1_669 ( .gnd(gnd), .vdd(vdd), .A(_10815_), .Y(_10816_) );
OAI21X1 OAI21X1_3022 ( .gnd(gnd), .vdd(vdd), .A(_10813_), .B(_10814_), .C(micro_hash_ucr_3_pipe26_bF_buf4), .Y(_10817_) );
OAI21X1 OAI21X1_3023 ( .gnd(gnd), .vdd(vdd), .A(_10816_), .B(_10817_), .C(_10812_), .Y(_10818_) );
OAI21X1 OAI21X1_3024 ( .gnd(gnd), .vdd(vdd), .A(_9217_), .B(_10519__bF_buf3), .C(_10592_), .Y(_10819_) );
OAI21X1 OAI21X1_3025 ( .gnd(gnd), .vdd(vdd), .A(_10737__bF_buf0), .B(_10738__bF_buf0), .C(_9220_), .Y(_10820_) );
NOR2X1 NOR2X1_1796 ( .gnd(gnd), .vdd(vdd), .A(_9220_), .B(_10798__bF_buf3), .Y(_10821_) );
INVX1 INVX1_670 ( .gnd(gnd), .vdd(vdd), .A(_10821_), .Y(_10822_) );
NAND2X1 NAND2X1_1441 ( .gnd(gnd), .vdd(vdd), .A(_10820_), .B(_10822_), .Y(_10823_) );
XOR2X1 XOR2X1_172 ( .gnd(gnd), .vdd(vdd), .A(_10823_), .B(_10819_), .Y(_10824_) );
AOI21X1 AOI21X1_1868 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe28_bF_buf4), .B(_10824_), .C(micro_hash_ucr_3_pipe30_bF_buf2), .Y(_10825_) );
OAI21X1 OAI21X1_3026 ( .gnd(gnd), .vdd(vdd), .A(_10818_), .B(micro_hash_ucr_3_pipe28_bF_buf3), .C(_10825_), .Y(_10826_) );
OAI21X1 OAI21X1_3027 ( .gnd(gnd), .vdd(vdd), .A(_10737__bF_buf3), .B(_10738__bF_buf3), .C(_9190_), .Y(_10827_) );
INVX1 INVX1_671 ( .gnd(gnd), .vdd(vdd), .A(_10827_), .Y(_10828_) );
NOR2X1 NOR2X1_1797 ( .gnd(gnd), .vdd(vdd), .A(_9190_), .B(_10798__bF_buf2), .Y(_10829_) );
NOR2X1 NOR2X1_1798 ( .gnd(gnd), .vdd(vdd), .A(_10828_), .B(_10829_), .Y(_10830_) );
OAI21X1 OAI21X1_3028 ( .gnd(gnd), .vdd(vdd), .A(_10597_), .B(_10599_), .C(_10830_), .Y(_10831_) );
NOR2X1 NOR2X1_1799 ( .gnd(gnd), .vdd(vdd), .A(_10597_), .B(_10599_), .Y(_10832_) );
OAI21X1 OAI21X1_3029 ( .gnd(gnd), .vdd(vdd), .A(_10828_), .B(_10829_), .C(_10832_), .Y(_10833_) );
NAND2X1 NAND2X1_1442 ( .gnd(gnd), .vdd(vdd), .A(_10833_), .B(_10831_), .Y(_10834_) );
OAI21X1 OAI21X1_3030 ( .gnd(gnd), .vdd(vdd), .A(_9322__bF_buf2), .B(_10834_), .C(_10826_), .Y(_10835_) );
OAI21X1 OAI21X1_3031 ( .gnd(gnd), .vdd(vdd), .A(_9043_), .B(_10519__bF_buf2), .C(_10604_), .Y(_10836_) );
OAI21X1 OAI21X1_3032 ( .gnd(gnd), .vdd(vdd), .A(_10737__bF_buf2), .B(_10738__bF_buf2), .C(_9047_), .Y(_10837_) );
NOR2X1 NOR2X1_1800 ( .gnd(gnd), .vdd(vdd), .A(_9047_), .B(_10798__bF_buf1), .Y(_10838_) );
INVX1 INVX1_672 ( .gnd(gnd), .vdd(vdd), .A(_10838_), .Y(_10839_) );
NAND2X1 NAND2X1_1443 ( .gnd(gnd), .vdd(vdd), .A(_10837_), .B(_10839_), .Y(_10840_) );
XNOR2X1 XNOR2X1_422 ( .gnd(gnd), .vdd(vdd), .A(_10840_), .B(_10836_), .Y(_10841_) );
MUX2X1 MUX2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_10835_), .B(_10841_), .S(_9317__bF_buf2), .Y(_10842_) );
NOR2X1 NOR2X1_1801 ( .gnd(gnd), .vdd(vdd), .A(_10610_), .B(_10612_), .Y(_10843_) );
OAI21X1 OAI21X1_3033 ( .gnd(gnd), .vdd(vdd), .A(_10737__bF_buf1), .B(_10738__bF_buf1), .C(_9142_), .Y(_10844_) );
INVX1 INVX1_673 ( .gnd(gnd), .vdd(vdd), .A(_10844_), .Y(_10845_) );
NOR2X1 NOR2X1_1802 ( .gnd(gnd), .vdd(vdd), .A(_9142_), .B(_10798__bF_buf0), .Y(_10846_) );
OAI21X1 OAI21X1_3034 ( .gnd(gnd), .vdd(vdd), .A(_10845_), .B(_10846_), .C(_10843_), .Y(_10847_) );
NOR2X1 NOR2X1_1803 ( .gnd(gnd), .vdd(vdd), .A(_10845_), .B(_10846_), .Y(_10848_) );
OAI21X1 OAI21X1_3035 ( .gnd(gnd), .vdd(vdd), .A(_10610_), .B(_10612_), .C(_10848_), .Y(_10849_) );
AOI21X1 AOI21X1_1869 ( .gnd(gnd), .vdd(vdd), .A(_10847_), .B(_10849_), .C(_9318__bF_buf4), .Y(_10850_) );
AOI21X1 AOI21X1_1870 ( .gnd(gnd), .vdd(vdd), .A(_9318__bF_buf3), .B(_10842_), .C(_10850_), .Y(_10851_) );
OAI21X1 OAI21X1_3036 ( .gnd(gnd), .vdd(vdd), .A(_9117_), .B(_10519__bF_buf1), .C(_10619_), .Y(_10852_) );
OAI21X1 OAI21X1_3037 ( .gnd(gnd), .vdd(vdd), .A(_10737__bF_buf0), .B(_10738__bF_buf0), .C(_9120_), .Y(_10853_) );
NOR2X1 NOR2X1_1804 ( .gnd(gnd), .vdd(vdd), .A(_9120_), .B(_10798__bF_buf5), .Y(_10854_) );
INVX1 INVX1_674 ( .gnd(gnd), .vdd(vdd), .A(_10854_), .Y(_10855_) );
NAND2X1 NAND2X1_1444 ( .gnd(gnd), .vdd(vdd), .A(_10853_), .B(_10855_), .Y(_10856_) );
XOR2X1 XOR2X1_173 ( .gnd(gnd), .vdd(vdd), .A(_10856_), .B(_10852_), .Y(_10857_) );
AOI21X1 AOI21X1_1871 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe36_bF_buf3), .B(_10857_), .C(micro_hash_ucr_3_pipe38_bF_buf2), .Y(_10858_) );
OAI21X1 OAI21X1_3038 ( .gnd(gnd), .vdd(vdd), .A(_10851_), .B(micro_hash_ucr_3_pipe36_bF_buf2), .C(_10858_), .Y(_10859_) );
AOI21X1 AOI21X1_1872 ( .gnd(gnd), .vdd(vdd), .A(_10453_), .B(_10529_), .C(_10528_), .Y(_10860_) );
OAI21X1 OAI21X1_3039 ( .gnd(gnd), .vdd(vdd), .A(_10737__bF_buf3), .B(_10738__bF_buf3), .C(_9024_), .Y(_10861_) );
INVX1 INVX1_675 ( .gnd(gnd), .vdd(vdd), .A(_10861_), .Y(_10862_) );
NOR2X1 NOR2X1_1805 ( .gnd(gnd), .vdd(vdd), .A(_9024_), .B(_10798__bF_buf4), .Y(_10863_) );
NOR2X1 NOR2X1_1806 ( .gnd(gnd), .vdd(vdd), .A(_10862_), .B(_10863_), .Y(_10864_) );
INVX1 INVX1_676 ( .gnd(gnd), .vdd(vdd), .A(_10864_), .Y(_10865_) );
NOR2X1 NOR2X1_1807 ( .gnd(gnd), .vdd(vdd), .A(_10860_), .B(_10865_), .Y(_10866_) );
INVX1 INVX1_677 ( .gnd(gnd), .vdd(vdd), .A(_10866_), .Y(_10867_) );
OAI21X1 OAI21X1_3040 ( .gnd(gnd), .vdd(vdd), .A(_10863_), .B(_10862_), .C(_10860_), .Y(_10868_) );
NAND2X1 NAND2X1_1445 ( .gnd(gnd), .vdd(vdd), .A(_10868_), .B(_10867_), .Y(_10869_) );
OAI21X1 OAI21X1_3041 ( .gnd(gnd), .vdd(vdd), .A(_9311__bF_buf1), .B(_10869_), .C(_10859_), .Y(_10870_) );
NOR2X1 NOR2X1_1808 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe40_bF_buf3), .B(_10870_), .Y(_10871_) );
OAI21X1 OAI21X1_3042 ( .gnd(gnd), .vdd(vdd), .A(_9072_), .B(_10519__bF_buf0), .C(_10626_), .Y(_10872_) );
OAI21X1 OAI21X1_3043 ( .gnd(gnd), .vdd(vdd), .A(_10737__bF_buf2), .B(_10738__bF_buf2), .C(_9076_), .Y(_10873_) );
NOR2X1 NOR2X1_1809 ( .gnd(gnd), .vdd(vdd), .A(_9076_), .B(_10798__bF_buf3), .Y(_10874_) );
INVX1 INVX1_678 ( .gnd(gnd), .vdd(vdd), .A(_10874_), .Y(_10875_) );
NAND2X1 NAND2X1_1446 ( .gnd(gnd), .vdd(vdd), .A(_10873_), .B(_10875_), .Y(_10876_) );
XNOR2X1 XNOR2X1_423 ( .gnd(gnd), .vdd(vdd), .A(_10876_), .B(_10872_), .Y(_10877_) );
OAI21X1 OAI21X1_3044 ( .gnd(gnd), .vdd(vdd), .A(_10877_), .B(_9312__bF_buf1), .C(_9310__bF_buf2), .Y(_10878_) );
NOR2X1 NOR2X1_1810 ( .gnd(gnd), .vdd(vdd), .A(_10631_), .B(_10633_), .Y(_10879_) );
OAI21X1 OAI21X1_3045 ( .gnd(gnd), .vdd(vdd), .A(_10737__bF_buf1), .B(_10738__bF_buf1), .C(_9191_), .Y(_10880_) );
INVX1 INVX1_679 ( .gnd(gnd), .vdd(vdd), .A(_10880_), .Y(_10881_) );
NOR2X1 NOR2X1_1811 ( .gnd(gnd), .vdd(vdd), .A(_9191_), .B(_10798__bF_buf2), .Y(_10882_) );
OAI21X1 OAI21X1_3046 ( .gnd(gnd), .vdd(vdd), .A(_10881_), .B(_10882_), .C(_10879_), .Y(_10883_) );
NOR2X1 NOR2X1_1812 ( .gnd(gnd), .vdd(vdd), .A(_10881_), .B(_10882_), .Y(_10884_) );
OAI21X1 OAI21X1_3047 ( .gnd(gnd), .vdd(vdd), .A(_10631_), .B(_10633_), .C(_10884_), .Y(_10885_) );
AND2X2 AND2X2_709 ( .gnd(gnd), .vdd(vdd), .A(_10885_), .B(micro_hash_ucr_3_pipe42_bF_buf1), .Y(_10886_) );
AOI21X1 AOI21X1_1873 ( .gnd(gnd), .vdd(vdd), .A(_10883_), .B(_10886_), .C(micro_hash_ucr_3_pipe44_bF_buf0), .Y(_10887_) );
OAI21X1 OAI21X1_3048 ( .gnd(gnd), .vdd(vdd), .A(_10871_), .B(_10878_), .C(_10887_), .Y(_10888_) );
OAI21X1 OAI21X1_3049 ( .gnd(gnd), .vdd(vdd), .A(_8936_), .B(_10519__bF_buf5), .C(_10640_), .Y(_10889_) );
OAI21X1 OAI21X1_3050 ( .gnd(gnd), .vdd(vdd), .A(_10737__bF_buf0), .B(_10738__bF_buf0), .C(_8940_), .Y(_10890_) );
NOR2X1 NOR2X1_1813 ( .gnd(gnd), .vdd(vdd), .A(_8940_), .B(_10798__bF_buf1), .Y(_10891_) );
INVX1 INVX1_680 ( .gnd(gnd), .vdd(vdd), .A(_10891_), .Y(_10892_) );
NAND2X1 NAND2X1_1447 ( .gnd(gnd), .vdd(vdd), .A(_10890_), .B(_10892_), .Y(_10893_) );
XOR2X1 XOR2X1_174 ( .gnd(gnd), .vdd(vdd), .A(_10893_), .B(_10889_), .Y(_10894_) );
AOI21X1 AOI21X1_1874 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe44_bF_buf3), .B(_10894_), .C(micro_hash_ucr_3_pipe46_bF_buf3), .Y(_10895_) );
AOI21X1 AOI21X1_1875 ( .gnd(gnd), .vdd(vdd), .A(_10469_), .B(_10525_), .C(_10524_), .Y(_10896_) );
INVX1 INVX1_681 ( .gnd(gnd), .vdd(vdd), .A(_10896_), .Y(_10897_) );
XNOR2X1 XNOR2X1_424 ( .gnd(gnd), .vdd(vdd), .A(_10739__bF_buf1), .B(_8997_), .Y(_10898_) );
NAND2X1 NAND2X1_1448 ( .gnd(gnd), .vdd(vdd), .A(_10898_), .B(_10897_), .Y(_10899_) );
NOR2X1 NOR2X1_1814 ( .gnd(gnd), .vdd(vdd), .A(_10898_), .B(_10897_), .Y(_10900_) );
NOR2X1 NOR2X1_1815 ( .gnd(gnd), .vdd(vdd), .A(_9306__bF_buf0), .B(_10900_), .Y(_10901_) );
AOI22X1 AOI22X1_78 ( .gnd(gnd), .vdd(vdd), .A(_10899_), .B(_10901_), .C(_10888_), .D(_10895_), .Y(_10902_) );
OAI21X1 OAI21X1_3051 ( .gnd(gnd), .vdd(vdd), .A(_8966_), .B(_10519__bF_buf4), .C(_10649_), .Y(_10903_) );
XNOR2X1 XNOR2X1_425 ( .gnd(gnd), .vdd(vdd), .A(_10739__bF_buf0), .B(_8970_), .Y(_10904_) );
XOR2X1 XOR2X1_175 ( .gnd(gnd), .vdd(vdd), .A(_10904_), .B(_10903_), .Y(_10905_) );
AOI21X1 AOI21X1_1876 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe48_bF_buf0), .B(_10905_), .C(micro_hash_ucr_3_pipe50_bF_buf1), .Y(_10906_) );
OAI21X1 OAI21X1_3052 ( .gnd(gnd), .vdd(vdd), .A(_10902_), .B(micro_hash_ucr_3_pipe48_bF_buf4), .C(_10906_), .Y(_10907_) );
OR2X2 OR2X2_74 ( .gnd(gnd), .vdd(vdd), .A(_10657_), .B(_10655_), .Y(_10908_) );
OAI21X1 OAI21X1_3053 ( .gnd(gnd), .vdd(vdd), .A(_10737__bF_buf3), .B(_10738__bF_buf3), .C(_8840_), .Y(_10909_) );
NOR2X1 NOR2X1_1816 ( .gnd(gnd), .vdd(vdd), .A(_8840_), .B(_10798__bF_buf0), .Y(_10910_) );
INVX1 INVX1_682 ( .gnd(gnd), .vdd(vdd), .A(_10910_), .Y(_10911_) );
NAND2X1 NAND2X1_1449 ( .gnd(gnd), .vdd(vdd), .A(_10909_), .B(_10911_), .Y(_10912_) );
XOR2X1 XOR2X1_176 ( .gnd(gnd), .vdd(vdd), .A(_10912_), .B(_10908_), .Y(_10913_) );
AOI21X1 AOI21X1_1877 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe50_bF_buf0), .B(_10913_), .C(micro_hash_ucr_3_pipe52_bF_buf3), .Y(_10914_) );
OAI21X1 OAI21X1_3054 ( .gnd(gnd), .vdd(vdd), .A(_9073_), .B(_10519__bF_buf3), .C(_10664_), .Y(_10915_) );
XNOR2X1 XNOR2X1_426 ( .gnd(gnd), .vdd(vdd), .A(_10739__bF_buf3), .B(_9077_), .Y(_10916_) );
NAND2X1 NAND2X1_1450 ( .gnd(gnd), .vdd(vdd), .A(_10915_), .B(_10916_), .Y(_10917_) );
INVX1 INVX1_683 ( .gnd(gnd), .vdd(vdd), .A(_10917_), .Y(_10918_) );
OAI21X1 OAI21X1_3055 ( .gnd(gnd), .vdd(vdd), .A(_10916_), .B(_10915_), .C(micro_hash_ucr_3_pipe52_bF_buf2), .Y(_10919_) );
OAI21X1 OAI21X1_3056 ( .gnd(gnd), .vdd(vdd), .A(_10918_), .B(_10919_), .C(_9298__bF_buf1), .Y(_10920_) );
AOI21X1 AOI21X1_1878 ( .gnd(gnd), .vdd(vdd), .A(_10914_), .B(_10907_), .C(_10920_), .Y(_10921_) );
NAND2X1 NAND2X1_1451 ( .gnd(gnd), .vdd(vdd), .A(_10482_), .B(_10667_), .Y(_10922_) );
OAI21X1 OAI21X1_3057 ( .gnd(gnd), .vdd(vdd), .A(_9044_), .B(_10519__bF_buf2), .C(_10922_), .Y(_10923_) );
OAI21X1 OAI21X1_3058 ( .gnd(gnd), .vdd(vdd), .A(_10737__bF_buf2), .B(_10738__bF_buf2), .C(_9048_), .Y(_10924_) );
NOR2X1 NOR2X1_1817 ( .gnd(gnd), .vdd(vdd), .A(_9048_), .B(_10798__bF_buf5), .Y(_10925_) );
INVX1 INVX1_684 ( .gnd(gnd), .vdd(vdd), .A(_10925_), .Y(_10926_) );
NAND2X1 NAND2X1_1452 ( .gnd(gnd), .vdd(vdd), .A(_10924_), .B(_10926_), .Y(_10927_) );
XNOR2X1 XNOR2X1_427 ( .gnd(gnd), .vdd(vdd), .A(_10927_), .B(_10923_), .Y(_10928_) );
OAI21X1 OAI21X1_3059 ( .gnd(gnd), .vdd(vdd), .A(_10928_), .B(_9298__bF_buf0), .C(_9293__bF_buf2), .Y(_10929_) );
XNOR2X1 XNOR2X1_428 ( .gnd(gnd), .vdd(vdd), .A(_10739__bF_buf2), .B(_8941_), .Y(_10930_) );
OAI21X1 OAI21X1_3060 ( .gnd(gnd), .vdd(vdd), .A(_10675_), .B(_10671_), .C(_10930_), .Y(_10931_) );
INVX1 INVX1_685 ( .gnd(gnd), .vdd(vdd), .A(_10931_), .Y(_10932_) );
OAI21X1 OAI21X1_3061 ( .gnd(gnd), .vdd(vdd), .A(_8937_), .B(_10519__bF_buf1), .C(_10674_), .Y(_10933_) );
OAI21X1 OAI21X1_3062 ( .gnd(gnd), .vdd(vdd), .A(_10933_), .B(_10930_), .C(micro_hash_ucr_3_pipe56_bF_buf1), .Y(_10934_) );
OAI22X1 OAI22X1_139 ( .gnd(gnd), .vdd(vdd), .A(_10932_), .B(_10934_), .C(_10921_), .D(_10929_), .Y(_10935_) );
OAI21X1 OAI21X1_3063 ( .gnd(gnd), .vdd(vdd), .A(_10680_), .B(_10679_), .C(_10681_), .Y(_10936_) );
OAI21X1 OAI21X1_3064 ( .gnd(gnd), .vdd(vdd), .A(_10737__bF_buf1), .B(_10738__bF_buf1), .C(_8998_), .Y(_10937_) );
NOR2X1 NOR2X1_1818 ( .gnd(gnd), .vdd(vdd), .A(_8998_), .B(_10798__bF_buf4), .Y(_10938_) );
INVX1 INVX1_686 ( .gnd(gnd), .vdd(vdd), .A(_10938_), .Y(_10939_) );
NAND2X1 NAND2X1_1453 ( .gnd(gnd), .vdd(vdd), .A(_10937_), .B(_10939_), .Y(_10940_) );
XOR2X1 XOR2X1_177 ( .gnd(gnd), .vdd(vdd), .A(_10940_), .B(_10936_), .Y(_10941_) );
AOI21X1 AOI21X1_1879 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe58_bF_buf0), .B(_10941_), .C(micro_hash_ucr_3_pipe60_bF_buf1), .Y(_10942_) );
OAI21X1 OAI21X1_3065 ( .gnd(gnd), .vdd(vdd), .A(_10935_), .B(micro_hash_ucr_3_pipe58_bF_buf3), .C(_10942_), .Y(_10943_) );
XNOR2X1 XNOR2X1_429 ( .gnd(gnd), .vdd(vdd), .A(_10739__bF_buf1), .B(_8971_), .Y(_10944_) );
OAI21X1 OAI21X1_3066 ( .gnd(gnd), .vdd(vdd), .A(_10693_), .B(_10690_), .C(_10944_), .Y(_10945_) );
INVX1 INVX1_687 ( .gnd(gnd), .vdd(vdd), .A(_10945_), .Y(_10946_) );
OAI21X1 OAI21X1_3067 ( .gnd(gnd), .vdd(vdd), .A(_8967_), .B(_10519__bF_buf0), .C(_10692_), .Y(_10947_) );
OAI21X1 OAI21X1_3068 ( .gnd(gnd), .vdd(vdd), .A(_10947_), .B(_10944_), .C(micro_hash_ucr_3_pipe60_bF_buf0), .Y(_10948_) );
OAI21X1 OAI21X1_3069 ( .gnd(gnd), .vdd(vdd), .A(_10946_), .B(_10948_), .C(_10943_), .Y(_10949_) );
NOR2X1 NOR2X1_1819 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe62_bF_buf2), .B(_10949_), .Y(_10950_) );
NAND2X1 NAND2X1_1454 ( .gnd(gnd), .vdd(vdd), .A(_10496_), .B(_10520_), .Y(_10951_) );
OAI21X1 OAI21X1_3070 ( .gnd(gnd), .vdd(vdd), .A(_8837_), .B(_10519__bF_buf5), .C(_10951_), .Y(_10952_) );
OAI21X1 OAI21X1_3071 ( .gnd(gnd), .vdd(vdd), .A(_10737__bF_buf0), .B(_10738__bF_buf0), .C(_8841_), .Y(_10953_) );
NOR2X1 NOR2X1_1820 ( .gnd(gnd), .vdd(vdd), .A(_8841_), .B(_10798__bF_buf3), .Y(_10954_) );
INVX1 INVX1_688 ( .gnd(gnd), .vdd(vdd), .A(_10954_), .Y(_10955_) );
NAND2X1 NAND2X1_1455 ( .gnd(gnd), .vdd(vdd), .A(_10953_), .B(_10955_), .Y(_10956_) );
XNOR2X1 XNOR2X1_430 ( .gnd(gnd), .vdd(vdd), .A(_10956_), .B(_10952_), .Y(_10957_) );
OAI21X1 OAI21X1_3072 ( .gnd(gnd), .vdd(vdd), .A(_10957_), .B(_9287__bF_buf1), .C(_9288__bF_buf2), .Y(_10958_) );
INVX2 INVX2_375 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_226_), .Y(_10959_) );
XNOR2X1 XNOR2X1_431 ( .gnd(gnd), .vdd(vdd), .A(_10739__bF_buf0), .B(_10959_), .Y(_10960_) );
OAI21X1 OAI21X1_3073 ( .gnd(gnd), .vdd(vdd), .A(_10703_), .B(_10700_), .C(_10960_), .Y(_10961_) );
INVX1 INVX1_689 ( .gnd(gnd), .vdd(vdd), .A(_10961_), .Y(_10962_) );
OAI21X1 OAI21X1_3074 ( .gnd(gnd), .vdd(vdd), .A(_10699_), .B(_10519__bF_buf4), .C(_10702_), .Y(_10963_) );
OAI21X1 OAI21X1_3075 ( .gnd(gnd), .vdd(vdd), .A(_10963_), .B(_10960_), .C(micro_hash_ucr_3_pipe64_bF_buf1), .Y(_10964_) );
OAI22X1 OAI22X1_140 ( .gnd(gnd), .vdd(vdd), .A(_10962_), .B(_10964_), .C(_10950_), .D(_10958_), .Y(_10965_) );
NOR2X1 NOR2X1_1821 ( .gnd(gnd), .vdd(vdd), .A(_10708_), .B(_10710_), .Y(_10966_) );
INVX2 INVX2_376 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_234_), .Y(_10967_) );
XNOR2X1 XNOR2X1_432 ( .gnd(gnd), .vdd(vdd), .A(_10739__bF_buf3), .B(_10967_), .Y(_10968_) );
XOR2X1 XOR2X1_178 ( .gnd(gnd), .vdd(vdd), .A(_10966_), .B(_10968_), .Y(_10969_) );
OAI21X1 OAI21X1_3076 ( .gnd(gnd), .vdd(vdd), .A(_10969_), .B(_9286__bF_buf1), .C(_9282__bF_buf2), .Y(_10970_) );
AOI21X1 AOI21X1_1880 ( .gnd(gnd), .vdd(vdd), .A(_9286__bF_buf0), .B(_10965_), .C(_10970_), .Y(_10971_) );
INVX1 INVX1_690 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_241_), .Y(_10972_) );
OAI21X1 OAI21X1_3077 ( .gnd(gnd), .vdd(vdd), .A(_10972_), .B(_10519__bF_buf3), .C(_10715_), .Y(_10973_) );
INVX2 INVX2_377 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_242_), .Y(_10974_) );
OAI21X1 OAI21X1_3078 ( .gnd(gnd), .vdd(vdd), .A(_10737__bF_buf3), .B(_10738__bF_buf3), .C(_10974_), .Y(_10975_) );
NOR2X1 NOR2X1_1822 ( .gnd(gnd), .vdd(vdd), .A(_10974_), .B(_10798__bF_buf2), .Y(_10976_) );
INVX1 INVX1_691 ( .gnd(gnd), .vdd(vdd), .A(_10976_), .Y(_10977_) );
NAND2X1 NAND2X1_1456 ( .gnd(gnd), .vdd(vdd), .A(_10975_), .B(_10977_), .Y(_10978_) );
XNOR2X1 XNOR2X1_433 ( .gnd(gnd), .vdd(vdd), .A(_10978_), .B(_10973_), .Y(_10979_) );
OAI21X1 OAI21X1_3079 ( .gnd(gnd), .vdd(vdd), .A(_10979_), .B(_9282__bF_buf1), .C(_10380_), .Y(_10980_) );
NAND2X1 NAND2X1_1457 ( .gnd(gnd), .vdd(vdd), .A(_10719_), .B(_10723_), .Y(_10981_) );
OAI21X1 OAI21X1_3080 ( .gnd(gnd), .vdd(vdd), .A(_10721_), .B(_10519__bF_buf2), .C(_10981_), .Y(_10982_) );
INVX1 INVX1_692 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_250_), .Y(_10983_) );
OAI21X1 OAI21X1_3081 ( .gnd(gnd), .vdd(vdd), .A(_10737__bF_buf2), .B(_10738__bF_buf2), .C(_10983_), .Y(_10984_) );
INVX1 INVX1_693 ( .gnd(gnd), .vdd(vdd), .A(_10984_), .Y(_10985_) );
NOR2X1 NOR2X1_1823 ( .gnd(gnd), .vdd(vdd), .A(_10983_), .B(_10798__bF_buf1), .Y(_10986_) );
NOR2X1 NOR2X1_1824 ( .gnd(gnd), .vdd(vdd), .A(_10985_), .B(_10986_), .Y(_10987_) );
AND2X2 AND2X2_710 ( .gnd(gnd), .vdd(vdd), .A(_10987_), .B(_10982_), .Y(_10988_) );
OAI21X1 OAI21X1_3082 ( .gnd(gnd), .vdd(vdd), .A(_10987_), .B(_10982_), .C(_8772_), .Y(_10989_) );
OAI22X1 OAI22X1_141 ( .gnd(gnd), .vdd(vdd), .A(_10988_), .B(_10989_), .C(_10971_), .D(_10980_), .Y(_8702__2_) );
OAI21X1 OAI21X1_3083 ( .gnd(gnd), .vdd(vdd), .A(_10710_), .B(_10708_), .C(_10968_), .Y(_10990_) );
OAI21X1 OAI21X1_3084 ( .gnd(gnd), .vdd(vdd), .A(_10967_), .B(_10798__bF_buf0), .C(_10990_), .Y(_10991_) );
XOR2X1 XOR2X1_179 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_k_3_), .B(micro_hash_ucr_3_x_3_), .Y(_10992_) );
OAI21X1 OAI21X1_3085 ( .gnd(gnd), .vdd(vdd), .A(_10737__bF_buf1), .B(_10734_), .C(_10992_), .Y(_10993_) );
INVX8 INVX8_280 ( .gnd(gnd), .vdd(vdd), .A(_10993_), .Y(_10994_) );
OAI21X1 OAI21X1_3086 ( .gnd(gnd), .vdd(vdd), .A(_10730_), .B(_10736_), .C(_10735_), .Y(_10995_) );
NOR2X1 NOR2X1_1825 ( .gnd(gnd), .vdd(vdd), .A(_10992_), .B(_10995_), .Y(_10996_) );
NOR2X1 NOR2X1_1826 ( .gnd(gnd), .vdd(vdd), .A(_10996__bF_buf4), .B(_10994__bF_buf4), .Y(_10997_) );
NOR2X1 NOR2X1_1827 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_235_), .B(_10997_), .Y(_10998_) );
INVX1 INVX1_694 ( .gnd(gnd), .vdd(vdd), .A(_10998_), .Y(_10999_) );
NAND2X1 NAND2X1_1458 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_235_), .B(_10997_), .Y(_11000_) );
NAND2X1 NAND2X1_1459 ( .gnd(gnd), .vdd(vdd), .A(_11000_), .B(_10999_), .Y(_11001_) );
XOR2X1 XOR2X1_180 ( .gnd(gnd), .vdd(vdd), .A(_11001_), .B(_10991_), .Y(_11002_) );
NAND2X1 NAND2X1_1460 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_26_), .B(_10739__bF_buf2), .Y(_11003_) );
OAI21X1 OAI21X1_3087 ( .gnd(gnd), .vdd(vdd), .A(_10765_), .B(_10764_), .C(_11003_), .Y(_11004_) );
INVX1 INVX1_695 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_27_), .Y(_11005_) );
OAI21X1 OAI21X1_3088 ( .gnd(gnd), .vdd(vdd), .A(_10994__bF_buf3), .B(_10996__bF_buf3), .C(_11005_), .Y(_11006_) );
INVX1 INVX1_696 ( .gnd(gnd), .vdd(vdd), .A(_11006_), .Y(_11007_) );
INVX8 INVX8_281 ( .gnd(gnd), .vdd(vdd), .A(_10997_), .Y(_11008_) );
NOR2X1 NOR2X1_1828 ( .gnd(gnd), .vdd(vdd), .A(_11005_), .B(_11008__bF_buf4), .Y(_11009_) );
NOR2X1 NOR2X1_1829 ( .gnd(gnd), .vdd(vdd), .A(_11007_), .B(_11009_), .Y(_11010_) );
XOR2X1 XOR2X1_181 ( .gnd(gnd), .vdd(vdd), .A(_11010_), .B(_11004_), .Y(_11011_) );
AOI21X1 AOI21X1_1881 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_2_), .B(_10739__bF_buf1), .C(_10753_), .Y(_11012_) );
INVX2 INVX2_378 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_3_), .Y(_11013_) );
XNOR2X1 XNOR2X1_434 ( .gnd(gnd), .vdd(vdd), .A(_10997_), .B(_11013_), .Y(_11014_) );
OAI21X1 OAI21X1_3089 ( .gnd(gnd), .vdd(vdd), .A(_11012_), .B(_11014_), .C(micro_hash_ucr_3_pipe8), .Y(_11015_) );
AOI21X1 AOI21X1_1882 ( .gnd(gnd), .vdd(vdd), .A(_11012_), .B(_11014_), .C(_11015_), .Y(_11016_) );
AND2X2 AND2X2_711 ( .gnd(gnd), .vdd(vdd), .A(H_3_19_), .B(micro_hash_ucr_3_pipe6_bF_buf3), .Y(_11017_) );
OAI21X1 OAI21X1_3090 ( .gnd(gnd), .vdd(vdd), .A(_9701__bF_buf2), .B(micro_hash_ucr_3_pipe6_bF_buf2), .C(_9341_), .Y(_11018_) );
OAI21X1 OAI21X1_3091 ( .gnd(gnd), .vdd(vdd), .A(_11018_), .B(_11017_), .C(_9342_), .Y(_11019_) );
NOR2X1 NOR2X1_1830 ( .gnd(gnd), .vdd(vdd), .A(_11019_), .B(_11016_), .Y(_11020_) );
OAI21X1 OAI21X1_3092 ( .gnd(gnd), .vdd(vdd), .A(_10745_), .B(_10798__bF_buf5), .C(_10747_), .Y(_11021_) );
INVX1 INVX1_697 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_11_), .Y(_11022_) );
OAI21X1 OAI21X1_3093 ( .gnd(gnd), .vdd(vdd), .A(_10994__bF_buf2), .B(_10996__bF_buf2), .C(_11022_), .Y(_11023_) );
NAND2X1 NAND2X1_1461 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_11_), .B(_10997_), .Y(_11024_) );
NAND2X1 NAND2X1_1462 ( .gnd(gnd), .vdd(vdd), .A(_11023_), .B(_11024_), .Y(_11025_) );
XOR2X1 XOR2X1_182 ( .gnd(gnd), .vdd(vdd), .A(_11025_), .B(_11021_), .Y(_11026_) );
OAI21X1 OAI21X1_3094 ( .gnd(gnd), .vdd(vdd), .A(_11026_), .B(_9342_), .C(_9340_), .Y(_11027_) );
AOI21X1 AOI21X1_1883 ( .gnd(gnd), .vdd(vdd), .A(_10728_), .B(_10742_), .C(_10741_), .Y(_11028_) );
INVX1 INVX1_698 ( .gnd(gnd), .vdd(vdd), .A(_11028_), .Y(_11029_) );
INVX1 INVX1_699 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_19_), .Y(_11030_) );
OAI21X1 OAI21X1_3095 ( .gnd(gnd), .vdd(vdd), .A(_10994__bF_buf1), .B(_10996__bF_buf1), .C(_11030_), .Y(_11031_) );
NOR2X1 NOR2X1_1831 ( .gnd(gnd), .vdd(vdd), .A(_11030_), .B(_11008__bF_buf3), .Y(_11032_) );
INVX1 INVX1_700 ( .gnd(gnd), .vdd(vdd), .A(_11032_), .Y(_11033_) );
NAND2X1 NAND2X1_1463 ( .gnd(gnd), .vdd(vdd), .A(_11031_), .B(_11033_), .Y(_11034_) );
AOI21X1 AOI21X1_1884 ( .gnd(gnd), .vdd(vdd), .A(_11029_), .B(_11034_), .C(_9340_), .Y(_11035_) );
OAI21X1 OAI21X1_3096 ( .gnd(gnd), .vdd(vdd), .A(_11029_), .B(_11034_), .C(_11035_), .Y(_11036_) );
OAI21X1 OAI21X1_3097 ( .gnd(gnd), .vdd(vdd), .A(_11020_), .B(_11027_), .C(_11036_), .Y(_11037_) );
NAND2X1 NAND2X1_1464 ( .gnd(gnd), .vdd(vdd), .A(_9335__bF_buf3), .B(_11037_), .Y(_11038_) );
OAI21X1 OAI21X1_3098 ( .gnd(gnd), .vdd(vdd), .A(_9335__bF_buf2), .B(_11011_), .C(_11038_), .Y(_11039_) );
NAND2X1 NAND2X1_1465 ( .gnd(gnd), .vdd(vdd), .A(_9336__bF_buf0), .B(_11039_), .Y(_11040_) );
OAI21X1 OAI21X1_3099 ( .gnd(gnd), .vdd(vdd), .A(_10771_), .B(_10798__bF_buf4), .C(_10774_), .Y(_11041_) );
INVX1 INVX1_701 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_35_), .Y(_11042_) );
OAI21X1 OAI21X1_3100 ( .gnd(gnd), .vdd(vdd), .A(_10994__bF_buf0), .B(_10996__bF_buf0), .C(_11042_), .Y(_11043_) );
NOR2X1 NOR2X1_1832 ( .gnd(gnd), .vdd(vdd), .A(_11042_), .B(_11008__bF_buf2), .Y(_11044_) );
INVX1 INVX1_702 ( .gnd(gnd), .vdd(vdd), .A(_11044_), .Y(_11045_) );
NAND2X1 NAND2X1_1466 ( .gnd(gnd), .vdd(vdd), .A(_11043_), .B(_11045_), .Y(_11046_) );
AOI21X1 AOI21X1_1885 ( .gnd(gnd), .vdd(vdd), .A(_11041_), .B(_11046_), .C(_9336__bF_buf3), .Y(_11047_) );
OAI21X1 OAI21X1_3101 ( .gnd(gnd), .vdd(vdd), .A(_11041_), .B(_11046_), .C(_11047_), .Y(_11048_) );
AND2X2 AND2X2_712 ( .gnd(gnd), .vdd(vdd), .A(_11048_), .B(_9334__bF_buf0), .Y(_11049_) );
OAI21X1 OAI21X1_3102 ( .gnd(gnd), .vdd(vdd), .A(_10779_), .B(_10798__bF_buf3), .C(_10782_), .Y(_11050_) );
INVX1 INVX1_703 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_43_), .Y(_11051_) );
OAI21X1 OAI21X1_3103 ( .gnd(gnd), .vdd(vdd), .A(_10994__bF_buf4), .B(_10996__bF_buf4), .C(_11051_), .Y(_11052_) );
NOR2X1 NOR2X1_1833 ( .gnd(gnd), .vdd(vdd), .A(_11051_), .B(_11008__bF_buf1), .Y(_11053_) );
INVX1 INVX1_704 ( .gnd(gnd), .vdd(vdd), .A(_11053_), .Y(_11054_) );
AOI21X1 AOI21X1_1886 ( .gnd(gnd), .vdd(vdd), .A(_11052_), .B(_11054_), .C(_11050_), .Y(_11055_) );
INVX1 INVX1_705 ( .gnd(gnd), .vdd(vdd), .A(_11050_), .Y(_11056_) );
NAND2X1 NAND2X1_1467 ( .gnd(gnd), .vdd(vdd), .A(_11052_), .B(_11054_), .Y(_11057_) );
OAI21X1 OAI21X1_3104 ( .gnd(gnd), .vdd(vdd), .A(_11057_), .B(_11056_), .C(micro_hash_ucr_3_pipe18_bF_buf0), .Y(_11058_) );
OAI21X1 OAI21X1_3105 ( .gnd(gnd), .vdd(vdd), .A(_11058_), .B(_11055_), .C(_9329__bF_buf4), .Y(_11059_) );
AOI21X1 AOI21X1_1887 ( .gnd(gnd), .vdd(vdd), .A(_11049_), .B(_11040_), .C(_11059_), .Y(_11060_) );
OAI21X1 OAI21X1_3106 ( .gnd(gnd), .vdd(vdd), .A(_10787_), .B(_10798__bF_buf2), .C(_10790_), .Y(_11061_) );
INVX1 INVX1_706 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_51_), .Y(_11062_) );
OAI21X1 OAI21X1_3107 ( .gnd(gnd), .vdd(vdd), .A(_10994__bF_buf3), .B(_10996__bF_buf3), .C(_11062_), .Y(_11063_) );
NOR2X1 NOR2X1_1834 ( .gnd(gnd), .vdd(vdd), .A(_11062_), .B(_11008__bF_buf0), .Y(_11064_) );
INVX1 INVX1_707 ( .gnd(gnd), .vdd(vdd), .A(_11064_), .Y(_11065_) );
NAND2X1 NAND2X1_1468 ( .gnd(gnd), .vdd(vdd), .A(_11063_), .B(_11065_), .Y(_11066_) );
XNOR2X1 XNOR2X1_435 ( .gnd(gnd), .vdd(vdd), .A(_11066_), .B(_11061_), .Y(_11067_) );
OAI21X1 OAI21X1_3108 ( .gnd(gnd), .vdd(vdd), .A(_11067_), .B(_9329__bF_buf3), .C(_9330__bF_buf3), .Y(_11068_) );
NOR2X1 NOR2X1_1835 ( .gnd(gnd), .vdd(vdd), .A(_10799_), .B(_10800_), .Y(_11069_) );
OAI21X1 OAI21X1_3109 ( .gnd(gnd), .vdd(vdd), .A(_10994__bF_buf2), .B(_10996__bF_buf2), .C(_9269_), .Y(_11070_) );
INVX1 INVX1_708 ( .gnd(gnd), .vdd(vdd), .A(_11070_), .Y(_11071_) );
NOR2X1 NOR2X1_1836 ( .gnd(gnd), .vdd(vdd), .A(_9269_), .B(_11008__bF_buf4), .Y(_11072_) );
NOR2X1 NOR2X1_1837 ( .gnd(gnd), .vdd(vdd), .A(_11071_), .B(_11072_), .Y(_11073_) );
XNOR2X1 XNOR2X1_436 ( .gnd(gnd), .vdd(vdd), .A(_11073_), .B(_11069_), .Y(_11074_) );
AOI21X1 AOI21X1_1888 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe22_bF_buf0), .B(_11074_), .C(micro_hash_ucr_3_pipe24_bF_buf0), .Y(_11075_) );
OAI21X1 OAI21X1_3110 ( .gnd(gnd), .vdd(vdd), .A(_11060_), .B(_11068_), .C(_11075_), .Y(_11076_) );
NAND3X1 NAND3X1_581 ( .gnd(gnd), .vdd(vdd), .A(_10805_), .B(_10806_), .C(_10808_), .Y(_11077_) );
OAI21X1 OAI21X1_3111 ( .gnd(gnd), .vdd(vdd), .A(_9243_), .B(_10798__bF_buf1), .C(_11077_), .Y(_11078_) );
OAI21X1 OAI21X1_3112 ( .gnd(gnd), .vdd(vdd), .A(_10994__bF_buf1), .B(_10996__bF_buf1), .C(_9246_), .Y(_11079_) );
NOR2X1 NOR2X1_1838 ( .gnd(gnd), .vdd(vdd), .A(_9246_), .B(_11008__bF_buf3), .Y(_11080_) );
INVX1 INVX1_709 ( .gnd(gnd), .vdd(vdd), .A(_11080_), .Y(_11081_) );
NAND2X1 NAND2X1_1469 ( .gnd(gnd), .vdd(vdd), .A(_11079_), .B(_11081_), .Y(_11082_) );
AOI21X1 AOI21X1_1889 ( .gnd(gnd), .vdd(vdd), .A(_11078_), .B(_11082_), .C(_9328__bF_buf0), .Y(_11083_) );
OAI21X1 OAI21X1_3113 ( .gnd(gnd), .vdd(vdd), .A(_11078_), .B(_11082_), .C(_11083_), .Y(_11084_) );
AND2X2 AND2X2_713 ( .gnd(gnd), .vdd(vdd), .A(_11084_), .B(_9323__bF_buf2), .Y(_11085_) );
OAI21X1 OAI21X1_3114 ( .gnd(gnd), .vdd(vdd), .A(_9165_), .B(_10798__bF_buf0), .C(_10815_), .Y(_11086_) );
OAI21X1 OAI21X1_3115 ( .gnd(gnd), .vdd(vdd), .A(_10994__bF_buf0), .B(_10996__bF_buf0), .C(_9168_), .Y(_11087_) );
NOR2X1 NOR2X1_1839 ( .gnd(gnd), .vdd(vdd), .A(_9168_), .B(_11008__bF_buf2), .Y(_11088_) );
INVX1 INVX1_710 ( .gnd(gnd), .vdd(vdd), .A(_11088_), .Y(_11089_) );
AOI21X1 AOI21X1_1890 ( .gnd(gnd), .vdd(vdd), .A(_11087_), .B(_11089_), .C(_11086_), .Y(_11090_) );
INVX1 INVX1_711 ( .gnd(gnd), .vdd(vdd), .A(_11086_), .Y(_11091_) );
NAND2X1 NAND2X1_1470 ( .gnd(gnd), .vdd(vdd), .A(_11087_), .B(_11089_), .Y(_11092_) );
OAI21X1 OAI21X1_3116 ( .gnd(gnd), .vdd(vdd), .A(_11092_), .B(_11091_), .C(micro_hash_ucr_3_pipe26_bF_buf3), .Y(_11093_) );
OAI21X1 OAI21X1_3117 ( .gnd(gnd), .vdd(vdd), .A(_11093_), .B(_11090_), .C(_9324__bF_buf2), .Y(_11094_) );
AOI21X1 AOI21X1_1891 ( .gnd(gnd), .vdd(vdd), .A(_11085_), .B(_11076_), .C(_11094_), .Y(_11095_) );
NAND3X1 NAND3X1_582 ( .gnd(gnd), .vdd(vdd), .A(_10819_), .B(_10820_), .C(_10822_), .Y(_11096_) );
OAI21X1 OAI21X1_3118 ( .gnd(gnd), .vdd(vdd), .A(_9220_), .B(_10798__bF_buf5), .C(_11096_), .Y(_11097_) );
OAI21X1 OAI21X1_3119 ( .gnd(gnd), .vdd(vdd), .A(_10994__bF_buf4), .B(_10996__bF_buf4), .C(_9223_), .Y(_11098_) );
NOR2X1 NOR2X1_1840 ( .gnd(gnd), .vdd(vdd), .A(_9223_), .B(_11008__bF_buf1), .Y(_11099_) );
INVX1 INVX1_712 ( .gnd(gnd), .vdd(vdd), .A(_11099_), .Y(_11100_) );
NAND2X1 NAND2X1_1471 ( .gnd(gnd), .vdd(vdd), .A(_11098_), .B(_11100_), .Y(_11101_) );
XNOR2X1 XNOR2X1_437 ( .gnd(gnd), .vdd(vdd), .A(_11101_), .B(_11097_), .Y(_11102_) );
OAI21X1 OAI21X1_3120 ( .gnd(gnd), .vdd(vdd), .A(_11102_), .B(_9324__bF_buf1), .C(_9322__bF_buf1), .Y(_11103_) );
OAI21X1 OAI21X1_3121 ( .gnd(gnd), .vdd(vdd), .A(_9190_), .B(_10798__bF_buf4), .C(_10831_), .Y(_11104_) );
OAI21X1 OAI21X1_3122 ( .gnd(gnd), .vdd(vdd), .A(_10994__bF_buf3), .B(_10996__bF_buf3), .C(_9194_), .Y(_11105_) );
INVX1 INVX1_713 ( .gnd(gnd), .vdd(vdd), .A(_11105_), .Y(_11106_) );
NOR2X1 NOR2X1_1841 ( .gnd(gnd), .vdd(vdd), .A(_9194_), .B(_11008__bF_buf0), .Y(_11107_) );
NOR2X1 NOR2X1_1842 ( .gnd(gnd), .vdd(vdd), .A(_11106_), .B(_11107_), .Y(_11108_) );
XOR2X1 XOR2X1_183 ( .gnd(gnd), .vdd(vdd), .A(_11108_), .B(_11104_), .Y(_11109_) );
AOI21X1 AOI21X1_1892 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe30_bF_buf1), .B(_11109_), .C(micro_hash_ucr_3_pipe32_bF_buf1), .Y(_11110_) );
OAI21X1 OAI21X1_3123 ( .gnd(gnd), .vdd(vdd), .A(_11095_), .B(_11103_), .C(_11110_), .Y(_11111_) );
NAND3X1 NAND3X1_583 ( .gnd(gnd), .vdd(vdd), .A(_10836_), .B(_10837_), .C(_10839_), .Y(_11112_) );
OAI21X1 OAI21X1_3124 ( .gnd(gnd), .vdd(vdd), .A(_9047_), .B(_10798__bF_buf3), .C(_11112_), .Y(_11113_) );
OAI21X1 OAI21X1_3125 ( .gnd(gnd), .vdd(vdd), .A(_10994__bF_buf2), .B(_10996__bF_buf2), .C(_9051_), .Y(_11114_) );
NOR2X1 NOR2X1_1843 ( .gnd(gnd), .vdd(vdd), .A(_9051_), .B(_11008__bF_buf4), .Y(_11115_) );
INVX1 INVX1_714 ( .gnd(gnd), .vdd(vdd), .A(_11115_), .Y(_11116_) );
NAND2X1 NAND2X1_1472 ( .gnd(gnd), .vdd(vdd), .A(_11114_), .B(_11116_), .Y(_11117_) );
AOI21X1 AOI21X1_1893 ( .gnd(gnd), .vdd(vdd), .A(_11113_), .B(_11117_), .C(_9317__bF_buf1), .Y(_11118_) );
OAI21X1 OAI21X1_3126 ( .gnd(gnd), .vdd(vdd), .A(_11113_), .B(_11117_), .C(_11118_), .Y(_11119_) );
AND2X2 AND2X2_714 ( .gnd(gnd), .vdd(vdd), .A(_11119_), .B(_9318__bF_buf2), .Y(_11120_) );
OAI21X1 OAI21X1_3127 ( .gnd(gnd), .vdd(vdd), .A(_9142_), .B(_10798__bF_buf2), .C(_10849_), .Y(_11121_) );
OAI21X1 OAI21X1_3128 ( .gnd(gnd), .vdd(vdd), .A(_10994__bF_buf1), .B(_10996__bF_buf1), .C(_9145_), .Y(_11122_) );
NOR2X1 NOR2X1_1844 ( .gnd(gnd), .vdd(vdd), .A(_9145_), .B(_11008__bF_buf3), .Y(_11123_) );
INVX1 INVX1_715 ( .gnd(gnd), .vdd(vdd), .A(_11123_), .Y(_11124_) );
NAND2X1 NAND2X1_1473 ( .gnd(gnd), .vdd(vdd), .A(_11122_), .B(_11124_), .Y(_11125_) );
XOR2X1 XOR2X1_184 ( .gnd(gnd), .vdd(vdd), .A(_11125_), .B(_11121_), .Y(_11126_) );
OAI21X1 OAI21X1_3129 ( .gnd(gnd), .vdd(vdd), .A(_11126_), .B(_9318__bF_buf1), .C(_9316__bF_buf1), .Y(_11127_) );
AOI21X1 AOI21X1_1894 ( .gnd(gnd), .vdd(vdd), .A(_11120_), .B(_11111_), .C(_11127_), .Y(_11128_) );
NAND3X1 NAND3X1_584 ( .gnd(gnd), .vdd(vdd), .A(_10852_), .B(_10853_), .C(_10855_), .Y(_11129_) );
OAI21X1 OAI21X1_3130 ( .gnd(gnd), .vdd(vdd), .A(_9120_), .B(_10798__bF_buf1), .C(_11129_), .Y(_11130_) );
OAI21X1 OAI21X1_3131 ( .gnd(gnd), .vdd(vdd), .A(_10994__bF_buf0), .B(_10996__bF_buf0), .C(_9123_), .Y(_11131_) );
NOR2X1 NOR2X1_1845 ( .gnd(gnd), .vdd(vdd), .A(_9123_), .B(_11008__bF_buf2), .Y(_11132_) );
INVX1 INVX1_716 ( .gnd(gnd), .vdd(vdd), .A(_11132_), .Y(_11133_) );
NAND2X1 NAND2X1_1474 ( .gnd(gnd), .vdd(vdd), .A(_11131_), .B(_11133_), .Y(_11134_) );
XNOR2X1 XNOR2X1_438 ( .gnd(gnd), .vdd(vdd), .A(_11134_), .B(_11130_), .Y(_11135_) );
OAI21X1 OAI21X1_3132 ( .gnd(gnd), .vdd(vdd), .A(_11135_), .B(_9316__bF_buf0), .C(_9311__bF_buf0), .Y(_11136_) );
OAI21X1 OAI21X1_3133 ( .gnd(gnd), .vdd(vdd), .A(_9024_), .B(_10798__bF_buf0), .C(_10867_), .Y(_11137_) );
OAI21X1 OAI21X1_3134 ( .gnd(gnd), .vdd(vdd), .A(_10994__bF_buf4), .B(_10996__bF_buf4), .C(_9027_), .Y(_11138_) );
NOR2X1 NOR2X1_1846 ( .gnd(gnd), .vdd(vdd), .A(_9027_), .B(_11008__bF_buf1), .Y(_11139_) );
INVX1 INVX1_717 ( .gnd(gnd), .vdd(vdd), .A(_11139_), .Y(_11140_) );
NAND2X1 NAND2X1_1475 ( .gnd(gnd), .vdd(vdd), .A(_11138_), .B(_11140_), .Y(_11141_) );
XNOR2X1 XNOR2X1_439 ( .gnd(gnd), .vdd(vdd), .A(_11137_), .B(_11141_), .Y(_11142_) );
AOI21X1 AOI21X1_1895 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe38_bF_buf1), .B(_11142_), .C(micro_hash_ucr_3_pipe40_bF_buf2), .Y(_11143_) );
OAI21X1 OAI21X1_3135 ( .gnd(gnd), .vdd(vdd), .A(_11128_), .B(_11136_), .C(_11143_), .Y(_11144_) );
NAND3X1 NAND3X1_585 ( .gnd(gnd), .vdd(vdd), .A(_10872_), .B(_10873_), .C(_10875_), .Y(_11145_) );
OAI21X1 OAI21X1_3136 ( .gnd(gnd), .vdd(vdd), .A(_9076_), .B(_10798__bF_buf5), .C(_11145_), .Y(_11146_) );
OAI21X1 OAI21X1_3137 ( .gnd(gnd), .vdd(vdd), .A(_10994__bF_buf3), .B(_10996__bF_buf3), .C(_9080_), .Y(_11147_) );
NOR2X1 NOR2X1_1847 ( .gnd(gnd), .vdd(vdd), .A(_9080_), .B(_11008__bF_buf0), .Y(_11148_) );
INVX1 INVX1_718 ( .gnd(gnd), .vdd(vdd), .A(_11148_), .Y(_11149_) );
NAND2X1 NAND2X1_1476 ( .gnd(gnd), .vdd(vdd), .A(_11147_), .B(_11149_), .Y(_11150_) );
AOI21X1 AOI21X1_1896 ( .gnd(gnd), .vdd(vdd), .A(_11146_), .B(_11150_), .C(_9312__bF_buf0), .Y(_11151_) );
OAI21X1 OAI21X1_3138 ( .gnd(gnd), .vdd(vdd), .A(_11146_), .B(_11150_), .C(_11151_), .Y(_11152_) );
AND2X2 AND2X2_715 ( .gnd(gnd), .vdd(vdd), .A(_11152_), .B(_9310__bF_buf1), .Y(_11153_) );
OAI21X1 OAI21X1_3139 ( .gnd(gnd), .vdd(vdd), .A(_9191_), .B(_10798__bF_buf4), .C(_10885_), .Y(_11154_) );
OAI21X1 OAI21X1_3140 ( .gnd(gnd), .vdd(vdd), .A(_10994__bF_buf2), .B(_10996__bF_buf2), .C(_9195_), .Y(_11155_) );
NOR2X1 NOR2X1_1848 ( .gnd(gnd), .vdd(vdd), .A(_9195_), .B(_11008__bF_buf4), .Y(_11156_) );
INVX1 INVX1_719 ( .gnd(gnd), .vdd(vdd), .A(_11156_), .Y(_11157_) );
NAND2X1 NAND2X1_1477 ( .gnd(gnd), .vdd(vdd), .A(_11155_), .B(_11157_), .Y(_11158_) );
XOR2X1 XOR2X1_185 ( .gnd(gnd), .vdd(vdd), .A(_11158_), .B(_11154_), .Y(_11159_) );
OAI21X1 OAI21X1_3141 ( .gnd(gnd), .vdd(vdd), .A(_11159_), .B(_9310__bF_buf0), .C(_9305__bF_buf3), .Y(_11160_) );
AOI21X1 AOI21X1_1897 ( .gnd(gnd), .vdd(vdd), .A(_11153_), .B(_11144_), .C(_11160_), .Y(_11161_) );
NAND3X1 NAND3X1_586 ( .gnd(gnd), .vdd(vdd), .A(_10889_), .B(_10890_), .C(_10892_), .Y(_11162_) );
OAI21X1 OAI21X1_3142 ( .gnd(gnd), .vdd(vdd), .A(_8940_), .B(_10798__bF_buf3), .C(_11162_), .Y(_11163_) );
OAI21X1 OAI21X1_3143 ( .gnd(gnd), .vdd(vdd), .A(_10994__bF_buf1), .B(_10996__bF_buf1), .C(_8944_), .Y(_11164_) );
NOR2X1 NOR2X1_1849 ( .gnd(gnd), .vdd(vdd), .A(_8944_), .B(_11008__bF_buf3), .Y(_11165_) );
INVX1 INVX1_720 ( .gnd(gnd), .vdd(vdd), .A(_11165_), .Y(_11166_) );
NAND2X1 NAND2X1_1478 ( .gnd(gnd), .vdd(vdd), .A(_11164_), .B(_11166_), .Y(_11167_) );
XNOR2X1 XNOR2X1_440 ( .gnd(gnd), .vdd(vdd), .A(_11167_), .B(_11163_), .Y(_11168_) );
OAI21X1 OAI21X1_3144 ( .gnd(gnd), .vdd(vdd), .A(_11168_), .B(_9305__bF_buf2), .C(_9306__bF_buf3), .Y(_11169_) );
OAI21X1 OAI21X1_3145 ( .gnd(gnd), .vdd(vdd), .A(_8997_), .B(_10798__bF_buf2), .C(_10899_), .Y(_11170_) );
OAI21X1 OAI21X1_3146 ( .gnd(gnd), .vdd(vdd), .A(_10994__bF_buf0), .B(_10996__bF_buf0), .C(_9001_), .Y(_11171_) );
INVX1 INVX1_721 ( .gnd(gnd), .vdd(vdd), .A(_11171_), .Y(_11172_) );
NOR2X1 NOR2X1_1850 ( .gnd(gnd), .vdd(vdd), .A(_9001_), .B(_11008__bF_buf2), .Y(_11173_) );
NOR2X1 NOR2X1_1851 ( .gnd(gnd), .vdd(vdd), .A(_11172_), .B(_11173_), .Y(_11174_) );
XOR2X1 XOR2X1_186 ( .gnd(gnd), .vdd(vdd), .A(_11174_), .B(_11170_), .Y(_11175_) );
AOI21X1 AOI21X1_1898 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe46_bF_buf2), .B(_11175_), .C(micro_hash_ucr_3_pipe48_bF_buf3), .Y(_11176_) );
OAI21X1 OAI21X1_3147 ( .gnd(gnd), .vdd(vdd), .A(_11161_), .B(_11169_), .C(_11176_), .Y(_11177_) );
OAI21X1 OAI21X1_3148 ( .gnd(gnd), .vdd(vdd), .A(_10650_), .B(_10646_), .C(_10904_), .Y(_11178_) );
OAI21X1 OAI21X1_3149 ( .gnd(gnd), .vdd(vdd), .A(_8970_), .B(_10798__bF_buf1), .C(_11178_), .Y(_11179_) );
OAI21X1 OAI21X1_3150 ( .gnd(gnd), .vdd(vdd), .A(_10994__bF_buf4), .B(_10996__bF_buf4), .C(_8974_), .Y(_11180_) );
NOR2X1 NOR2X1_1852 ( .gnd(gnd), .vdd(vdd), .A(_8974_), .B(_11008__bF_buf1), .Y(_11181_) );
INVX1 INVX1_722 ( .gnd(gnd), .vdd(vdd), .A(_11181_), .Y(_11182_) );
NAND2X1 NAND2X1_1479 ( .gnd(gnd), .vdd(vdd), .A(_11180_), .B(_11182_), .Y(_11183_) );
AOI21X1 AOI21X1_1899 ( .gnd(gnd), .vdd(vdd), .A(_11179_), .B(_11183_), .C(_9304__bF_buf2), .Y(_11184_) );
OAI21X1 OAI21X1_3151 ( .gnd(gnd), .vdd(vdd), .A(_11179_), .B(_11183_), .C(_11184_), .Y(_11185_) );
AND2X2 AND2X2_716 ( .gnd(gnd), .vdd(vdd), .A(_11185_), .B(_9299__bF_buf2), .Y(_11186_) );
NAND3X1 NAND3X1_587 ( .gnd(gnd), .vdd(vdd), .A(_10909_), .B(_10911_), .C(_10908_), .Y(_11187_) );
OAI21X1 OAI21X1_3152 ( .gnd(gnd), .vdd(vdd), .A(_8840_), .B(_10798__bF_buf0), .C(_11187_), .Y(_11188_) );
OAI21X1 OAI21X1_3153 ( .gnd(gnd), .vdd(vdd), .A(_10994__bF_buf3), .B(_10996__bF_buf3), .C(_8844_), .Y(_11189_) );
NOR2X1 NOR2X1_1853 ( .gnd(gnd), .vdd(vdd), .A(_8844_), .B(_11008__bF_buf0), .Y(_11190_) );
INVX1 INVX1_723 ( .gnd(gnd), .vdd(vdd), .A(_11190_), .Y(_11191_) );
NAND2X1 NAND2X1_1480 ( .gnd(gnd), .vdd(vdd), .A(_11189_), .B(_11191_), .Y(_11192_) );
XOR2X1 XOR2X1_187 ( .gnd(gnd), .vdd(vdd), .A(_11192_), .B(_11188_), .Y(_11193_) );
OAI21X1 OAI21X1_3154 ( .gnd(gnd), .vdd(vdd), .A(_11193_), .B(_9299__bF_buf1), .C(_9300__bF_buf0), .Y(_11194_) );
AOI21X1 AOI21X1_1900 ( .gnd(gnd), .vdd(vdd), .A(_11186_), .B(_11177_), .C(_11194_), .Y(_11195_) );
OAI21X1 OAI21X1_3155 ( .gnd(gnd), .vdd(vdd), .A(_9077_), .B(_10798__bF_buf5), .C(_10917_), .Y(_11196_) );
OAI21X1 OAI21X1_3156 ( .gnd(gnd), .vdd(vdd), .A(_10994__bF_buf2), .B(_10996__bF_buf2), .C(_9081_), .Y(_11197_) );
NOR2X1 NOR2X1_1854 ( .gnd(gnd), .vdd(vdd), .A(_9081_), .B(_11008__bF_buf4), .Y(_11198_) );
INVX1 INVX1_724 ( .gnd(gnd), .vdd(vdd), .A(_11198_), .Y(_11199_) );
NAND2X1 NAND2X1_1481 ( .gnd(gnd), .vdd(vdd), .A(_11197_), .B(_11199_), .Y(_11200_) );
XNOR2X1 XNOR2X1_441 ( .gnd(gnd), .vdd(vdd), .A(_11200_), .B(_11196_), .Y(_11201_) );
OAI21X1 OAI21X1_3157 ( .gnd(gnd), .vdd(vdd), .A(_11201_), .B(_9300__bF_buf3), .C(_9298__bF_buf4), .Y(_11202_) );
NAND3X1 NAND3X1_588 ( .gnd(gnd), .vdd(vdd), .A(_10923_), .B(_10924_), .C(_10926_), .Y(_11203_) );
OAI21X1 OAI21X1_3158 ( .gnd(gnd), .vdd(vdd), .A(_9048_), .B(_10798__bF_buf4), .C(_11203_), .Y(_11204_) );
OAI21X1 OAI21X1_3159 ( .gnd(gnd), .vdd(vdd), .A(_10994__bF_buf1), .B(_10996__bF_buf1), .C(_9052_), .Y(_11205_) );
INVX1 INVX1_725 ( .gnd(gnd), .vdd(vdd), .A(_11205_), .Y(_11206_) );
NOR2X1 NOR2X1_1855 ( .gnd(gnd), .vdd(vdd), .A(_9052_), .B(_11008__bF_buf3), .Y(_11207_) );
NOR2X1 NOR2X1_1856 ( .gnd(gnd), .vdd(vdd), .A(_11206_), .B(_11207_), .Y(_11208_) );
XOR2X1 XOR2X1_188 ( .gnd(gnd), .vdd(vdd), .A(_11208_), .B(_11204_), .Y(_11209_) );
AOI21X1 AOI21X1_1901 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe54_bF_buf2), .B(_11209_), .C(micro_hash_ucr_3_pipe56_bF_buf0), .Y(_11210_) );
OAI21X1 OAI21X1_3160 ( .gnd(gnd), .vdd(vdd), .A(_11195_), .B(_11202_), .C(_11210_), .Y(_11211_) );
OAI21X1 OAI21X1_3161 ( .gnd(gnd), .vdd(vdd), .A(_8941_), .B(_10798__bF_buf3), .C(_10931_), .Y(_11212_) );
OAI21X1 OAI21X1_3162 ( .gnd(gnd), .vdd(vdd), .A(_10994__bF_buf0), .B(_10996__bF_buf0), .C(_8945_), .Y(_11213_) );
NOR2X1 NOR2X1_1857 ( .gnd(gnd), .vdd(vdd), .A(_8945_), .B(_11008__bF_buf2), .Y(_11214_) );
INVX1 INVX1_726 ( .gnd(gnd), .vdd(vdd), .A(_11214_), .Y(_11215_) );
NAND2X1 NAND2X1_1482 ( .gnd(gnd), .vdd(vdd), .A(_11213_), .B(_11215_), .Y(_11216_) );
AOI21X1 AOI21X1_1902 ( .gnd(gnd), .vdd(vdd), .A(_11212_), .B(_11216_), .C(_9293__bF_buf1), .Y(_11217_) );
OAI21X1 OAI21X1_3163 ( .gnd(gnd), .vdd(vdd), .A(_11212_), .B(_11216_), .C(_11217_), .Y(_11218_) );
AND2X2 AND2X2_717 ( .gnd(gnd), .vdd(vdd), .A(_11218_), .B(_9294__bF_buf3), .Y(_11219_) );
NAND3X1 NAND3X1_589 ( .gnd(gnd), .vdd(vdd), .A(_10936_), .B(_10937_), .C(_10939_), .Y(_11220_) );
OAI21X1 OAI21X1_3164 ( .gnd(gnd), .vdd(vdd), .A(_8998_), .B(_10798__bF_buf2), .C(_11220_), .Y(_11221_) );
OAI21X1 OAI21X1_3165 ( .gnd(gnd), .vdd(vdd), .A(_10994__bF_buf4), .B(_10996__bF_buf4), .C(_9002_), .Y(_11222_) );
NOR2X1 NOR2X1_1858 ( .gnd(gnd), .vdd(vdd), .A(_9002_), .B(_11008__bF_buf1), .Y(_11223_) );
INVX1 INVX1_727 ( .gnd(gnd), .vdd(vdd), .A(_11223_), .Y(_11224_) );
NAND2X1 NAND2X1_1483 ( .gnd(gnd), .vdd(vdd), .A(_11222_), .B(_11224_), .Y(_11225_) );
XOR2X1 XOR2X1_189 ( .gnd(gnd), .vdd(vdd), .A(_11225_), .B(_11221_), .Y(_11226_) );
OAI21X1 OAI21X1_3166 ( .gnd(gnd), .vdd(vdd), .A(_11226_), .B(_9294__bF_buf2), .C(_9292__bF_buf2), .Y(_11227_) );
AOI21X1 AOI21X1_1903 ( .gnd(gnd), .vdd(vdd), .A(_11219_), .B(_11211_), .C(_11227_), .Y(_11228_) );
OAI21X1 OAI21X1_3167 ( .gnd(gnd), .vdd(vdd), .A(_8971_), .B(_10798__bF_buf1), .C(_10945_), .Y(_11229_) );
OAI21X1 OAI21X1_3168 ( .gnd(gnd), .vdd(vdd), .A(_10994__bF_buf3), .B(_10996__bF_buf3), .C(_8975_), .Y(_11230_) );
NOR2X1 NOR2X1_1859 ( .gnd(gnd), .vdd(vdd), .A(_8975_), .B(_11008__bF_buf0), .Y(_11231_) );
INVX1 INVX1_728 ( .gnd(gnd), .vdd(vdd), .A(_11231_), .Y(_11232_) );
NAND2X1 NAND2X1_1484 ( .gnd(gnd), .vdd(vdd), .A(_11230_), .B(_11232_), .Y(_11233_) );
XNOR2X1 XNOR2X1_442 ( .gnd(gnd), .vdd(vdd), .A(_11233_), .B(_11229_), .Y(_11234_) );
OAI21X1 OAI21X1_3169 ( .gnd(gnd), .vdd(vdd), .A(_11234_), .B(_9292__bF_buf1), .C(_9287__bF_buf0), .Y(_11235_) );
NAND3X1 NAND3X1_590 ( .gnd(gnd), .vdd(vdd), .A(_10952_), .B(_10953_), .C(_10955_), .Y(_11236_) );
OAI21X1 OAI21X1_3170 ( .gnd(gnd), .vdd(vdd), .A(_8841_), .B(_10798__bF_buf0), .C(_11236_), .Y(_11237_) );
OAI21X1 OAI21X1_3171 ( .gnd(gnd), .vdd(vdd), .A(_10994__bF_buf2), .B(_10996__bF_buf2), .C(_8845_), .Y(_11238_) );
INVX1 INVX1_729 ( .gnd(gnd), .vdd(vdd), .A(_11238_), .Y(_11239_) );
NOR2X1 NOR2X1_1860 ( .gnd(gnd), .vdd(vdd), .A(_8845_), .B(_11008__bF_buf4), .Y(_11240_) );
NOR2X1 NOR2X1_1861 ( .gnd(gnd), .vdd(vdd), .A(_11239_), .B(_11240_), .Y(_11241_) );
XOR2X1 XOR2X1_190 ( .gnd(gnd), .vdd(vdd), .A(_11241_), .B(_11237_), .Y(_11242_) );
AOI21X1 AOI21X1_1904 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe62_bF_buf1), .B(_11242_), .C(micro_hash_ucr_3_pipe64_bF_buf0), .Y(_11243_) );
OAI21X1 OAI21X1_3172 ( .gnd(gnd), .vdd(vdd), .A(_11228_), .B(_11235_), .C(_11243_), .Y(_11244_) );
OAI21X1 OAI21X1_3173 ( .gnd(gnd), .vdd(vdd), .A(_10959_), .B(_10798__bF_buf5), .C(_10961_), .Y(_11245_) );
INVX1 INVX1_730 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_227_), .Y(_11246_) );
OAI21X1 OAI21X1_3174 ( .gnd(gnd), .vdd(vdd), .A(_10994__bF_buf1), .B(_10996__bF_buf1), .C(_11246_), .Y(_11247_) );
NOR2X1 NOR2X1_1862 ( .gnd(gnd), .vdd(vdd), .A(_11246_), .B(_11008__bF_buf3), .Y(_11248_) );
INVX1 INVX1_731 ( .gnd(gnd), .vdd(vdd), .A(_11248_), .Y(_11249_) );
NAND2X1 NAND2X1_1485 ( .gnd(gnd), .vdd(vdd), .A(_11247_), .B(_11249_), .Y(_11250_) );
AOI21X1 AOI21X1_1905 ( .gnd(gnd), .vdd(vdd), .A(_11245_), .B(_11250_), .C(_9288__bF_buf1), .Y(_11251_) );
OAI21X1 OAI21X1_3175 ( .gnd(gnd), .vdd(vdd), .A(_11245_), .B(_11250_), .C(_11251_), .Y(_11252_) );
AOI21X1 AOI21X1_1906 ( .gnd(gnd), .vdd(vdd), .A(_11252_), .B(_11244_), .C(micro_hash_ucr_3_pipe66_bF_buf2), .Y(_11253_) );
AOI21X1 AOI21X1_1907 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe66_bF_buf1), .B(_11002_), .C(_11253_), .Y(_11254_) );
NAND3X1 NAND3X1_591 ( .gnd(gnd), .vdd(vdd), .A(_10973_), .B(_10975_), .C(_10977_), .Y(_11255_) );
OAI21X1 OAI21X1_3176 ( .gnd(gnd), .vdd(vdd), .A(_10974_), .B(_10798__bF_buf4), .C(_11255_), .Y(_11256_) );
INVX1 INVX1_732 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_243_), .Y(_11257_) );
OAI21X1 OAI21X1_3177 ( .gnd(gnd), .vdd(vdd), .A(_10994__bF_buf0), .B(_10996__bF_buf0), .C(_11257_), .Y(_11258_) );
INVX1 INVX1_733 ( .gnd(gnd), .vdd(vdd), .A(_11258_), .Y(_11259_) );
NOR2X1 NOR2X1_1863 ( .gnd(gnd), .vdd(vdd), .A(_11257_), .B(_11008__bF_buf2), .Y(_11260_) );
NOR2X1 NOR2X1_1864 ( .gnd(gnd), .vdd(vdd), .A(_11259_), .B(_11260_), .Y(_11261_) );
XOR2X1 XOR2X1_191 ( .gnd(gnd), .vdd(vdd), .A(_11261_), .B(_11256_), .Y(_11262_) );
MUX2X1 MUX2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_11254_), .B(_11262_), .S(_9282__bF_buf0), .Y(_11263_) );
NOR2X1 NOR2X1_1865 ( .gnd(gnd), .vdd(vdd), .A(_10986_), .B(_10988_), .Y(_11264_) );
INVX2 INVX2_379 ( .gnd(gnd), .vdd(vdd), .A(_11264_), .Y(_11265_) );
INVX1 INVX1_734 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_251_), .Y(_11266_) );
OAI21X1 OAI21X1_3178 ( .gnd(gnd), .vdd(vdd), .A(_10994__bF_buf4), .B(_10996__bF_buf4), .C(_11266_), .Y(_11267_) );
INVX1 INVX1_735 ( .gnd(gnd), .vdd(vdd), .A(_11267_), .Y(_11268_) );
NOR2X1 NOR2X1_1866 ( .gnd(gnd), .vdd(vdd), .A(_11266_), .B(_11008__bF_buf1), .Y(_11269_) );
NOR2X1 NOR2X1_1867 ( .gnd(gnd), .vdd(vdd), .A(_11268_), .B(_11269_), .Y(_11270_) );
AND2X2 AND2X2_718 ( .gnd(gnd), .vdd(vdd), .A(_11265_), .B(_11270_), .Y(_11271_) );
OAI21X1 OAI21X1_3179 ( .gnd(gnd), .vdd(vdd), .A(_11265_), .B(_11270_), .C(_8772_), .Y(_11272_) );
OAI22X1 OAI22X1_142 ( .gnd(gnd), .vdd(vdd), .A(_11271_), .B(_11272_), .C(_11263_), .D(_10381_), .Y(_8702__3_) );
AOI21X1 AOI21X1_1908 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_k_3_), .B(micro_hash_ucr_3_x_3_), .C(_10994__bF_buf3), .Y(_11273_) );
NOR2X1 NOR2X1_1868 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_k_4_), .B(micro_hash_ucr_3_x_4_), .Y(_11274_) );
INVX1 INVX1_736 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_k_4_), .Y(_11275_) );
INVX1 INVX1_737 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_x_4_), .Y(_11276_) );
NOR2X1 NOR2X1_1869 ( .gnd(gnd), .vdd(vdd), .A(_11275_), .B(_11276_), .Y(_11277_) );
NOR2X1 NOR2X1_1870 ( .gnd(gnd), .vdd(vdd), .A(_11274_), .B(_11277_), .Y(_11278_) );
INVX1 INVX1_738 ( .gnd(gnd), .vdd(vdd), .A(_11278_), .Y(_11279_) );
NOR2X1 NOR2X1_1871 ( .gnd(gnd), .vdd(vdd), .A(_11279_), .B(_11273_), .Y(_11280_) );
INVX1 INVX1_739 ( .gnd(gnd), .vdd(vdd), .A(_11280_), .Y(_11281_) );
OAI21X1 OAI21X1_3180 ( .gnd(gnd), .vdd(vdd), .A(_11274_), .B(_11277_), .C(_11273_), .Y(_11282_) );
NAND2X1 NAND2X1_1486 ( .gnd(gnd), .vdd(vdd), .A(_11282_), .B(_11281_), .Y(_11283_) );
XNOR2X1 XNOR2X1_443 ( .gnd(gnd), .vdd(vdd), .A(_11283__bF_buf5), .B(micro_hash_ucr_3_Wx_36_), .Y(_11284_) );
INVX1 INVX1_740 ( .gnd(gnd), .vdd(vdd), .A(_11284_), .Y(_11285_) );
AOI21X1 AOI21X1_1909 ( .gnd(gnd), .vdd(vdd), .A(_11043_), .B(_11041_), .C(_11044_), .Y(_11286_) );
AND2X2 AND2X2_719 ( .gnd(gnd), .vdd(vdd), .A(_11285_), .B(_11286_), .Y(_11287_) );
NOR2X1 NOR2X1_1872 ( .gnd(gnd), .vdd(vdd), .A(_11286_), .B(_11285_), .Y(_11288_) );
OAI21X1 OAI21X1_3181 ( .gnd(gnd), .vdd(vdd), .A(_11287_), .B(_11288_), .C(micro_hash_ucr_3_pipe16_bF_buf4), .Y(_11289_) );
INVX1 INVX1_741 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_20_), .Y(_11290_) );
XNOR2X1 XNOR2X1_444 ( .gnd(gnd), .vdd(vdd), .A(_11283__bF_buf4), .B(_11290_), .Y(_11291_) );
INVX1 INVX1_742 ( .gnd(gnd), .vdd(vdd), .A(_11031_), .Y(_11292_) );
OAI21X1 OAI21X1_3182 ( .gnd(gnd), .vdd(vdd), .A(_11028_), .B(_11292_), .C(_11033_), .Y(_11293_) );
INVX1 INVX1_743 ( .gnd(gnd), .vdd(vdd), .A(_11293_), .Y(_11294_) );
AND2X2 AND2X2_720 ( .gnd(gnd), .vdd(vdd), .A(_11291_), .B(_11294_), .Y(_11295_) );
NOR2X1 NOR2X1_1873 ( .gnd(gnd), .vdd(vdd), .A(_11294_), .B(_11291_), .Y(_11296_) );
OAI21X1 OAI21X1_3183 ( .gnd(gnd), .vdd(vdd), .A(_11295_), .B(_11296_), .C(micro_hash_ucr_3_pipe12), .Y(_11297_) );
XOR2X1 XOR2X1_192 ( .gnd(gnd), .vdd(vdd), .A(_11283__bF_buf3), .B(micro_hash_ucr_3_Wx_12_), .Y(_11298_) );
INVX1 INVX1_744 ( .gnd(gnd), .vdd(vdd), .A(_11024_), .Y(_11299_) );
AOI21X1 AOI21X1_1910 ( .gnd(gnd), .vdd(vdd), .A(_11023_), .B(_11021_), .C(_11299_), .Y(_11300_) );
AOI21X1 AOI21X1_1911 ( .gnd(gnd), .vdd(vdd), .A(_11300_), .B(_11298_), .C(_9342_), .Y(_11301_) );
OAI21X1 OAI21X1_3184 ( .gnd(gnd), .vdd(vdd), .A(_11298_), .B(_11300_), .C(_11301_), .Y(_11302_) );
XNOR2X1 XNOR2X1_445 ( .gnd(gnd), .vdd(vdd), .A(_11283__bF_buf2), .B(micro_hash_ucr_3_Wx_4_), .Y(_11303_) );
INVX1 INVX1_745 ( .gnd(gnd), .vdd(vdd), .A(_11303_), .Y(_11304_) );
OAI21X1 OAI21X1_3185 ( .gnd(gnd), .vdd(vdd), .A(_11013_), .B(_11008__bF_buf0), .C(_11012_), .Y(_11305_) );
OAI21X1 OAI21X1_3186 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_3_), .B(_10997_), .C(_11305_), .Y(_11306_) );
OR2X2 OR2X2_75 ( .gnd(gnd), .vdd(vdd), .A(_11304_), .B(_11306_), .Y(_11307_) );
NAND2X1 NAND2X1_1487 ( .gnd(gnd), .vdd(vdd), .A(_11306_), .B(_11304_), .Y(_11308_) );
AOI21X1 AOI21X1_1912 ( .gnd(gnd), .vdd(vdd), .A(_11308_), .B(_11307_), .C(_9341_), .Y(_11309_) );
INVX1 INVX1_746 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_4_), .Y(_11310_) );
NAND2X1 NAND2X1_1488 ( .gnd(gnd), .vdd(vdd), .A(H_3_20_), .B(micro_hash_ucr_3_pipe6_bF_buf1), .Y(_11311_) );
OAI21X1 OAI21X1_3187 ( .gnd(gnd), .vdd(vdd), .A(_11310_), .B(micro_hash_ucr_3_pipe6_bF_buf0), .C(_11311_), .Y(_11312_) );
OAI21X1 OAI21X1_3188 ( .gnd(gnd), .vdd(vdd), .A(_11312_), .B(micro_hash_ucr_3_pipe8), .C(_9342_), .Y(_11313_) );
OAI21X1 OAI21X1_3189 ( .gnd(gnd), .vdd(vdd), .A(_11309_), .B(_11313_), .C(_11302_), .Y(_11314_) );
OAI21X1 OAI21X1_3190 ( .gnd(gnd), .vdd(vdd), .A(_11314_), .B(micro_hash_ucr_3_pipe12), .C(_11297_), .Y(_11315_) );
XNOR2X1 XNOR2X1_446 ( .gnd(gnd), .vdd(vdd), .A(_11283__bF_buf1), .B(micro_hash_ucr_3_Wx_28_), .Y(_11316_) );
INVX1 INVX1_747 ( .gnd(gnd), .vdd(vdd), .A(_11316_), .Y(_11317_) );
AOI21X1 AOI21X1_1913 ( .gnd(gnd), .vdd(vdd), .A(_11006_), .B(_11004_), .C(_11009_), .Y(_11318_) );
NOR2X1 NOR2X1_1874 ( .gnd(gnd), .vdd(vdd), .A(_11318_), .B(_11317_), .Y(_11319_) );
INVX1 INVX1_748 ( .gnd(gnd), .vdd(vdd), .A(_11319_), .Y(_11320_) );
NAND2X1 NAND2X1_1489 ( .gnd(gnd), .vdd(vdd), .A(_11318_), .B(_11317_), .Y(_11321_) );
NAND3X1 NAND3X1_592 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe14_bF_buf0), .B(_11321_), .C(_11320_), .Y(_11322_) );
OAI21X1 OAI21X1_3191 ( .gnd(gnd), .vdd(vdd), .A(_11315_), .B(micro_hash_ucr_3_pipe14_bF_buf3), .C(_11322_), .Y(_11323_) );
OAI21X1 OAI21X1_3192 ( .gnd(gnd), .vdd(vdd), .A(_11323_), .B(micro_hash_ucr_3_pipe16_bF_buf3), .C(_11289_), .Y(_11324_) );
XNOR2X1 XNOR2X1_447 ( .gnd(gnd), .vdd(vdd), .A(_11283__bF_buf0), .B(micro_hash_ucr_3_Wx_44_), .Y(_11325_) );
INVX1 INVX1_749 ( .gnd(gnd), .vdd(vdd), .A(_11325_), .Y(_11326_) );
AOI21X1 AOI21X1_1914 ( .gnd(gnd), .vdd(vdd), .A(_11052_), .B(_11050_), .C(_11053_), .Y(_11327_) );
NOR2X1 NOR2X1_1875 ( .gnd(gnd), .vdd(vdd), .A(_11327_), .B(_11326_), .Y(_11328_) );
INVX1 INVX1_750 ( .gnd(gnd), .vdd(vdd), .A(_11328_), .Y(_11329_) );
NAND2X1 NAND2X1_1490 ( .gnd(gnd), .vdd(vdd), .A(_11327_), .B(_11326_), .Y(_11330_) );
NAND3X1 NAND3X1_593 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe18_bF_buf4), .B(_11330_), .C(_11329_), .Y(_11331_) );
OAI21X1 OAI21X1_3193 ( .gnd(gnd), .vdd(vdd), .A(_11324_), .B(micro_hash_ucr_3_pipe18_bF_buf3), .C(_11331_), .Y(_11332_) );
XNOR2X1 XNOR2X1_448 ( .gnd(gnd), .vdd(vdd), .A(_11283__bF_buf5), .B(micro_hash_ucr_3_Wx_52_), .Y(_11333_) );
INVX1 INVX1_751 ( .gnd(gnd), .vdd(vdd), .A(_11333_), .Y(_11334_) );
AOI21X1 AOI21X1_1915 ( .gnd(gnd), .vdd(vdd), .A(_11063_), .B(_11061_), .C(_11064_), .Y(_11335_) );
NAND2X1 NAND2X1_1491 ( .gnd(gnd), .vdd(vdd), .A(_11335_), .B(_11334_), .Y(_11336_) );
NOR2X1 NOR2X1_1876 ( .gnd(gnd), .vdd(vdd), .A(_11335_), .B(_11334_), .Y(_11337_) );
INVX1 INVX1_752 ( .gnd(gnd), .vdd(vdd), .A(_11337_), .Y(_11338_) );
NAND2X1 NAND2X1_1492 ( .gnd(gnd), .vdd(vdd), .A(_11336_), .B(_11338_), .Y(_11339_) );
AOI21X1 AOI21X1_1916 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe20_bF_buf4), .B(_11339_), .C(micro_hash_ucr_3_pipe22_bF_buf4), .Y(_11340_) );
OAI21X1 OAI21X1_3194 ( .gnd(gnd), .vdd(vdd), .A(_11332_), .B(micro_hash_ucr_3_pipe20_bF_buf3), .C(_11340_), .Y(_11341_) );
XNOR2X1 XNOR2X1_449 ( .gnd(gnd), .vdd(vdd), .A(_11283__bF_buf4), .B(micro_hash_ucr_3_Wx_60_), .Y(_11342_) );
INVX1 INVX1_753 ( .gnd(gnd), .vdd(vdd), .A(_11072_), .Y(_11343_) );
OAI21X1 OAI21X1_3195 ( .gnd(gnd), .vdd(vdd), .A(_11069_), .B(_11071_), .C(_11343_), .Y(_11344_) );
NAND2X1 NAND2X1_1493 ( .gnd(gnd), .vdd(vdd), .A(_11344_), .B(_11342_), .Y(_11345_) );
INVX1 INVX1_754 ( .gnd(gnd), .vdd(vdd), .A(_11345_), .Y(_11346_) );
OAI21X1 OAI21X1_3196 ( .gnd(gnd), .vdd(vdd), .A(_11342_), .B(_11344_), .C(micro_hash_ucr_3_pipe22_bF_buf3), .Y(_11347_) );
OAI21X1 OAI21X1_3197 ( .gnd(gnd), .vdd(vdd), .A(_11346_), .B(_11347_), .C(_11341_), .Y(_11348_) );
XNOR2X1 XNOR2X1_450 ( .gnd(gnd), .vdd(vdd), .A(_11283__bF_buf3), .B(micro_hash_ucr_3_Wx_68_), .Y(_11349_) );
INVX1 INVX1_755 ( .gnd(gnd), .vdd(vdd), .A(_11349_), .Y(_11350_) );
AOI21X1 AOI21X1_1917 ( .gnd(gnd), .vdd(vdd), .A(_11079_), .B(_11078_), .C(_11080_), .Y(_11351_) );
AND2X2 AND2X2_721 ( .gnd(gnd), .vdd(vdd), .A(_11350_), .B(_11351_), .Y(_11352_) );
NOR2X1 NOR2X1_1877 ( .gnd(gnd), .vdd(vdd), .A(_11351_), .B(_11350_), .Y(_11353_) );
OAI21X1 OAI21X1_3198 ( .gnd(gnd), .vdd(vdd), .A(_11352_), .B(_11353_), .C(micro_hash_ucr_3_pipe24_bF_buf4), .Y(_11354_) );
OAI21X1 OAI21X1_3199 ( .gnd(gnd), .vdd(vdd), .A(_11348_), .B(micro_hash_ucr_3_pipe24_bF_buf3), .C(_11354_), .Y(_11355_) );
NOR2X1 NOR2X1_1878 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe26_bF_buf2), .B(_11355_), .Y(_11356_) );
XNOR2X1 XNOR2X1_451 ( .gnd(gnd), .vdd(vdd), .A(_11283__bF_buf2), .B(micro_hash_ucr_3_Wx_76_), .Y(_11357_) );
INVX1 INVX1_756 ( .gnd(gnd), .vdd(vdd), .A(_11357_), .Y(_11358_) );
AOI21X1 AOI21X1_1918 ( .gnd(gnd), .vdd(vdd), .A(_11087_), .B(_11086_), .C(_11088_), .Y(_11359_) );
NOR2X1 NOR2X1_1879 ( .gnd(gnd), .vdd(vdd), .A(_11359_), .B(_11358_), .Y(_11360_) );
INVX1 INVX1_757 ( .gnd(gnd), .vdd(vdd), .A(_11360_), .Y(_11361_) );
AOI21X1 AOI21X1_1919 ( .gnd(gnd), .vdd(vdd), .A(_11359_), .B(_11358_), .C(_9323__bF_buf1), .Y(_11362_) );
AOI21X1 AOI21X1_1920 ( .gnd(gnd), .vdd(vdd), .A(_11361_), .B(_11362_), .C(_11356_), .Y(_11363_) );
XNOR2X1 XNOR2X1_452 ( .gnd(gnd), .vdd(vdd), .A(_11283__bF_buf1), .B(micro_hash_ucr_3_Wx_84_), .Y(_11364_) );
INVX1 INVX1_758 ( .gnd(gnd), .vdd(vdd), .A(_11364_), .Y(_11365_) );
AOI21X1 AOI21X1_1921 ( .gnd(gnd), .vdd(vdd), .A(_11098_), .B(_11097_), .C(_11099_), .Y(_11366_) );
NAND2X1 NAND2X1_1494 ( .gnd(gnd), .vdd(vdd), .A(_11366_), .B(_11365_), .Y(_11367_) );
NOR2X1 NOR2X1_1880 ( .gnd(gnd), .vdd(vdd), .A(_11366_), .B(_11365_), .Y(_11368_) );
INVX1 INVX1_759 ( .gnd(gnd), .vdd(vdd), .A(_11368_), .Y(_11369_) );
NAND3X1 NAND3X1_594 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe28_bF_buf2), .B(_11367_), .C(_11369_), .Y(_11370_) );
OAI21X1 OAI21X1_3200 ( .gnd(gnd), .vdd(vdd), .A(_11363_), .B(micro_hash_ucr_3_pipe28_bF_buf1), .C(_11370_), .Y(_11371_) );
XNOR2X1 XNOR2X1_453 ( .gnd(gnd), .vdd(vdd), .A(_11283__bF_buf0), .B(micro_hash_ucr_3_Wx_92_), .Y(_11372_) );
INVX1 INVX1_760 ( .gnd(gnd), .vdd(vdd), .A(_11372_), .Y(_11373_) );
AOI21X1 AOI21X1_1922 ( .gnd(gnd), .vdd(vdd), .A(_11105_), .B(_11104_), .C(_11107_), .Y(_11374_) );
NOR2X1 NOR2X1_1881 ( .gnd(gnd), .vdd(vdd), .A(_11374_), .B(_11373_), .Y(_11375_) );
INVX1 INVX1_761 ( .gnd(gnd), .vdd(vdd), .A(_11375_), .Y(_11376_) );
AOI21X1 AOI21X1_1923 ( .gnd(gnd), .vdd(vdd), .A(_11374_), .B(_11373_), .C(_9322__bF_buf0), .Y(_11377_) );
AOI22X1 AOI22X1_79 ( .gnd(gnd), .vdd(vdd), .A(_11376_), .B(_11377_), .C(_11371_), .D(_9322__bF_buf3), .Y(_11378_) );
XNOR2X1 XNOR2X1_454 ( .gnd(gnd), .vdd(vdd), .A(_11283__bF_buf5), .B(micro_hash_ucr_3_Wx_100_), .Y(_11379_) );
INVX1 INVX1_762 ( .gnd(gnd), .vdd(vdd), .A(_11379_), .Y(_11380_) );
AOI21X1 AOI21X1_1924 ( .gnd(gnd), .vdd(vdd), .A(_11114_), .B(_11113_), .C(_11115_), .Y(_11381_) );
NAND2X1 NAND2X1_1495 ( .gnd(gnd), .vdd(vdd), .A(_11381_), .B(_11380_), .Y(_11382_) );
NOR2X1 NOR2X1_1882 ( .gnd(gnd), .vdd(vdd), .A(_11381_), .B(_11380_), .Y(_11383_) );
NOR2X1 NOR2X1_1883 ( .gnd(gnd), .vdd(vdd), .A(_9317__bF_buf0), .B(_11383_), .Y(_11384_) );
AOI21X1 AOI21X1_1925 ( .gnd(gnd), .vdd(vdd), .A(_11382_), .B(_11384_), .C(micro_hash_ucr_3_pipe34_bF_buf2), .Y(_11385_) );
OAI21X1 OAI21X1_3201 ( .gnd(gnd), .vdd(vdd), .A(_11378_), .B(micro_hash_ucr_3_pipe32_bF_buf0), .C(_11385_), .Y(_11386_) );
XNOR2X1 XNOR2X1_455 ( .gnd(gnd), .vdd(vdd), .A(_11283__bF_buf4), .B(micro_hash_ucr_3_Wx_108_), .Y(_11387_) );
INVX1 INVX1_763 ( .gnd(gnd), .vdd(vdd), .A(_11387_), .Y(_11388_) );
AOI21X1 AOI21X1_1926 ( .gnd(gnd), .vdd(vdd), .A(_11122_), .B(_11121_), .C(_11123_), .Y(_11389_) );
AND2X2 AND2X2_722 ( .gnd(gnd), .vdd(vdd), .A(_11388_), .B(_11389_), .Y(_11390_) );
NOR2X1 NOR2X1_1884 ( .gnd(gnd), .vdd(vdd), .A(_11389_), .B(_11388_), .Y(_11391_) );
OAI21X1 OAI21X1_3202 ( .gnd(gnd), .vdd(vdd), .A(_11390_), .B(_11391_), .C(micro_hash_ucr_3_pipe34_bF_buf1), .Y(_11392_) );
AOI21X1 AOI21X1_1927 ( .gnd(gnd), .vdd(vdd), .A(_11392_), .B(_11386_), .C(micro_hash_ucr_3_pipe36_bF_buf1), .Y(_11393_) );
XNOR2X1 XNOR2X1_456 ( .gnd(gnd), .vdd(vdd), .A(_11283__bF_buf3), .B(micro_hash_ucr_3_Wx_116_), .Y(_11394_) );
INVX1 INVX1_764 ( .gnd(gnd), .vdd(vdd), .A(_11394_), .Y(_11395_) );
AOI21X1 AOI21X1_1928 ( .gnd(gnd), .vdd(vdd), .A(_11131_), .B(_11130_), .C(_11132_), .Y(_11396_) );
NOR2X1 NOR2X1_1885 ( .gnd(gnd), .vdd(vdd), .A(_11396_), .B(_11395_), .Y(_11397_) );
INVX1 INVX1_765 ( .gnd(gnd), .vdd(vdd), .A(_11397_), .Y(_11398_) );
NAND2X1 NAND2X1_1496 ( .gnd(gnd), .vdd(vdd), .A(_11396_), .B(_11395_), .Y(_11399_) );
AOI21X1 AOI21X1_1929 ( .gnd(gnd), .vdd(vdd), .A(_11399_), .B(_11398_), .C(_9316__bF_buf3), .Y(_11400_) );
OAI21X1 OAI21X1_3203 ( .gnd(gnd), .vdd(vdd), .A(_11393_), .B(_11400_), .C(_9311__bF_buf4), .Y(_11401_) );
XNOR2X1 XNOR2X1_457 ( .gnd(gnd), .vdd(vdd), .A(_11283__bF_buf2), .B(_8978_), .Y(_11402_) );
AOI21X1 AOI21X1_1930 ( .gnd(gnd), .vdd(vdd), .A(_11138_), .B(_11137_), .C(_11139_), .Y(_11403_) );
AND2X2 AND2X2_723 ( .gnd(gnd), .vdd(vdd), .A(_11403_), .B(_11402_), .Y(_11404_) );
NOR2X1 NOR2X1_1886 ( .gnd(gnd), .vdd(vdd), .A(_11402_), .B(_11403_), .Y(_11405_) );
OAI21X1 OAI21X1_3204 ( .gnd(gnd), .vdd(vdd), .A(_11404_), .B(_11405_), .C(micro_hash_ucr_3_pipe38_bF_buf0), .Y(_11406_) );
AOI21X1 AOI21X1_1931 ( .gnd(gnd), .vdd(vdd), .A(_11406_), .B(_11401_), .C(micro_hash_ucr_3_pipe40_bF_buf1), .Y(_11407_) );
XNOR2X1 XNOR2X1_458 ( .gnd(gnd), .vdd(vdd), .A(_11283__bF_buf1), .B(micro_hash_ucr_3_Wx_132_), .Y(_11408_) );
INVX1 INVX1_766 ( .gnd(gnd), .vdd(vdd), .A(_11408_), .Y(_11409_) );
AOI21X1 AOI21X1_1932 ( .gnd(gnd), .vdd(vdd), .A(_11147_), .B(_11146_), .C(_11148_), .Y(_11410_) );
NAND2X1 NAND2X1_1497 ( .gnd(gnd), .vdd(vdd), .A(_11410_), .B(_11409_), .Y(_11411_) );
NOR2X1 NOR2X1_1887 ( .gnd(gnd), .vdd(vdd), .A(_11410_), .B(_11409_), .Y(_11412_) );
INVX1 INVX1_767 ( .gnd(gnd), .vdd(vdd), .A(_11412_), .Y(_11413_) );
AOI21X1 AOI21X1_1933 ( .gnd(gnd), .vdd(vdd), .A(_11411_), .B(_11413_), .C(_9312__bF_buf3), .Y(_11414_) );
OAI21X1 OAI21X1_3205 ( .gnd(gnd), .vdd(vdd), .A(_11407_), .B(_11414_), .C(_9310__bF_buf4), .Y(_11415_) );
XNOR2X1 XNOR2X1_459 ( .gnd(gnd), .vdd(vdd), .A(_11283__bF_buf0), .B(micro_hash_ucr_3_Wx_140_), .Y(_11416_) );
INVX1 INVX1_768 ( .gnd(gnd), .vdd(vdd), .A(_11416_), .Y(_11417_) );
AOI21X1 AOI21X1_1934 ( .gnd(gnd), .vdd(vdd), .A(_11155_), .B(_11154_), .C(_11156_), .Y(_11418_) );
AND2X2 AND2X2_724 ( .gnd(gnd), .vdd(vdd), .A(_11417_), .B(_11418_), .Y(_11419_) );
NOR2X1 NOR2X1_1888 ( .gnd(gnd), .vdd(vdd), .A(_11418_), .B(_11417_), .Y(_11420_) );
OAI21X1 OAI21X1_3206 ( .gnd(gnd), .vdd(vdd), .A(_11419_), .B(_11420_), .C(micro_hash_ucr_3_pipe42_bF_buf0), .Y(_11421_) );
NAND3X1 NAND3X1_595 ( .gnd(gnd), .vdd(vdd), .A(_9305__bF_buf1), .B(_11421_), .C(_11415_), .Y(_11422_) );
XNOR2X1 XNOR2X1_460 ( .gnd(gnd), .vdd(vdd), .A(_11283__bF_buf5), .B(micro_hash_ucr_3_Wx_148_), .Y(_11423_) );
INVX1 INVX1_769 ( .gnd(gnd), .vdd(vdd), .A(_11423_), .Y(_11424_) );
AOI21X1 AOI21X1_1935 ( .gnd(gnd), .vdd(vdd), .A(_11164_), .B(_11163_), .C(_11165_), .Y(_11425_) );
NOR2X1 NOR2X1_1889 ( .gnd(gnd), .vdd(vdd), .A(_11425_), .B(_11424_), .Y(_11426_) );
INVX1 INVX1_770 ( .gnd(gnd), .vdd(vdd), .A(_11426_), .Y(_11427_) );
NAND2X1 NAND2X1_1498 ( .gnd(gnd), .vdd(vdd), .A(_11425_), .B(_11424_), .Y(_11428_) );
NAND2X1 NAND2X1_1499 ( .gnd(gnd), .vdd(vdd), .A(_11428_), .B(_11427_), .Y(_11429_) );
OAI21X1 OAI21X1_3207 ( .gnd(gnd), .vdd(vdd), .A(_9305__bF_buf0), .B(_11429_), .C(_11422_), .Y(_11430_) );
NOR2X1 NOR2X1_1890 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe46_bF_buf1), .B(_11430_), .Y(_11431_) );
XNOR2X1 XNOR2X1_461 ( .gnd(gnd), .vdd(vdd), .A(_11283__bF_buf4), .B(micro_hash_ucr_3_Wx_156_), .Y(_11432_) );
INVX1 INVX1_771 ( .gnd(gnd), .vdd(vdd), .A(_11432_), .Y(_11433_) );
AOI21X1 AOI21X1_1936 ( .gnd(gnd), .vdd(vdd), .A(_11171_), .B(_11170_), .C(_11173_), .Y(_11434_) );
NAND2X1 NAND2X1_1500 ( .gnd(gnd), .vdd(vdd), .A(_11434_), .B(_11433_), .Y(_11435_) );
NOR2X1 NOR2X1_1891 ( .gnd(gnd), .vdd(vdd), .A(_11434_), .B(_11433_), .Y(_11436_) );
INVX1 INVX1_772 ( .gnd(gnd), .vdd(vdd), .A(_11436_), .Y(_11437_) );
AOI21X1 AOI21X1_1937 ( .gnd(gnd), .vdd(vdd), .A(_11435_), .B(_11437_), .C(_9306__bF_buf2), .Y(_11438_) );
OAI21X1 OAI21X1_3208 ( .gnd(gnd), .vdd(vdd), .A(_11431_), .B(_11438_), .C(_9304__bF_buf1), .Y(_11439_) );
XNOR2X1 XNOR2X1_462 ( .gnd(gnd), .vdd(vdd), .A(_11283__bF_buf3), .B(micro_hash_ucr_3_Wx_164_), .Y(_11440_) );
INVX1 INVX1_773 ( .gnd(gnd), .vdd(vdd), .A(_11440_), .Y(_11441_) );
AOI21X1 AOI21X1_1938 ( .gnd(gnd), .vdd(vdd), .A(_11180_), .B(_11179_), .C(_11181_), .Y(_11442_) );
AND2X2 AND2X2_725 ( .gnd(gnd), .vdd(vdd), .A(_11441_), .B(_11442_), .Y(_11443_) );
NOR2X1 NOR2X1_1892 ( .gnd(gnd), .vdd(vdd), .A(_11442_), .B(_11441_), .Y(_11444_) );
OAI21X1 OAI21X1_3209 ( .gnd(gnd), .vdd(vdd), .A(_11443_), .B(_11444_), .C(micro_hash_ucr_3_pipe48_bF_buf2), .Y(_11445_) );
NAND3X1 NAND3X1_596 ( .gnd(gnd), .vdd(vdd), .A(_9299__bF_buf0), .B(_11445_), .C(_11439_), .Y(_11446_) );
XNOR2X1 XNOR2X1_463 ( .gnd(gnd), .vdd(vdd), .A(_11283__bF_buf2), .B(micro_hash_ucr_3_Wx_172_), .Y(_11447_) );
INVX1 INVX1_774 ( .gnd(gnd), .vdd(vdd), .A(_11447_), .Y(_11448_) );
AOI21X1 AOI21X1_1939 ( .gnd(gnd), .vdd(vdd), .A(_11189_), .B(_11188_), .C(_11190_), .Y(_11449_) );
NOR2X1 NOR2X1_1893 ( .gnd(gnd), .vdd(vdd), .A(_11449_), .B(_11448_), .Y(_11450_) );
INVX1 INVX1_775 ( .gnd(gnd), .vdd(vdd), .A(_11450_), .Y(_11451_) );
NAND2X1 NAND2X1_1501 ( .gnd(gnd), .vdd(vdd), .A(_11449_), .B(_11448_), .Y(_11452_) );
NAND2X1 NAND2X1_1502 ( .gnd(gnd), .vdd(vdd), .A(_11452_), .B(_11451_), .Y(_11453_) );
OAI21X1 OAI21X1_3210 ( .gnd(gnd), .vdd(vdd), .A(_9299__bF_buf3), .B(_11453_), .C(_11446_), .Y(_11454_) );
XNOR2X1 XNOR2X1_464 ( .gnd(gnd), .vdd(vdd), .A(_11283__bF_buf1), .B(_9085_), .Y(_11455_) );
AOI21X1 AOI21X1_1940 ( .gnd(gnd), .vdd(vdd), .A(_11197_), .B(_11196_), .C(_11198_), .Y(_11456_) );
AND2X2 AND2X2_726 ( .gnd(gnd), .vdd(vdd), .A(_11455_), .B(_11456_), .Y(_11457_) );
NOR2X1 NOR2X1_1894 ( .gnd(gnd), .vdd(vdd), .A(_11456_), .B(_11455_), .Y(_11458_) );
OAI21X1 OAI21X1_3211 ( .gnd(gnd), .vdd(vdd), .A(_11457_), .B(_11458_), .C(micro_hash_ucr_3_pipe52_bF_buf1), .Y(_11459_) );
OAI21X1 OAI21X1_3212 ( .gnd(gnd), .vdd(vdd), .A(_11454_), .B(micro_hash_ucr_3_pipe52_bF_buf0), .C(_11459_), .Y(_11460_) );
NAND2X1 NAND2X1_1503 ( .gnd(gnd), .vdd(vdd), .A(_9298__bF_buf3), .B(_11460_), .Y(_11461_) );
XNOR2X1 XNOR2X1_465 ( .gnd(gnd), .vdd(vdd), .A(_11283__bF_buf0), .B(micro_hash_ucr_3_Wx_188_), .Y(_11462_) );
INVX1 INVX1_776 ( .gnd(gnd), .vdd(vdd), .A(_11462_), .Y(_11463_) );
AOI21X1 AOI21X1_1941 ( .gnd(gnd), .vdd(vdd), .A(_11205_), .B(_11204_), .C(_11207_), .Y(_11464_) );
AND2X2 AND2X2_727 ( .gnd(gnd), .vdd(vdd), .A(_11463_), .B(_11464_), .Y(_11465_) );
NOR2X1 NOR2X1_1895 ( .gnd(gnd), .vdd(vdd), .A(_11464_), .B(_11463_), .Y(_11466_) );
OAI21X1 OAI21X1_3213 ( .gnd(gnd), .vdd(vdd), .A(_11465_), .B(_11466_), .C(micro_hash_ucr_3_pipe54_bF_buf1), .Y(_11467_) );
AND2X2 AND2X2_728 ( .gnd(gnd), .vdd(vdd), .A(_11467_), .B(_9293__bF_buf0), .Y(_11468_) );
XNOR2X1 XNOR2X1_466 ( .gnd(gnd), .vdd(vdd), .A(_11283__bF_buf5), .B(micro_hash_ucr_3_Wx_196_), .Y(_11469_) );
INVX1 INVX1_777 ( .gnd(gnd), .vdd(vdd), .A(_11469_), .Y(_11470_) );
AOI21X1 AOI21X1_1942 ( .gnd(gnd), .vdd(vdd), .A(_11213_), .B(_11212_), .C(_11214_), .Y(_11471_) );
NOR2X1 NOR2X1_1896 ( .gnd(gnd), .vdd(vdd), .A(_11471_), .B(_11470_), .Y(_11472_) );
INVX1 INVX1_778 ( .gnd(gnd), .vdd(vdd), .A(_11472_), .Y(_11473_) );
AOI21X1 AOI21X1_1943 ( .gnd(gnd), .vdd(vdd), .A(_11471_), .B(_11470_), .C(_9293__bF_buf3), .Y(_11474_) );
AOI22X1 AOI22X1_80 ( .gnd(gnd), .vdd(vdd), .A(_11473_), .B(_11474_), .C(_11461_), .D(_11468_), .Y(_11475_) );
XNOR2X1 XNOR2X1_467 ( .gnd(gnd), .vdd(vdd), .A(_11283__bF_buf4), .B(micro_hash_ucr_3_Wx_204_), .Y(_11476_) );
INVX1 INVX1_779 ( .gnd(gnd), .vdd(vdd), .A(_11476_), .Y(_11477_) );
AOI21X1 AOI21X1_1944 ( .gnd(gnd), .vdd(vdd), .A(_11222_), .B(_11221_), .C(_11223_), .Y(_11478_) );
NAND2X1 NAND2X1_1504 ( .gnd(gnd), .vdd(vdd), .A(_11478_), .B(_11477_), .Y(_11479_) );
NOR2X1 NOR2X1_1897 ( .gnd(gnd), .vdd(vdd), .A(_11478_), .B(_11477_), .Y(_11480_) );
NOR2X1 NOR2X1_1898 ( .gnd(gnd), .vdd(vdd), .A(_9294__bF_buf1), .B(_11480_), .Y(_11481_) );
AOI21X1 AOI21X1_1945 ( .gnd(gnd), .vdd(vdd), .A(_11479_), .B(_11481_), .C(micro_hash_ucr_3_pipe60_bF_buf4), .Y(_11482_) );
OAI21X1 OAI21X1_3214 ( .gnd(gnd), .vdd(vdd), .A(_11475_), .B(micro_hash_ucr_3_pipe58_bF_buf2), .C(_11482_), .Y(_11483_) );
XNOR2X1 XNOR2X1_468 ( .gnd(gnd), .vdd(vdd), .A(_11283__bF_buf3), .B(micro_hash_ucr_3_Wx_212_), .Y(_11484_) );
INVX1 INVX1_780 ( .gnd(gnd), .vdd(vdd), .A(_11484_), .Y(_11485_) );
AOI21X1 AOI21X1_1946 ( .gnd(gnd), .vdd(vdd), .A(_11230_), .B(_11229_), .C(_11231_), .Y(_11486_) );
AND2X2 AND2X2_729 ( .gnd(gnd), .vdd(vdd), .A(_11485_), .B(_11486_), .Y(_11487_) );
NOR2X1 NOR2X1_1899 ( .gnd(gnd), .vdd(vdd), .A(_11486_), .B(_11485_), .Y(_11488_) );
OAI21X1 OAI21X1_3215 ( .gnd(gnd), .vdd(vdd), .A(_11487_), .B(_11488_), .C(micro_hash_ucr_3_pipe60_bF_buf3), .Y(_11489_) );
NAND3X1 NAND3X1_597 ( .gnd(gnd), .vdd(vdd), .A(_9287__bF_buf4), .B(_11489_), .C(_11483_), .Y(_11490_) );
XNOR2X1 XNOR2X1_469 ( .gnd(gnd), .vdd(vdd), .A(_11283__bF_buf2), .B(micro_hash_ucr_3_Wx_220_), .Y(_11491_) );
INVX1 INVX1_781 ( .gnd(gnd), .vdd(vdd), .A(_11491_), .Y(_11492_) );
AOI21X1 AOI21X1_1947 ( .gnd(gnd), .vdd(vdd), .A(_11238_), .B(_11237_), .C(_11240_), .Y(_11493_) );
NOR2X1 NOR2X1_1900 ( .gnd(gnd), .vdd(vdd), .A(_11493_), .B(_11492_), .Y(_11494_) );
NAND2X1 NAND2X1_1505 ( .gnd(gnd), .vdd(vdd), .A(_11493_), .B(_11492_), .Y(_11495_) );
NAND2X1 NAND2X1_1506 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe62_bF_buf0), .B(_11495_), .Y(_11496_) );
OAI21X1 OAI21X1_3216 ( .gnd(gnd), .vdd(vdd), .A(_11494_), .B(_11496_), .C(_11490_), .Y(_11497_) );
XNOR2X1 XNOR2X1_470 ( .gnd(gnd), .vdd(vdd), .A(_11283__bF_buf1), .B(micro_hash_ucr_3_Wx_228_), .Y(_11498_) );
INVX2 INVX2_380 ( .gnd(gnd), .vdd(vdd), .A(_11498_), .Y(_11499_) );
AOI21X1 AOI21X1_1948 ( .gnd(gnd), .vdd(vdd), .A(_11247_), .B(_11245_), .C(_11248_), .Y(_11500_) );
AND2X2 AND2X2_730 ( .gnd(gnd), .vdd(vdd), .A(_11499_), .B(_11500_), .Y(_11501_) );
OAI21X1 OAI21X1_3217 ( .gnd(gnd), .vdd(vdd), .A(_11499_), .B(_11500_), .C(micro_hash_ucr_3_pipe64_bF_buf4), .Y(_11502_) );
OAI21X1 OAI21X1_3218 ( .gnd(gnd), .vdd(vdd), .A(_11501_), .B(_11502_), .C(_9286__bF_buf3), .Y(_11503_) );
AOI21X1 AOI21X1_1949 ( .gnd(gnd), .vdd(vdd), .A(_9288__bF_buf0), .B(_11497_), .C(_11503_), .Y(_11504_) );
XNOR2X1 XNOR2X1_471 ( .gnd(gnd), .vdd(vdd), .A(_11283__bF_buf0), .B(micro_hash_ucr_3_Wx_236_), .Y(_11505_) );
INVX1 INVX1_782 ( .gnd(gnd), .vdd(vdd), .A(_10991_), .Y(_11506_) );
OAI21X1 OAI21X1_3219 ( .gnd(gnd), .vdd(vdd), .A(_11506_), .B(_10998_), .C(_11000_), .Y(_11507_) );
OR2X2 OR2X2_76 ( .gnd(gnd), .vdd(vdd), .A(_11505_), .B(_11507_), .Y(_11508_) );
NAND2X1 NAND2X1_1507 ( .gnd(gnd), .vdd(vdd), .A(_11507_), .B(_11505_), .Y(_11509_) );
AOI21X1 AOI21X1_1950 ( .gnd(gnd), .vdd(vdd), .A(_11509_), .B(_11508_), .C(_9286__bF_buf2), .Y(_11510_) );
OAI21X1 OAI21X1_3220 ( .gnd(gnd), .vdd(vdd), .A(_11504_), .B(_11510_), .C(_9282__bF_buf4), .Y(_11511_) );
XNOR2X1 XNOR2X1_472 ( .gnd(gnd), .vdd(vdd), .A(_11283__bF_buf5), .B(micro_hash_ucr_3_Wx_244_), .Y(_11512_) );
INVX1 INVX1_783 ( .gnd(gnd), .vdd(vdd), .A(_11512_), .Y(_11513_) );
AOI21X1 AOI21X1_1951 ( .gnd(gnd), .vdd(vdd), .A(_11258_), .B(_11256_), .C(_11260_), .Y(_11514_) );
AND2X2 AND2X2_731 ( .gnd(gnd), .vdd(vdd), .A(_11513_), .B(_11514_), .Y(_11515_) );
NOR2X1 NOR2X1_1901 ( .gnd(gnd), .vdd(vdd), .A(_11514_), .B(_11513_), .Y(_11516_) );
OAI21X1 OAI21X1_3221 ( .gnd(gnd), .vdd(vdd), .A(_11515_), .B(_11516_), .C(micro_hash_ucr_3_pipe68_bF_buf0), .Y(_11517_) );
NAND2X1 NAND2X1_1508 ( .gnd(gnd), .vdd(vdd), .A(_11517_), .B(_11511_), .Y(_11518_) );
XNOR2X1 XNOR2X1_473 ( .gnd(gnd), .vdd(vdd), .A(_11283__bF_buf4), .B(micro_hash_ucr_3_Wx_252_), .Y(_11519_) );
INVX2 INVX2_381 ( .gnd(gnd), .vdd(vdd), .A(_11519_), .Y(_11520_) );
AOI21X1 AOI21X1_1952 ( .gnd(gnd), .vdd(vdd), .A(_11267_), .B(_11265_), .C(_11269_), .Y(_11521_) );
AOI21X1 AOI21X1_1953 ( .gnd(gnd), .vdd(vdd), .A(_11521_), .B(_11520_), .C(_8800__bF_buf3), .Y(_11522_) );
OAI21X1 OAI21X1_3222 ( .gnd(gnd), .vdd(vdd), .A(_11520_), .B(_11521_), .C(_11522_), .Y(_11523_) );
AOI22X1 AOI22X1_81 ( .gnd(gnd), .vdd(vdd), .A(_10381_), .B(_11523_), .C(_11518_), .D(_9283__bF_buf2), .Y(_8702__4_) );
INVX4 INVX4_153 ( .gnd(gnd), .vdd(vdd), .A(_8772_), .Y(_11524_) );
INVX1 INVX1_784 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_236_), .Y(_11525_) );
OAI21X1 OAI21X1_3223 ( .gnd(gnd), .vdd(vdd), .A(_11525_), .B(_11283__bF_buf3), .C(_11509_), .Y(_11526_) );
INVX2 INVX2_382 ( .gnd(gnd), .vdd(vdd), .A(_11526_), .Y(_11527_) );
INVX2 INVX2_383 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_x_5_), .Y(_11528_) );
NAND2X1 NAND2X1_1509 ( .gnd(gnd), .vdd(vdd), .A(_10255_), .B(_11528_), .Y(_11529_) );
NOR2X1 NOR2X1_1902 ( .gnd(gnd), .vdd(vdd), .A(_10255_), .B(_11528_), .Y(_11530_) );
INVX1 INVX1_785 ( .gnd(gnd), .vdd(vdd), .A(_11530_), .Y(_11531_) );
AND2X2 AND2X2_732 ( .gnd(gnd), .vdd(vdd), .A(_11531_), .B(_11529_), .Y(_11532_) );
OAI21X1 OAI21X1_3224 ( .gnd(gnd), .vdd(vdd), .A(_11280_), .B(_11277_), .C(_11532_), .Y(_11533_) );
INVX8 INVX8_282 ( .gnd(gnd), .vdd(vdd), .A(_11533_), .Y(_11534_) );
OAI21X1 OAI21X1_3225 ( .gnd(gnd), .vdd(vdd), .A(_11275_), .B(_11276_), .C(_11281_), .Y(_11535_) );
NOR2X1 NOR2X1_1903 ( .gnd(gnd), .vdd(vdd), .A(_11532_), .B(_11535_), .Y(_11536_) );
NOR2X1 NOR2X1_1904 ( .gnd(gnd), .vdd(vdd), .A(_11534__bF_buf3), .B(_11536__bF_buf3), .Y(_11537_) );
NOR2X1 NOR2X1_1905 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_237_), .B(_11537__bF_buf4), .Y(_11538_) );
INVX1 INVX1_786 ( .gnd(gnd), .vdd(vdd), .A(_11538_), .Y(_11539_) );
NAND2X1 NAND2X1_1510 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_237_), .B(_11537__bF_buf3), .Y(_11540_) );
NAND2X1 NAND2X1_1511 ( .gnd(gnd), .vdd(vdd), .A(_11540_), .B(_11539_), .Y(_11541_) );
XNOR2X1 XNOR2X1_474 ( .gnd(gnd), .vdd(vdd), .A(_11541_), .B(_11527_), .Y(_11542_) );
INVX8 INVX8_283 ( .gnd(gnd), .vdd(vdd), .A(_11283__bF_buf2), .Y(_11543_) );
AOI21X1 AOI21X1_1954 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_188_), .B(_11543__bF_buf3), .C(_11466_), .Y(_11544_) );
NOR2X1 NOR2X1_1906 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_189_), .B(_11537__bF_buf2), .Y(_11545_) );
INVX1 INVX1_787 ( .gnd(gnd), .vdd(vdd), .A(_11545_), .Y(_11546_) );
NAND2X1 NAND2X1_1512 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_189_), .B(_11537__bF_buf1), .Y(_11547_) );
NAND2X1 NAND2X1_1513 ( .gnd(gnd), .vdd(vdd), .A(_11547_), .B(_11546_), .Y(_11548_) );
XOR2X1 XOR2X1_193 ( .gnd(gnd), .vdd(vdd), .A(_11548_), .B(_11544_), .Y(_11549_) );
AOI21X1 AOI21X1_1955 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_28_), .B(_11543__bF_buf2), .C(_11319_), .Y(_11550_) );
NOR2X1 NOR2X1_1907 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_29_), .B(_11537__bF_buf0), .Y(_11551_) );
INVX1 INVX1_788 ( .gnd(gnd), .vdd(vdd), .A(_11551_), .Y(_11552_) );
NAND2X1 NAND2X1_1514 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_29_), .B(_11537__bF_buf4), .Y(_11553_) );
NAND2X1 NAND2X1_1515 ( .gnd(gnd), .vdd(vdd), .A(_11553_), .B(_11552_), .Y(_11554_) );
XOR2X1 XOR2X1_194 ( .gnd(gnd), .vdd(vdd), .A(_11554_), .B(_11550_), .Y(_11555_) );
INVX1 INVX1_789 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_4_), .Y(_11556_) );
OAI21X1 OAI21X1_3226 ( .gnd(gnd), .vdd(vdd), .A(_11556_), .B(_11283__bF_buf1), .C(_11307_), .Y(_11557_) );
INVX1 INVX1_790 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_5_), .Y(_11558_) );
OAI21X1 OAI21X1_3227 ( .gnd(gnd), .vdd(vdd), .A(_11536__bF_buf2), .B(_11534__bF_buf2), .C(_11558_), .Y(_11559_) );
INVX8 INVX8_284 ( .gnd(gnd), .vdd(vdd), .A(_11537__bF_buf3), .Y(_11560_) );
NOR2X1 NOR2X1_1908 ( .gnd(gnd), .vdd(vdd), .A(_11558_), .B(_11560__bF_buf3), .Y(_11561_) );
INVX1 INVX1_791 ( .gnd(gnd), .vdd(vdd), .A(_11561_), .Y(_11562_) );
NAND2X1 NAND2X1_1516 ( .gnd(gnd), .vdd(vdd), .A(_11559_), .B(_11562_), .Y(_11563_) );
AOI21X1 AOI21X1_1956 ( .gnd(gnd), .vdd(vdd), .A(_11557_), .B(_11563_), .C(_9341_), .Y(_11564_) );
OAI21X1 OAI21X1_3228 ( .gnd(gnd), .vdd(vdd), .A(_11557_), .B(_11563_), .C(_11564_), .Y(_11565_) );
AOI21X1 AOI21X1_1957 ( .gnd(gnd), .vdd(vdd), .A(_9932_), .B(_9345_), .C(micro_hash_ucr_3_pipe10_bF_buf2), .Y(_11566_) );
OAI21X1 OAI21X1_3229 ( .gnd(gnd), .vdd(vdd), .A(H_3_21_), .B(_9345_), .C(_11566_), .Y(_11567_) );
OAI21X1 OAI21X1_3230 ( .gnd(gnd), .vdd(vdd), .A(_9341_), .B(micro_hash_ucr_3_pipe10_bF_buf1), .C(_11567_), .Y(_11568_) );
NOR2X1 NOR2X1_1909 ( .gnd(gnd), .vdd(vdd), .A(_11300_), .B(_11298_), .Y(_11569_) );
AOI21X1 AOI21X1_1958 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_12_), .B(_11543__bF_buf1), .C(_11569_), .Y(_11570_) );
NOR2X1 NOR2X1_1910 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_13_), .B(_11537__bF_buf2), .Y(_11571_) );
INVX1 INVX1_792 ( .gnd(gnd), .vdd(vdd), .A(_11571_), .Y(_11572_) );
NAND2X1 NAND2X1_1517 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_13_), .B(_11537__bF_buf1), .Y(_11573_) );
NAND2X1 NAND2X1_1518 ( .gnd(gnd), .vdd(vdd), .A(_11573_), .B(_11572_), .Y(_11574_) );
XNOR2X1 XNOR2X1_475 ( .gnd(gnd), .vdd(vdd), .A(_11574_), .B(_11570_), .Y(_11575_) );
OAI21X1 OAI21X1_3231 ( .gnd(gnd), .vdd(vdd), .A(_11575_), .B(_9342_), .C(_9340_), .Y(_11576_) );
AOI21X1 AOI21X1_1959 ( .gnd(gnd), .vdd(vdd), .A(_11568_), .B(_11565_), .C(_11576_), .Y(_11577_) );
AOI21X1 AOI21X1_1960 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_20_), .B(_11543__bF_buf0), .C(_11296_), .Y(_11578_) );
INVX1 INVX1_793 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_21_), .Y(_11579_) );
OAI21X1 OAI21X1_3232 ( .gnd(gnd), .vdd(vdd), .A(_11536__bF_buf1), .B(_11534__bF_buf1), .C(_11579_), .Y(_11580_) );
INVX1 INVX1_794 ( .gnd(gnd), .vdd(vdd), .A(_11580_), .Y(_11581_) );
NOR2X1 NOR2X1_1911 ( .gnd(gnd), .vdd(vdd), .A(_11579_), .B(_11560__bF_buf2), .Y(_11582_) );
NOR2X1 NOR2X1_1912 ( .gnd(gnd), .vdd(vdd), .A(_11581_), .B(_11582_), .Y(_11583_) );
OAI21X1 OAI21X1_3233 ( .gnd(gnd), .vdd(vdd), .A(_11583_), .B(_11578_), .C(micro_hash_ucr_3_pipe12), .Y(_11584_) );
AOI21X1 AOI21X1_1961 ( .gnd(gnd), .vdd(vdd), .A(_11578_), .B(_11583_), .C(_11584_), .Y(_11585_) );
OAI21X1 OAI21X1_3234 ( .gnd(gnd), .vdd(vdd), .A(_11577_), .B(_11585_), .C(_9335__bF_buf1), .Y(_11586_) );
OAI21X1 OAI21X1_3235 ( .gnd(gnd), .vdd(vdd), .A(_9335__bF_buf0), .B(_11555_), .C(_11586_), .Y(_11587_) );
NAND2X1 NAND2X1_1519 ( .gnd(gnd), .vdd(vdd), .A(_9336__bF_buf2), .B(_11587_), .Y(_11588_) );
AOI21X1 AOI21X1_1962 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_36_), .B(_11543__bF_buf3), .C(_11288_), .Y(_11589_) );
INVX2 INVX2_384 ( .gnd(gnd), .vdd(vdd), .A(_11589_), .Y(_11590_) );
INVX1 INVX1_795 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_37_), .Y(_11591_) );
OAI21X1 OAI21X1_3236 ( .gnd(gnd), .vdd(vdd), .A(_11536__bF_buf0), .B(_11534__bF_buf0), .C(_11591_), .Y(_11592_) );
NOR2X1 NOR2X1_1913 ( .gnd(gnd), .vdd(vdd), .A(_11591_), .B(_11560__bF_buf1), .Y(_11593_) );
INVX1 INVX1_796 ( .gnd(gnd), .vdd(vdd), .A(_11593_), .Y(_11594_) );
NAND2X1 NAND2X1_1520 ( .gnd(gnd), .vdd(vdd), .A(_11592_), .B(_11594_), .Y(_11595_) );
AOI21X1 AOI21X1_1963 ( .gnd(gnd), .vdd(vdd), .A(_11590_), .B(_11595_), .C(_9336__bF_buf1), .Y(_11596_) );
OAI21X1 OAI21X1_3237 ( .gnd(gnd), .vdd(vdd), .A(_11590_), .B(_11595_), .C(_11596_), .Y(_11597_) );
AND2X2 AND2X2_733 ( .gnd(gnd), .vdd(vdd), .A(_11597_), .B(_9334__bF_buf3), .Y(_11598_) );
AOI21X1 AOI21X1_1964 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_44_), .B(_11543__bF_buf2), .C(_11328_), .Y(_11599_) );
NOR2X1 NOR2X1_1914 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_45_), .B(_11537__bF_buf0), .Y(_11600_) );
INVX1 INVX1_797 ( .gnd(gnd), .vdd(vdd), .A(_11600_), .Y(_11601_) );
NAND2X1 NAND2X1_1521 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_45_), .B(_11537__bF_buf4), .Y(_11602_) );
NAND2X1 NAND2X1_1522 ( .gnd(gnd), .vdd(vdd), .A(_11602_), .B(_11601_), .Y(_11603_) );
AND2X2 AND2X2_734 ( .gnd(gnd), .vdd(vdd), .A(_11603_), .B(_11599_), .Y(_11604_) );
OAI21X1 OAI21X1_3238 ( .gnd(gnd), .vdd(vdd), .A(_11603_), .B(_11599_), .C(micro_hash_ucr_3_pipe18_bF_buf2), .Y(_11605_) );
OAI21X1 OAI21X1_3239 ( .gnd(gnd), .vdd(vdd), .A(_11604_), .B(_11605_), .C(_9329__bF_buf2), .Y(_11606_) );
AOI21X1 AOI21X1_1965 ( .gnd(gnd), .vdd(vdd), .A(_11598_), .B(_11588_), .C(_11606_), .Y(_11607_) );
AOI21X1 AOI21X1_1966 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_52_), .B(_11543__bF_buf1), .C(_11337_), .Y(_11608_) );
NOR2X1 NOR2X1_1915 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_53_), .B(_11537__bF_buf3), .Y(_11609_) );
INVX1 INVX1_798 ( .gnd(gnd), .vdd(vdd), .A(_11609_), .Y(_11610_) );
NAND2X1 NAND2X1_1523 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_53_), .B(_11537__bF_buf2), .Y(_11611_) );
NAND2X1 NAND2X1_1524 ( .gnd(gnd), .vdd(vdd), .A(_11611_), .B(_11610_), .Y(_11612_) );
XOR2X1 XOR2X1_195 ( .gnd(gnd), .vdd(vdd), .A(_11612_), .B(_11608_), .Y(_11613_) );
OAI21X1 OAI21X1_3240 ( .gnd(gnd), .vdd(vdd), .A(_11613_), .B(_9329__bF_buf1), .C(_9330__bF_buf2), .Y(_11614_) );
OAI21X1 OAI21X1_3241 ( .gnd(gnd), .vdd(vdd), .A(_9272_), .B(_11283__bF_buf0), .C(_11345_), .Y(_11615_) );
XNOR2X1 XNOR2X1_476 ( .gnd(gnd), .vdd(vdd), .A(_11537__bF_buf1), .B(micro_hash_ucr_3_Wx_61_), .Y(_11616_) );
XNOR2X1 XNOR2X1_477 ( .gnd(gnd), .vdd(vdd), .A(_11616_), .B(_11615_), .Y(_11617_) );
AOI21X1 AOI21X1_1967 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe22_bF_buf2), .B(_11617_), .C(micro_hash_ucr_3_pipe24_bF_buf2), .Y(_11618_) );
OAI21X1 OAI21X1_3242 ( .gnd(gnd), .vdd(vdd), .A(_11607_), .B(_11614_), .C(_11618_), .Y(_11619_) );
AOI21X1 AOI21X1_1968 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_68_), .B(_11543__bF_buf0), .C(_11353_), .Y(_11620_) );
XNOR2X1 XNOR2X1_478 ( .gnd(gnd), .vdd(vdd), .A(_11537__bF_buf0), .B(micro_hash_ucr_3_Wx_69_), .Y(_11621_) );
XNOR2X1 XNOR2X1_479 ( .gnd(gnd), .vdd(vdd), .A(_11620_), .B(_11621_), .Y(_11622_) );
AOI21X1 AOI21X1_1969 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe24_bF_buf1), .B(_11622_), .C(micro_hash_ucr_3_pipe26_bF_buf1), .Y(_11623_) );
OAI21X1 OAI21X1_3243 ( .gnd(gnd), .vdd(vdd), .A(_9171_), .B(_11283__bF_buf5), .C(_11361_), .Y(_11624_) );
OAI21X1 OAI21X1_3244 ( .gnd(gnd), .vdd(vdd), .A(_11536__bF_buf3), .B(_11534__bF_buf3), .C(_9174_), .Y(_11625_) );
NAND2X1 NAND2X1_1525 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_77_), .B(_11537__bF_buf4), .Y(_11626_) );
AOI21X1 AOI21X1_1970 ( .gnd(gnd), .vdd(vdd), .A(_11625_), .B(_11626_), .C(_11624_), .Y(_11627_) );
INVX1 INVX1_799 ( .gnd(gnd), .vdd(vdd), .A(_11624_), .Y(_11628_) );
NAND2X1 NAND2X1_1526 ( .gnd(gnd), .vdd(vdd), .A(_11625_), .B(_11626_), .Y(_11629_) );
OAI21X1 OAI21X1_3245 ( .gnd(gnd), .vdd(vdd), .A(_11628_), .B(_11629_), .C(micro_hash_ucr_3_pipe26_bF_buf0), .Y(_11630_) );
OAI21X1 OAI21X1_3246 ( .gnd(gnd), .vdd(vdd), .A(_11630_), .B(_11627_), .C(_9324__bF_buf0), .Y(_11631_) );
AOI21X1 AOI21X1_1971 ( .gnd(gnd), .vdd(vdd), .A(_11623_), .B(_11619_), .C(_11631_), .Y(_11632_) );
OAI21X1 OAI21X1_3247 ( .gnd(gnd), .vdd(vdd), .A(_9226_), .B(_11283__bF_buf4), .C(_11369_), .Y(_11633_) );
OAI21X1 OAI21X1_3248 ( .gnd(gnd), .vdd(vdd), .A(_11536__bF_buf2), .B(_11534__bF_buf2), .C(_9229_), .Y(_11634_) );
NOR2X1 NOR2X1_1916 ( .gnd(gnd), .vdd(vdd), .A(_9229_), .B(_11560__bF_buf0), .Y(_11635_) );
INVX1 INVX1_800 ( .gnd(gnd), .vdd(vdd), .A(_11635_), .Y(_11636_) );
NAND2X1 NAND2X1_1527 ( .gnd(gnd), .vdd(vdd), .A(_11634_), .B(_11636_), .Y(_11637_) );
XNOR2X1 XNOR2X1_480 ( .gnd(gnd), .vdd(vdd), .A(_11637_), .B(_11633_), .Y(_11638_) );
OAI21X1 OAI21X1_3249 ( .gnd(gnd), .vdd(vdd), .A(_11638_), .B(_9324__bF_buf4), .C(_9322__bF_buf2), .Y(_11639_) );
OAI21X1 OAI21X1_3250 ( .gnd(gnd), .vdd(vdd), .A(_9198_), .B(_11283__bF_buf3), .C(_11376_), .Y(_11640_) );
XNOR2X1 XNOR2X1_481 ( .gnd(gnd), .vdd(vdd), .A(_11537__bF_buf3), .B(micro_hash_ucr_3_Wx_93_), .Y(_11641_) );
XNOR2X1 XNOR2X1_482 ( .gnd(gnd), .vdd(vdd), .A(_11640_), .B(_11641_), .Y(_11642_) );
AOI21X1 AOI21X1_1972 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe30_bF_buf0), .B(_11642_), .C(micro_hash_ucr_3_pipe32_bF_buf3), .Y(_11643_) );
OAI21X1 OAI21X1_3251 ( .gnd(gnd), .vdd(vdd), .A(_11632_), .B(_11639_), .C(_11643_), .Y(_11644_) );
INVX1 INVX1_801 ( .gnd(gnd), .vdd(vdd), .A(_11383_), .Y(_11645_) );
OAI21X1 OAI21X1_3252 ( .gnd(gnd), .vdd(vdd), .A(_9055_), .B(_11283__bF_buf2), .C(_11645_), .Y(_11646_) );
XNOR2X1 XNOR2X1_483 ( .gnd(gnd), .vdd(vdd), .A(_11537__bF_buf2), .B(micro_hash_ucr_3_Wx_101_), .Y(_11647_) );
AOI21X1 AOI21X1_1973 ( .gnd(gnd), .vdd(vdd), .A(_11647_), .B(_11646_), .C(_9317__bF_buf4), .Y(_11648_) );
OAI21X1 OAI21X1_3253 ( .gnd(gnd), .vdd(vdd), .A(_11646_), .B(_11647_), .C(_11648_), .Y(_11649_) );
AND2X2 AND2X2_735 ( .gnd(gnd), .vdd(vdd), .A(_11649_), .B(_9318__bF_buf0), .Y(_11650_) );
AOI21X1 AOI21X1_1974 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_108_), .B(_11543__bF_buf3), .C(_11391_), .Y(_11651_) );
OAI21X1 OAI21X1_3254 ( .gnd(gnd), .vdd(vdd), .A(_11536__bF_buf1), .B(_11534__bF_buf1), .C(_9151_), .Y(_11652_) );
NAND2X1 NAND2X1_1528 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_109_), .B(_11537__bF_buf1), .Y(_11653_) );
NAND2X1 NAND2X1_1529 ( .gnd(gnd), .vdd(vdd), .A(_11652_), .B(_11653_), .Y(_11654_) );
AND2X2 AND2X2_736 ( .gnd(gnd), .vdd(vdd), .A(_11651_), .B(_11654_), .Y(_11655_) );
OAI21X1 OAI21X1_3255 ( .gnd(gnd), .vdd(vdd), .A(_11651_), .B(_11654_), .C(micro_hash_ucr_3_pipe34_bF_buf0), .Y(_11656_) );
OAI21X1 OAI21X1_3256 ( .gnd(gnd), .vdd(vdd), .A(_11655_), .B(_11656_), .C(_9316__bF_buf2), .Y(_11657_) );
AOI21X1 AOI21X1_1975 ( .gnd(gnd), .vdd(vdd), .A(_11650_), .B(_11644_), .C(_11657_), .Y(_11658_) );
OAI21X1 OAI21X1_3257 ( .gnd(gnd), .vdd(vdd), .A(_9126_), .B(_11283__bF_buf1), .C(_11398_), .Y(_11659_) );
XNOR2X1 XNOR2X1_484 ( .gnd(gnd), .vdd(vdd), .A(_11537__bF_buf0), .B(micro_hash_ucr_3_Wx_117_), .Y(_11660_) );
XNOR2X1 XNOR2X1_485 ( .gnd(gnd), .vdd(vdd), .A(_11659_), .B(_11660_), .Y(_11661_) );
OAI21X1 OAI21X1_3258 ( .gnd(gnd), .vdd(vdd), .A(_11661_), .B(_9316__bF_buf1), .C(_9311__bF_buf3), .Y(_11662_) );
AOI21X1 AOI21X1_1976 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_124_), .B(_11543__bF_buf2), .C(_11405_), .Y(_11663_) );
OAI21X1 OAI21X1_3259 ( .gnd(gnd), .vdd(vdd), .A(_11536__bF_buf0), .B(_11534__bF_buf0), .C(_9032_), .Y(_11664_) );
NAND2X1 NAND2X1_1530 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_125_), .B(_11537__bF_buf4), .Y(_11665_) );
NAND2X1 NAND2X1_1531 ( .gnd(gnd), .vdd(vdd), .A(_11664_), .B(_11665_), .Y(_11666_) );
XOR2X1 XOR2X1_196 ( .gnd(gnd), .vdd(vdd), .A(_11663_), .B(_11666_), .Y(_11667_) );
AOI21X1 AOI21X1_1977 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe38_bF_buf3), .B(_11667_), .C(micro_hash_ucr_3_pipe40_bF_buf0), .Y(_11668_) );
OAI21X1 OAI21X1_3260 ( .gnd(gnd), .vdd(vdd), .A(_11658_), .B(_11662_), .C(_11668_), .Y(_11669_) );
OAI21X1 OAI21X1_3261 ( .gnd(gnd), .vdd(vdd), .A(_9084_), .B(_11283__bF_buf0), .C(_11413_), .Y(_11670_) );
XNOR2X1 XNOR2X1_486 ( .gnd(gnd), .vdd(vdd), .A(_11537__bF_buf3), .B(micro_hash_ucr_3_Wx_133_), .Y(_11671_) );
AOI21X1 AOI21X1_1978 ( .gnd(gnd), .vdd(vdd), .A(_11671_), .B(_11670_), .C(_9312__bF_buf2), .Y(_11672_) );
OAI21X1 OAI21X1_3262 ( .gnd(gnd), .vdd(vdd), .A(_11670_), .B(_11671_), .C(_11672_), .Y(_11673_) );
AND2X2 AND2X2_737 ( .gnd(gnd), .vdd(vdd), .A(_11673_), .B(_9310__bF_buf3), .Y(_11674_) );
AOI21X1 AOI21X1_1979 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_140_), .B(_11543__bF_buf1), .C(_11420_), .Y(_11675_) );
OAI21X1 OAI21X1_3263 ( .gnd(gnd), .vdd(vdd), .A(_11536__bF_buf3), .B(_11534__bF_buf3), .C(_9203_), .Y(_11676_) );
NAND2X1 NAND2X1_1532 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_141_), .B(_11537__bF_buf2), .Y(_11677_) );
NAND2X1 NAND2X1_1533 ( .gnd(gnd), .vdd(vdd), .A(_11676_), .B(_11677_), .Y(_11678_) );
AND2X2 AND2X2_738 ( .gnd(gnd), .vdd(vdd), .A(_11675_), .B(_11678_), .Y(_11679_) );
OAI21X1 OAI21X1_3264 ( .gnd(gnd), .vdd(vdd), .A(_11675_), .B(_11678_), .C(micro_hash_ucr_3_pipe42_bF_buf3), .Y(_11680_) );
OAI21X1 OAI21X1_3265 ( .gnd(gnd), .vdd(vdd), .A(_11679_), .B(_11680_), .C(_9305__bF_buf4), .Y(_11681_) );
AOI21X1 AOI21X1_1980 ( .gnd(gnd), .vdd(vdd), .A(_11674_), .B(_11669_), .C(_11681_), .Y(_11682_) );
OAI21X1 OAI21X1_3266 ( .gnd(gnd), .vdd(vdd), .A(_8948_), .B(_11283__bF_buf5), .C(_11427_), .Y(_11683_) );
OAI21X1 OAI21X1_3267 ( .gnd(gnd), .vdd(vdd), .A(_11536__bF_buf2), .B(_11534__bF_buf2), .C(_8951_), .Y(_11684_) );
NOR2X1 NOR2X1_1917 ( .gnd(gnd), .vdd(vdd), .A(_8951_), .B(_11560__bF_buf3), .Y(_11685_) );
INVX1 INVX1_802 ( .gnd(gnd), .vdd(vdd), .A(_11685_), .Y(_11686_) );
NAND2X1 NAND2X1_1534 ( .gnd(gnd), .vdd(vdd), .A(_11684_), .B(_11686_), .Y(_11687_) );
XNOR2X1 XNOR2X1_487 ( .gnd(gnd), .vdd(vdd), .A(_11687_), .B(_11683_), .Y(_11688_) );
OAI21X1 OAI21X1_3268 ( .gnd(gnd), .vdd(vdd), .A(_11688_), .B(_9305__bF_buf3), .C(_9306__bF_buf1), .Y(_11689_) );
OAI21X1 OAI21X1_3269 ( .gnd(gnd), .vdd(vdd), .A(_9005_), .B(_11283__bF_buf4), .C(_11437_), .Y(_11690_) );
OAI21X1 OAI21X1_3270 ( .gnd(gnd), .vdd(vdd), .A(_11536__bF_buf1), .B(_11534__bF_buf1), .C(_9008_), .Y(_11691_) );
INVX1 INVX1_803 ( .gnd(gnd), .vdd(vdd), .A(_11691_), .Y(_11692_) );
NOR2X1 NOR2X1_1918 ( .gnd(gnd), .vdd(vdd), .A(_9008_), .B(_11560__bF_buf2), .Y(_11693_) );
NOR2X1 NOR2X1_1919 ( .gnd(gnd), .vdd(vdd), .A(_11692_), .B(_11693_), .Y(_11694_) );
XOR2X1 XOR2X1_197 ( .gnd(gnd), .vdd(vdd), .A(_11690_), .B(_11694_), .Y(_11695_) );
AOI21X1 AOI21X1_1981 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe46_bF_buf0), .B(_11695_), .C(micro_hash_ucr_3_pipe48_bF_buf1), .Y(_11696_) );
OAI21X1 OAI21X1_3271 ( .gnd(gnd), .vdd(vdd), .A(_11682_), .B(_11689_), .C(_11696_), .Y(_11697_) );
AOI21X1 AOI21X1_1982 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_164_), .B(_11543__bF_buf0), .C(_11444_), .Y(_11698_) );
INVX2 INVX2_385 ( .gnd(gnd), .vdd(vdd), .A(_11698_), .Y(_11699_) );
OAI21X1 OAI21X1_3272 ( .gnd(gnd), .vdd(vdd), .A(_11536__bF_buf0), .B(_11534__bF_buf0), .C(_8981_), .Y(_11700_) );
NOR2X1 NOR2X1_1920 ( .gnd(gnd), .vdd(vdd), .A(_8981_), .B(_11560__bF_buf1), .Y(_11701_) );
INVX1 INVX1_804 ( .gnd(gnd), .vdd(vdd), .A(_11701_), .Y(_11702_) );
NAND2X1 NAND2X1_1535 ( .gnd(gnd), .vdd(vdd), .A(_11700_), .B(_11702_), .Y(_11703_) );
AOI21X1 AOI21X1_1983 ( .gnd(gnd), .vdd(vdd), .A(_11699_), .B(_11703_), .C(_9304__bF_buf0), .Y(_11704_) );
OAI21X1 OAI21X1_3273 ( .gnd(gnd), .vdd(vdd), .A(_11699_), .B(_11703_), .C(_11704_), .Y(_11705_) );
AND2X2 AND2X2_739 ( .gnd(gnd), .vdd(vdd), .A(_11705_), .B(_9299__bF_buf2), .Y(_11706_) );
OAI21X1 OAI21X1_3274 ( .gnd(gnd), .vdd(vdd), .A(_8848_), .B(_11283__bF_buf3), .C(_11451_), .Y(_11707_) );
OAI21X1 OAI21X1_3275 ( .gnd(gnd), .vdd(vdd), .A(_11536__bF_buf3), .B(_11534__bF_buf3), .C(_8851_), .Y(_11708_) );
NOR2X1 NOR2X1_1921 ( .gnd(gnd), .vdd(vdd), .A(_8851_), .B(_11560__bF_buf0), .Y(_11709_) );
INVX1 INVX1_805 ( .gnd(gnd), .vdd(vdd), .A(_11709_), .Y(_11710_) );
NAND2X1 NAND2X1_1536 ( .gnd(gnd), .vdd(vdd), .A(_11708_), .B(_11710_), .Y(_11711_) );
XOR2X1 XOR2X1_198 ( .gnd(gnd), .vdd(vdd), .A(_11711_), .B(_11707_), .Y(_11712_) );
OAI21X1 OAI21X1_3276 ( .gnd(gnd), .vdd(vdd), .A(_11712_), .B(_9299__bF_buf1), .C(_9300__bF_buf2), .Y(_11713_) );
AOI21X1 AOI21X1_1984 ( .gnd(gnd), .vdd(vdd), .A(_11706_), .B(_11697_), .C(_11713_), .Y(_11714_) );
AOI21X1 AOI21X1_1985 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_180_), .B(_11543__bF_buf3), .C(_11458_), .Y(_11715_) );
NOR2X1 NOR2X1_1922 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_181_), .B(_11537__bF_buf1), .Y(_11716_) );
NOR2X1 NOR2X1_1923 ( .gnd(gnd), .vdd(vdd), .A(_9089_), .B(_11560__bF_buf3), .Y(_11717_) );
NOR2X1 NOR2X1_1924 ( .gnd(gnd), .vdd(vdd), .A(_11716_), .B(_11717_), .Y(_11718_) );
OAI21X1 OAI21X1_3277 ( .gnd(gnd), .vdd(vdd), .A(_11718_), .B(_11715_), .C(micro_hash_ucr_3_pipe52_bF_buf4), .Y(_11719_) );
AOI21X1 AOI21X1_1986 ( .gnd(gnd), .vdd(vdd), .A(_11715_), .B(_11718_), .C(_11719_), .Y(_11720_) );
OAI21X1 OAI21X1_3278 ( .gnd(gnd), .vdd(vdd), .A(_11714_), .B(_11720_), .C(_9298__bF_buf2), .Y(_11721_) );
OAI21X1 OAI21X1_3279 ( .gnd(gnd), .vdd(vdd), .A(_9298__bF_buf1), .B(_11549_), .C(_11721_), .Y(_11722_) );
NAND2X1 NAND2X1_1537 ( .gnd(gnd), .vdd(vdd), .A(_9293__bF_buf2), .B(_11722_), .Y(_11723_) );
AOI21X1 AOI21X1_1987 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_196_), .B(_11543__bF_buf2), .C(_11472_), .Y(_11724_) );
INVX2 INVX2_386 ( .gnd(gnd), .vdd(vdd), .A(_11724_), .Y(_11725_) );
OAI21X1 OAI21X1_3280 ( .gnd(gnd), .vdd(vdd), .A(_11536__bF_buf2), .B(_11534__bF_buf2), .C(_8952_), .Y(_11726_) );
NOR2X1 NOR2X1_1925 ( .gnd(gnd), .vdd(vdd), .A(_8952_), .B(_11560__bF_buf2), .Y(_11727_) );
INVX1 INVX1_806 ( .gnd(gnd), .vdd(vdd), .A(_11727_), .Y(_11728_) );
NAND2X1 NAND2X1_1538 ( .gnd(gnd), .vdd(vdd), .A(_11726_), .B(_11728_), .Y(_11729_) );
AOI21X1 AOI21X1_1988 ( .gnd(gnd), .vdd(vdd), .A(_11725_), .B(_11729_), .C(_9293__bF_buf1), .Y(_11730_) );
OAI21X1 OAI21X1_3281 ( .gnd(gnd), .vdd(vdd), .A(_11725_), .B(_11729_), .C(_11730_), .Y(_11731_) );
AND2X2 AND2X2_740 ( .gnd(gnd), .vdd(vdd), .A(_11731_), .B(_9294__bF_buf0), .Y(_11732_) );
AOI21X1 AOI21X1_1989 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_204_), .B(_11543__bF_buf1), .C(_11480_), .Y(_11733_) );
NOR2X1 NOR2X1_1926 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_205_), .B(_11537__bF_buf0), .Y(_11734_) );
INVX1 INVX1_807 ( .gnd(gnd), .vdd(vdd), .A(_11734_), .Y(_11735_) );
NAND2X1 NAND2X1_1539 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_205_), .B(_11537__bF_buf4), .Y(_11736_) );
NAND2X1 NAND2X1_1540 ( .gnd(gnd), .vdd(vdd), .A(_11736_), .B(_11735_), .Y(_11737_) );
AND2X2 AND2X2_741 ( .gnd(gnd), .vdd(vdd), .A(_11737_), .B(_11733_), .Y(_11738_) );
OAI21X1 OAI21X1_3282 ( .gnd(gnd), .vdd(vdd), .A(_11737_), .B(_11733_), .C(micro_hash_ucr_3_pipe58_bF_buf1), .Y(_11739_) );
OAI21X1 OAI21X1_3283 ( .gnd(gnd), .vdd(vdd), .A(_11738_), .B(_11739_), .C(_9292__bF_buf0), .Y(_11740_) );
AOI21X1 AOI21X1_1990 ( .gnd(gnd), .vdd(vdd), .A(_11732_), .B(_11723_), .C(_11740_), .Y(_11741_) );
AOI21X1 AOI21X1_1991 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_212_), .B(_11543__bF_buf0), .C(_11488_), .Y(_11742_) );
OAI21X1 OAI21X1_3284 ( .gnd(gnd), .vdd(vdd), .A(_11536__bF_buf1), .B(_11534__bF_buf1), .C(_8982_), .Y(_11743_) );
INVX1 INVX1_808 ( .gnd(gnd), .vdd(vdd), .A(_11743_), .Y(_11744_) );
NOR2X1 NOR2X1_1927 ( .gnd(gnd), .vdd(vdd), .A(_8982_), .B(_11560__bF_buf1), .Y(_11745_) );
NOR2X1 NOR2X1_1928 ( .gnd(gnd), .vdd(vdd), .A(_11744_), .B(_11745_), .Y(_11746_) );
XNOR2X1 XNOR2X1_488 ( .gnd(gnd), .vdd(vdd), .A(_11746_), .B(_11742_), .Y(_11747_) );
OAI21X1 OAI21X1_3285 ( .gnd(gnd), .vdd(vdd), .A(_11747_), .B(_9292__bF_buf3), .C(_9287__bF_buf3), .Y(_11748_) );
AOI21X1 AOI21X1_1992 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_220_), .B(_11543__bF_buf3), .C(_11494_), .Y(_11749_) );
NOR2X1 NOR2X1_1929 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_221_), .B(_11537__bF_buf3), .Y(_11750_) );
INVX1 INVX1_809 ( .gnd(gnd), .vdd(vdd), .A(_11750_), .Y(_11751_) );
NAND2X1 NAND2X1_1541 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_221_), .B(_11537__bF_buf2), .Y(_11752_) );
NAND2X1 NAND2X1_1542 ( .gnd(gnd), .vdd(vdd), .A(_11752_), .B(_11751_), .Y(_11753_) );
XOR2X1 XOR2X1_199 ( .gnd(gnd), .vdd(vdd), .A(_11753_), .B(_11749_), .Y(_11754_) );
AOI21X1 AOI21X1_1993 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe62_bF_buf3), .B(_11754_), .C(micro_hash_ucr_3_pipe64_bF_buf3), .Y(_11755_) );
OAI21X1 OAI21X1_3286 ( .gnd(gnd), .vdd(vdd), .A(_11741_), .B(_11748_), .C(_11755_), .Y(_11756_) );
NOR2X1 NOR2X1_1930 ( .gnd(gnd), .vdd(vdd), .A(_11500_), .B(_11499_), .Y(_11757_) );
AOI21X1 AOI21X1_1994 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_228_), .B(_11543__bF_buf2), .C(_11757_), .Y(_11758_) );
INVX2 INVX2_387 ( .gnd(gnd), .vdd(vdd), .A(_11758_), .Y(_11759_) );
INVX1 INVX1_810 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_229_), .Y(_11760_) );
OAI21X1 OAI21X1_3287 ( .gnd(gnd), .vdd(vdd), .A(_11536__bF_buf0), .B(_11534__bF_buf0), .C(_11760_), .Y(_11761_) );
NOR2X1 NOR2X1_1931 ( .gnd(gnd), .vdd(vdd), .A(_11760_), .B(_11560__bF_buf0), .Y(_11762_) );
INVX1 INVX1_811 ( .gnd(gnd), .vdd(vdd), .A(_11762_), .Y(_11763_) );
NAND2X1 NAND2X1_1543 ( .gnd(gnd), .vdd(vdd), .A(_11761_), .B(_11763_), .Y(_11764_) );
AOI21X1 AOI21X1_1995 ( .gnd(gnd), .vdd(vdd), .A(_11759_), .B(_11764_), .C(_9288__bF_buf3), .Y(_11765_) );
OAI21X1 OAI21X1_3288 ( .gnd(gnd), .vdd(vdd), .A(_11759_), .B(_11764_), .C(_11765_), .Y(_11766_) );
AOI21X1 AOI21X1_1996 ( .gnd(gnd), .vdd(vdd), .A(_11766_), .B(_11756_), .C(micro_hash_ucr_3_pipe66_bF_buf0), .Y(_11767_) );
AOI21X1 AOI21X1_1997 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe66_bF_buf4), .B(_11542_), .C(_11767_), .Y(_11768_) );
AOI21X1 AOI21X1_1998 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_244_), .B(_11543__bF_buf1), .C(_11516_), .Y(_11769_) );
INVX1 INVX1_812 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_245_), .Y(_11770_) );
OAI21X1 OAI21X1_3289 ( .gnd(gnd), .vdd(vdd), .A(_11536__bF_buf3), .B(_11534__bF_buf3), .C(_11770_), .Y(_11771_) );
INVX1 INVX1_813 ( .gnd(gnd), .vdd(vdd), .A(_11771_), .Y(_11772_) );
NOR2X1 NOR2X1_1932 ( .gnd(gnd), .vdd(vdd), .A(_11770_), .B(_11560__bF_buf3), .Y(_11773_) );
NOR2X1 NOR2X1_1933 ( .gnd(gnd), .vdd(vdd), .A(_11772_), .B(_11773_), .Y(_11774_) );
AND2X2 AND2X2_742 ( .gnd(gnd), .vdd(vdd), .A(_11774_), .B(_11769_), .Y(_11775_) );
OAI21X1 OAI21X1_3290 ( .gnd(gnd), .vdd(vdd), .A(_11774_), .B(_11769_), .C(micro_hash_ucr_3_pipe68_bF_buf3), .Y(_11776_) );
OAI22X1 OAI22X1_143 ( .gnd(gnd), .vdd(vdd), .A(_11775_), .B(_11776_), .C(_11768_), .D(micro_hash_ucr_3_pipe68_bF_buf2), .Y(_11777_) );
NAND2X1 NAND2X1_1544 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_252_), .B(_11543__bF_buf0), .Y(_11778_) );
OAI21X1 OAI21X1_3291 ( .gnd(gnd), .vdd(vdd), .A(_11521_), .B(_11520_), .C(_11778_), .Y(_11779_) );
INVX1 INVX1_814 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_253_), .Y(_11780_) );
OAI21X1 OAI21X1_3292 ( .gnd(gnd), .vdd(vdd), .A(_11536__bF_buf2), .B(_11534__bF_buf2), .C(_11780_), .Y(_11781_) );
NOR2X1 NOR2X1_1934 ( .gnd(gnd), .vdd(vdd), .A(_11780_), .B(_11560__bF_buf2), .Y(_11782_) );
INVX1 INVX1_815 ( .gnd(gnd), .vdd(vdd), .A(_11782_), .Y(_11783_) );
NAND2X1 NAND2X1_1545 ( .gnd(gnd), .vdd(vdd), .A(_11781_), .B(_11783_), .Y(_11784_) );
XOR2X1 XOR2X1_200 ( .gnd(gnd), .vdd(vdd), .A(_11784_), .B(_11779_), .Y(_11785_) );
OAI22X1 OAI22X1_144 ( .gnd(gnd), .vdd(vdd), .A(_11524_), .B(_11785_), .C(_11777_), .D(_10381_), .Y(_8702__5_) );
OAI21X1 OAI21X1_3293 ( .gnd(gnd), .vdd(vdd), .A(_10255_), .B(_11528_), .C(_11533_), .Y(_11786_) );
XOR2X1 XOR2X1_201 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_k_6_), .B(micro_hash_ucr_3_x_6_), .Y(_11787_) );
NOR2X1 NOR2X1_1935 ( .gnd(gnd), .vdd(vdd), .A(_11787_), .B(_11786_), .Y(_11788_) );
OAI21X1 OAI21X1_3294 ( .gnd(gnd), .vdd(vdd), .A(_11534__bF_buf1), .B(_11530_), .C(_11787_), .Y(_11789_) );
INVX4 INVX4_154 ( .gnd(gnd), .vdd(vdd), .A(_11789_), .Y(_11790_) );
NOR2X1 NOR2X1_1936 ( .gnd(gnd), .vdd(vdd), .A(_11788_), .B(_11790_), .Y(_11791_) );
XOR2X1 XOR2X1_202 ( .gnd(gnd), .vdd(vdd), .A(_11791__bF_buf5), .B(micro_hash_ucr_3_Wx_14_), .Y(_11792_) );
OAI21X1 OAI21X1_3295 ( .gnd(gnd), .vdd(vdd), .A(_11570_), .B(_11571_), .C(_11573_), .Y(_11793_) );
XNOR2X1 XNOR2X1_489 ( .gnd(gnd), .vdd(vdd), .A(_11793_), .B(_11792_), .Y(_11794_) );
NAND2X1 NAND2X1_1546 ( .gnd(gnd), .vdd(vdd), .A(H_3_22_), .B(micro_hash_ucr_3_pipe6_bF_buf3), .Y(_11795_) );
OAI21X1 OAI21X1_3296 ( .gnd(gnd), .vdd(vdd), .A(_12893_), .B(micro_hash_ucr_3_pipe6_bF_buf2), .C(_11795_), .Y(_11796_) );
XNOR2X1 XNOR2X1_490 ( .gnd(gnd), .vdd(vdd), .A(_11791__bF_buf4), .B(micro_hash_ucr_3_Wx_6_), .Y(_11797_) );
AOI21X1 AOI21X1_1999 ( .gnd(gnd), .vdd(vdd), .A(_11559_), .B(_11557_), .C(_11561_), .Y(_11798_) );
AND2X2 AND2X2_743 ( .gnd(gnd), .vdd(vdd), .A(_11798_), .B(_11797_), .Y(_11799_) );
NOR2X1 NOR2X1_1937 ( .gnd(gnd), .vdd(vdd), .A(_11797_), .B(_11798_), .Y(_11800_) );
OAI21X1 OAI21X1_3297 ( .gnd(gnd), .vdd(vdd), .A(_11799_), .B(_11800_), .C(micro_hash_ucr_3_pipe8), .Y(_11801_) );
OAI21X1 OAI21X1_3298 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe8), .B(_11796_), .C(_11801_), .Y(_11802_) );
MUX2X1 MUX2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_11802_), .B(_11794_), .S(_9342_), .Y(_11803_) );
INVX2 INVX2_388 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_22_), .Y(_11804_) );
XNOR2X1 XNOR2X1_491 ( .gnd(gnd), .vdd(vdd), .A(_11791__bF_buf3), .B(_11804_), .Y(_11805_) );
INVX1 INVX1_816 ( .gnd(gnd), .vdd(vdd), .A(_11582_), .Y(_11806_) );
OAI21X1 OAI21X1_3299 ( .gnd(gnd), .vdd(vdd), .A(_11578_), .B(_11581_), .C(_11806_), .Y(_11807_) );
NAND2X1 NAND2X1_1547 ( .gnd(gnd), .vdd(vdd), .A(_11805_), .B(_11807_), .Y(_11808_) );
INVX1 INVX1_817 ( .gnd(gnd), .vdd(vdd), .A(_11808_), .Y(_11809_) );
NOR2X1 NOR2X1_1938 ( .gnd(gnd), .vdd(vdd), .A(_11805_), .B(_11807_), .Y(_11810_) );
OAI21X1 OAI21X1_3300 ( .gnd(gnd), .vdd(vdd), .A(_11809_), .B(_11810_), .C(micro_hash_ucr_3_pipe12), .Y(_11811_) );
OAI21X1 OAI21X1_3301 ( .gnd(gnd), .vdd(vdd), .A(_11803_), .B(micro_hash_ucr_3_pipe12), .C(_11811_), .Y(_11812_) );
INVX2 INVX2_389 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_30_), .Y(_11813_) );
XNOR2X1 XNOR2X1_492 ( .gnd(gnd), .vdd(vdd), .A(_11791__bF_buf2), .B(_11813_), .Y(_11814_) );
OAI21X1 OAI21X1_3302 ( .gnd(gnd), .vdd(vdd), .A(_11550_), .B(_11551_), .C(_11553_), .Y(_11815_) );
XNOR2X1 XNOR2X1_493 ( .gnd(gnd), .vdd(vdd), .A(_11815_), .B(_11814_), .Y(_11816_) );
MUX2X1 MUX2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_11812_), .B(_11816_), .S(_9335__bF_buf3), .Y(_11817_) );
NAND2X1 NAND2X1_1548 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_38_), .B(_11791__bF_buf1), .Y(_11818_) );
INVX1 INVX1_818 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_38_), .Y(_11819_) );
OAI21X1 OAI21X1_3303 ( .gnd(gnd), .vdd(vdd), .A(_11790_), .B(_11788_), .C(_11819_), .Y(_11820_) );
AND2X2 AND2X2_744 ( .gnd(gnd), .vdd(vdd), .A(_11818_), .B(_11820_), .Y(_11821_) );
AOI21X1 AOI21X1_2000 ( .gnd(gnd), .vdd(vdd), .A(_11592_), .B(_11590_), .C(_11593_), .Y(_11822_) );
XNOR2X1 XNOR2X1_494 ( .gnd(gnd), .vdd(vdd), .A(_11822_), .B(_11821_), .Y(_11823_) );
MUX2X1 MUX2X1_33 ( .gnd(gnd), .vdd(vdd), .A(_11817_), .B(_11823_), .S(_9336__bF_buf0), .Y(_11824_) );
INVX2 INVX2_390 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_46_), .Y(_11825_) );
XNOR2X1 XNOR2X1_495 ( .gnd(gnd), .vdd(vdd), .A(_11791__bF_buf0), .B(_11825_), .Y(_11826_) );
OAI21X1 OAI21X1_3304 ( .gnd(gnd), .vdd(vdd), .A(_11599_), .B(_11600_), .C(_11602_), .Y(_11827_) );
OR2X2 OR2X2_77 ( .gnd(gnd), .vdd(vdd), .A(_11827_), .B(_11826_), .Y(_11828_) );
NAND2X1 NAND2X1_1549 ( .gnd(gnd), .vdd(vdd), .A(_11826_), .B(_11827_), .Y(_11829_) );
NAND3X1 NAND3X1_598 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe18_bF_buf1), .B(_11829_), .C(_11828_), .Y(_11830_) );
OAI21X1 OAI21X1_3305 ( .gnd(gnd), .vdd(vdd), .A(_11824_), .B(micro_hash_ucr_3_pipe18_bF_buf0), .C(_11830_), .Y(_11831_) );
INVX2 INVX2_391 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_54_), .Y(_11832_) );
XNOR2X1 XNOR2X1_496 ( .gnd(gnd), .vdd(vdd), .A(_11791__bF_buf5), .B(_11832_), .Y(_11833_) );
OAI21X1 OAI21X1_3306 ( .gnd(gnd), .vdd(vdd), .A(_11608_), .B(_11609_), .C(_11611_), .Y(_11834_) );
OAI21X1 OAI21X1_3307 ( .gnd(gnd), .vdd(vdd), .A(_11834_), .B(_11833_), .C(micro_hash_ucr_3_pipe20_bF_buf2), .Y(_11835_) );
AOI21X1 AOI21X1_2001 ( .gnd(gnd), .vdd(vdd), .A(_11833_), .B(_11834_), .C(_11835_), .Y(_11836_) );
AOI21X1 AOI21X1_2002 ( .gnd(gnd), .vdd(vdd), .A(_9329__bF_buf0), .B(_11831_), .C(_11836_), .Y(_11837_) );
XNOR2X1 XNOR2X1_497 ( .gnd(gnd), .vdd(vdd), .A(_11791__bF_buf4), .B(_9278_), .Y(_11838_) );
OAI21X1 OAI21X1_3308 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_61_), .B(_11537__bF_buf1), .C(_11615_), .Y(_11839_) );
OAI21X1 OAI21X1_3309 ( .gnd(gnd), .vdd(vdd), .A(_9275_), .B(_11560__bF_buf1), .C(_11839_), .Y(_11840_) );
OR2X2 OR2X2_78 ( .gnd(gnd), .vdd(vdd), .A(_11840_), .B(_11838_), .Y(_11841_) );
NAND2X1 NAND2X1_1550 ( .gnd(gnd), .vdd(vdd), .A(_11838_), .B(_11840_), .Y(_11842_) );
AND2X2 AND2X2_745 ( .gnd(gnd), .vdd(vdd), .A(_11841_), .B(_11842_), .Y(_11843_) );
OAI21X1 OAI21X1_3310 ( .gnd(gnd), .vdd(vdd), .A(_11843_), .B(_9330__bF_buf1), .C(_9328__bF_buf3), .Y(_11844_) );
AOI21X1 AOI21X1_2003 ( .gnd(gnd), .vdd(vdd), .A(_9330__bF_buf0), .B(_11837_), .C(_11844_), .Y(_11845_) );
XNOR2X1 XNOR2X1_498 ( .gnd(gnd), .vdd(vdd), .A(_11791__bF_buf3), .B(micro_hash_ucr_3_Wx_70_), .Y(_11846_) );
OAI21X1 OAI21X1_3311 ( .gnd(gnd), .vdd(vdd), .A(_9251_), .B(_11560__bF_buf0), .C(_11620_), .Y(_11847_) );
OAI21X1 OAI21X1_3312 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_69_), .B(_11537__bF_buf0), .C(_11847_), .Y(_11848_) );
AOI21X1 AOI21X1_2004 ( .gnd(gnd), .vdd(vdd), .A(_11846_), .B(_11848_), .C(_9328__bF_buf2), .Y(_11849_) );
OAI21X1 OAI21X1_3313 ( .gnd(gnd), .vdd(vdd), .A(_11846_), .B(_11848_), .C(_11849_), .Y(_11850_) );
NAND2X1 NAND2X1_1551 ( .gnd(gnd), .vdd(vdd), .A(_9323__bF_buf0), .B(_11850_), .Y(_11851_) );
INVX8 INVX8_285 ( .gnd(gnd), .vdd(vdd), .A(_11791__bF_buf2), .Y(_11852_) );
NOR2X1 NOR2X1_1939 ( .gnd(gnd), .vdd(vdd), .A(_9177_), .B(_11852__bF_buf3), .Y(_11853_) );
INVX1 INVX1_819 ( .gnd(gnd), .vdd(vdd), .A(_11853_), .Y(_11854_) );
OAI21X1 OAI21X1_3314 ( .gnd(gnd), .vdd(vdd), .A(_11790_), .B(_11788_), .C(_9177_), .Y(_11855_) );
NAND2X1 NAND2X1_1552 ( .gnd(gnd), .vdd(vdd), .A(_11855_), .B(_11854_), .Y(_11856_) );
INVX1 INVX1_820 ( .gnd(gnd), .vdd(vdd), .A(_11625_), .Y(_11857_) );
OAI21X1 OAI21X1_3315 ( .gnd(gnd), .vdd(vdd), .A(_11628_), .B(_11857_), .C(_11626_), .Y(_11858_) );
XOR2X1 XOR2X1_203 ( .gnd(gnd), .vdd(vdd), .A(_11858_), .B(_11856_), .Y(_11859_) );
AOI21X1 AOI21X1_2005 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe26_bF_buf4), .B(_11859_), .C(micro_hash_ucr_3_pipe28_bF_buf0), .Y(_11860_) );
OAI21X1 OAI21X1_3316 ( .gnd(gnd), .vdd(vdd), .A(_11845_), .B(_11851_), .C(_11860_), .Y(_11861_) );
XNOR2X1 XNOR2X1_499 ( .gnd(gnd), .vdd(vdd), .A(_11791__bF_buf1), .B(_9232_), .Y(_11862_) );
AOI21X1 AOI21X1_2006 ( .gnd(gnd), .vdd(vdd), .A(_11634_), .B(_11633_), .C(_11635_), .Y(_11863_) );
INVX1 INVX1_821 ( .gnd(gnd), .vdd(vdd), .A(_11863_), .Y(_11864_) );
NAND2X1 NAND2X1_1553 ( .gnd(gnd), .vdd(vdd), .A(_11862_), .B(_11864_), .Y(_11865_) );
INVX1 INVX1_822 ( .gnd(gnd), .vdd(vdd), .A(_11865_), .Y(_11866_) );
OAI21X1 OAI21X1_3317 ( .gnd(gnd), .vdd(vdd), .A(_11864_), .B(_11862_), .C(micro_hash_ucr_3_pipe28_bF_buf4), .Y(_11867_) );
OAI21X1 OAI21X1_3318 ( .gnd(gnd), .vdd(vdd), .A(_11866_), .B(_11867_), .C(_11861_), .Y(_11868_) );
NOR2X1 NOR2X1_1940 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe30_bF_buf4), .B(_11868_), .Y(_11869_) );
XNOR2X1 XNOR2X1_500 ( .gnd(gnd), .vdd(vdd), .A(_11791__bF_buf0), .B(_9206_), .Y(_11870_) );
OAI21X1 OAI21X1_3319 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_93_), .B(_11537__bF_buf4), .C(_11640_), .Y(_11871_) );
OAI21X1 OAI21X1_3320 ( .gnd(gnd), .vdd(vdd), .A(_9202_), .B(_11560__bF_buf3), .C(_11871_), .Y(_11872_) );
XOR2X1 XOR2X1_204 ( .gnd(gnd), .vdd(vdd), .A(_11872_), .B(_11870_), .Y(_11873_) );
OAI21X1 OAI21X1_3321 ( .gnd(gnd), .vdd(vdd), .A(_11873_), .B(_9322__bF_buf1), .C(_9317__bF_buf3), .Y(_11874_) );
XNOR2X1 XNOR2X1_501 ( .gnd(gnd), .vdd(vdd), .A(_11791__bF_buf5), .B(_9061_), .Y(_11875_) );
OAI21X1 OAI21X1_3322 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_101_), .B(_11537__bF_buf3), .C(_11646_), .Y(_11876_) );
OAI21X1 OAI21X1_3323 ( .gnd(gnd), .vdd(vdd), .A(_9058_), .B(_11560__bF_buf2), .C(_11876_), .Y(_11877_) );
XOR2X1 XOR2X1_205 ( .gnd(gnd), .vdd(vdd), .A(_11877_), .B(_11875_), .Y(_11878_) );
AOI21X1 AOI21X1_2007 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe32_bF_buf2), .B(_11878_), .C(micro_hash_ucr_3_pipe34_bF_buf4), .Y(_11879_) );
OAI21X1 OAI21X1_3324 ( .gnd(gnd), .vdd(vdd), .A(_11869_), .B(_11874_), .C(_11879_), .Y(_11880_) );
NOR2X1 NOR2X1_1941 ( .gnd(gnd), .vdd(vdd), .A(_9154_), .B(_11852__bF_buf2), .Y(_11881_) );
INVX1 INVX1_823 ( .gnd(gnd), .vdd(vdd), .A(_11881_), .Y(_11882_) );
OAI21X1 OAI21X1_3325 ( .gnd(gnd), .vdd(vdd), .A(_11790_), .B(_11788_), .C(_9154_), .Y(_11883_) );
NAND2X1 NAND2X1_1554 ( .gnd(gnd), .vdd(vdd), .A(_11883_), .B(_11882_), .Y(_11884_) );
INVX1 INVX1_824 ( .gnd(gnd), .vdd(vdd), .A(_11652_), .Y(_11885_) );
OAI21X1 OAI21X1_3326 ( .gnd(gnd), .vdd(vdd), .A(_11651_), .B(_11885_), .C(_11653_), .Y(_11886_) );
XOR2X1 XOR2X1_206 ( .gnd(gnd), .vdd(vdd), .A(_11884_), .B(_11886_), .Y(_11887_) );
AOI21X1 AOI21X1_2008 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe34_bF_buf3), .B(_11887_), .C(micro_hash_ucr_3_pipe36_bF_buf0), .Y(_11888_) );
XNOR2X1 XNOR2X1_502 ( .gnd(gnd), .vdd(vdd), .A(_11791__bF_buf4), .B(_9132_), .Y(_11889_) );
OAI21X1 OAI21X1_3327 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_117_), .B(_11537__bF_buf2), .C(_11659_), .Y(_11890_) );
OAI21X1 OAI21X1_3328 ( .gnd(gnd), .vdd(vdd), .A(_9129_), .B(_11560__bF_buf1), .C(_11890_), .Y(_11891_) );
OAI21X1 OAI21X1_3329 ( .gnd(gnd), .vdd(vdd), .A(_11891_), .B(_11889_), .C(micro_hash_ucr_3_pipe36_bF_buf4), .Y(_11892_) );
AOI21X1 AOI21X1_2009 ( .gnd(gnd), .vdd(vdd), .A(_11889_), .B(_11891_), .C(_11892_), .Y(_11893_) );
AOI21X1 AOI21X1_2010 ( .gnd(gnd), .vdd(vdd), .A(_11888_), .B(_11880_), .C(_11893_), .Y(_11894_) );
NAND2X1 NAND2X1_1555 ( .gnd(gnd), .vdd(vdd), .A(_9311__bF_buf2), .B(_11894_), .Y(_11895_) );
XNOR2X1 XNOR2X1_503 ( .gnd(gnd), .vdd(vdd), .A(_11791__bF_buf3), .B(_8985_), .Y(_11896_) );
INVX1 INVX1_825 ( .gnd(gnd), .vdd(vdd), .A(_11664_), .Y(_11897_) );
OAI21X1 OAI21X1_3330 ( .gnd(gnd), .vdd(vdd), .A(_11663_), .B(_11897_), .C(_11665_), .Y(_11898_) );
XOR2X1 XOR2X1_207 ( .gnd(gnd), .vdd(vdd), .A(_11898_), .B(_11896_), .Y(_11899_) );
OAI21X1 OAI21X1_3331 ( .gnd(gnd), .vdd(vdd), .A(_9311__bF_buf1), .B(_11899_), .C(_11895_), .Y(_11900_) );
XNOR2X1 XNOR2X1_504 ( .gnd(gnd), .vdd(vdd), .A(_11791__bF_buf2), .B(_9092_), .Y(_11901_) );
OAI21X1 OAI21X1_3332 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_133_), .B(_11537__bF_buf1), .C(_11670_), .Y(_11902_) );
OAI21X1 OAI21X1_3333 ( .gnd(gnd), .vdd(vdd), .A(_9088_), .B(_11560__bF_buf0), .C(_11902_), .Y(_11903_) );
XOR2X1 XOR2X1_208 ( .gnd(gnd), .vdd(vdd), .A(_11903_), .B(_11901_), .Y(_11904_) );
AOI21X1 AOI21X1_2011 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe40_bF_buf4), .B(_11904_), .C(micro_hash_ucr_3_pipe42_bF_buf2), .Y(_11905_) );
OAI21X1 OAI21X1_3334 ( .gnd(gnd), .vdd(vdd), .A(_11900_), .B(micro_hash_ucr_3_pipe40_bF_buf3), .C(_11905_), .Y(_11906_) );
XNOR2X1 XNOR2X1_505 ( .gnd(gnd), .vdd(vdd), .A(_11791__bF_buf1), .B(_9207_), .Y(_11907_) );
INVX1 INVX1_826 ( .gnd(gnd), .vdd(vdd), .A(_11676_), .Y(_11908_) );
OAI21X1 OAI21X1_3335 ( .gnd(gnd), .vdd(vdd), .A(_11675_), .B(_11908_), .C(_11677_), .Y(_11909_) );
XNOR2X1 XNOR2X1_506 ( .gnd(gnd), .vdd(vdd), .A(_11909_), .B(_11907_), .Y(_11910_) );
AOI21X1 AOI21X1_2012 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe42_bF_buf1), .B(_11910_), .C(micro_hash_ucr_3_pipe44_bF_buf2), .Y(_11911_) );
XNOR2X1 XNOR2X1_507 ( .gnd(gnd), .vdd(vdd), .A(_11791__bF_buf0), .B(_8955_), .Y(_11912_) );
AOI21X1 AOI21X1_2013 ( .gnd(gnd), .vdd(vdd), .A(_11684_), .B(_11683_), .C(_11685_), .Y(_11913_) );
INVX1 INVX1_827 ( .gnd(gnd), .vdd(vdd), .A(_11913_), .Y(_11914_) );
NAND2X1 NAND2X1_1556 ( .gnd(gnd), .vdd(vdd), .A(_11912_), .B(_11914_), .Y(_11915_) );
INVX1 INVX1_828 ( .gnd(gnd), .vdd(vdd), .A(_11912_), .Y(_11916_) );
AOI21X1 AOI21X1_2014 ( .gnd(gnd), .vdd(vdd), .A(_11916_), .B(_11913_), .C(_9305__bF_buf2), .Y(_11917_) );
AOI22X1 AOI22X1_82 ( .gnd(gnd), .vdd(vdd), .A(_11915_), .B(_11917_), .C(_11906_), .D(_11911_), .Y(_11918_) );
NAND2X1 NAND2X1_1557 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_158_), .B(_11791__bF_buf5), .Y(_11919_) );
OAI21X1 OAI21X1_3336 ( .gnd(gnd), .vdd(vdd), .A(_11790_), .B(_11788_), .C(_9011_), .Y(_11920_) );
AND2X2 AND2X2_746 ( .gnd(gnd), .vdd(vdd), .A(_11919_), .B(_11920_), .Y(_11921_) );
AOI21X1 AOI21X1_2015 ( .gnd(gnd), .vdd(vdd), .A(_11691_), .B(_11690_), .C(_11693_), .Y(_11922_) );
XNOR2X1 XNOR2X1_508 ( .gnd(gnd), .vdd(vdd), .A(_11922_), .B(_11921_), .Y(_11923_) );
AOI21X1 AOI21X1_2016 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe46_bF_buf4), .B(_11923_), .C(micro_hash_ucr_3_pipe48_bF_buf0), .Y(_11924_) );
OAI21X1 OAI21X1_3337 ( .gnd(gnd), .vdd(vdd), .A(_11918_), .B(micro_hash_ucr_3_pipe46_bF_buf3), .C(_11924_), .Y(_11925_) );
XNOR2X1 XNOR2X1_509 ( .gnd(gnd), .vdd(vdd), .A(_11791__bF_buf4), .B(micro_hash_ucr_3_Wx_166_), .Y(_11926_) );
AOI21X1 AOI21X1_2017 ( .gnd(gnd), .vdd(vdd), .A(_11700_), .B(_11699_), .C(_11701_), .Y(_11927_) );
XNOR2X1 XNOR2X1_510 ( .gnd(gnd), .vdd(vdd), .A(_11927_), .B(_11926_), .Y(_11928_) );
AOI21X1 AOI21X1_2018 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe48_bF_buf4), .B(_11928_), .C(micro_hash_ucr_3_pipe50_bF_buf4), .Y(_11929_) );
XNOR2X1 XNOR2X1_511 ( .gnd(gnd), .vdd(vdd), .A(_11791__bF_buf3), .B(_8854_), .Y(_11930_) );
AOI21X1 AOI21X1_2019 ( .gnd(gnd), .vdd(vdd), .A(_11708_), .B(_11707_), .C(_11709_), .Y(_11931_) );
INVX1 INVX1_829 ( .gnd(gnd), .vdd(vdd), .A(_11931_), .Y(_11932_) );
NAND2X1 NAND2X1_1558 ( .gnd(gnd), .vdd(vdd), .A(_11930_), .B(_11932_), .Y(_11933_) );
INVX1 INVX1_830 ( .gnd(gnd), .vdd(vdd), .A(_11930_), .Y(_11934_) );
AOI21X1 AOI21X1_2020 ( .gnd(gnd), .vdd(vdd), .A(_11934_), .B(_11931_), .C(_9299__bF_buf0), .Y(_11935_) );
AOI22X1 AOI22X1_83 ( .gnd(gnd), .vdd(vdd), .A(_11933_), .B(_11935_), .C(_11925_), .D(_11929_), .Y(_11936_) );
XNOR2X1 XNOR2X1_512 ( .gnd(gnd), .vdd(vdd), .A(_11791__bF_buf2), .B(_9093_), .Y(_11937_) );
INVX1 INVX1_831 ( .gnd(gnd), .vdd(vdd), .A(_11717_), .Y(_11938_) );
OAI21X1 OAI21X1_3338 ( .gnd(gnd), .vdd(vdd), .A(_11715_), .B(_11716_), .C(_11938_), .Y(_11939_) );
XOR2X1 XOR2X1_209 ( .gnd(gnd), .vdd(vdd), .A(_11939_), .B(_11937_), .Y(_11940_) );
AOI21X1 AOI21X1_2021 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe52_bF_buf3), .B(_11940_), .C(micro_hash_ucr_3_pipe54_bF_buf0), .Y(_11941_) );
OAI21X1 OAI21X1_3339 ( .gnd(gnd), .vdd(vdd), .A(_11936_), .B(micro_hash_ucr_3_pipe52_bF_buf2), .C(_11941_), .Y(_11942_) );
XNOR2X1 XNOR2X1_513 ( .gnd(gnd), .vdd(vdd), .A(_11791__bF_buf1), .B(_9062_), .Y(_11943_) );
OAI21X1 OAI21X1_3340 ( .gnd(gnd), .vdd(vdd), .A(_11544_), .B(_11545_), .C(_11547_), .Y(_11944_) );
XNOR2X1 XNOR2X1_514 ( .gnd(gnd), .vdd(vdd), .A(_11944_), .B(_11943_), .Y(_11945_) );
AOI21X1 AOI21X1_2022 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe54_bF_buf3), .B(_11945_), .C(micro_hash_ucr_3_pipe56_bF_buf4), .Y(_11946_) );
XNOR2X1 XNOR2X1_515 ( .gnd(gnd), .vdd(vdd), .A(_11791__bF_buf0), .B(_8956_), .Y(_11947_) );
AOI21X1 AOI21X1_2023 ( .gnd(gnd), .vdd(vdd), .A(_11726_), .B(_11725_), .C(_11727_), .Y(_11948_) );
INVX1 INVX1_832 ( .gnd(gnd), .vdd(vdd), .A(_11948_), .Y(_11949_) );
NAND2X1 NAND2X1_1559 ( .gnd(gnd), .vdd(vdd), .A(_11947_), .B(_11949_), .Y(_11950_) );
INVX1 INVX1_833 ( .gnd(gnd), .vdd(vdd), .A(_11947_), .Y(_11951_) );
AOI21X1 AOI21X1_2024 ( .gnd(gnd), .vdd(vdd), .A(_11951_), .B(_11948_), .C(_9293__bF_buf0), .Y(_11952_) );
AOI22X1 AOI22X1_84 ( .gnd(gnd), .vdd(vdd), .A(_11950_), .B(_11952_), .C(_11942_), .D(_11946_), .Y(_11953_) );
XNOR2X1 XNOR2X1_516 ( .gnd(gnd), .vdd(vdd), .A(_11791__bF_buf5), .B(_9012_), .Y(_11954_) );
OAI21X1 OAI21X1_3341 ( .gnd(gnd), .vdd(vdd), .A(_11733_), .B(_11734_), .C(_11736_), .Y(_11955_) );
XOR2X1 XOR2X1_210 ( .gnd(gnd), .vdd(vdd), .A(_11955_), .B(_11954_), .Y(_11956_) );
AOI21X1 AOI21X1_2025 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe58_bF_buf0), .B(_11956_), .C(micro_hash_ucr_3_pipe60_bF_buf2), .Y(_11957_) );
OAI21X1 OAI21X1_3342 ( .gnd(gnd), .vdd(vdd), .A(_11953_), .B(micro_hash_ucr_3_pipe58_bF_buf3), .C(_11957_), .Y(_11958_) );
XNOR2X1 XNOR2X1_517 ( .gnd(gnd), .vdd(vdd), .A(_11791__bF_buf4), .B(micro_hash_ucr_3_Wx_214_), .Y(_11959_) );
INVX1 INVX1_834 ( .gnd(gnd), .vdd(vdd), .A(_11745_), .Y(_11960_) );
OAI21X1 OAI21X1_3343 ( .gnd(gnd), .vdd(vdd), .A(_11742_), .B(_11744_), .C(_11960_), .Y(_11961_) );
XOR2X1 XOR2X1_211 ( .gnd(gnd), .vdd(vdd), .A(_11961_), .B(_11959_), .Y(_11962_) );
AOI21X1 AOI21X1_2026 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe60_bF_buf1), .B(_11962_), .C(micro_hash_ucr_3_pipe62_bF_buf2), .Y(_11963_) );
XNOR2X1 XNOR2X1_518 ( .gnd(gnd), .vdd(vdd), .A(_11791__bF_buf3), .B(_8855_), .Y(_11964_) );
OAI21X1 OAI21X1_3344 ( .gnd(gnd), .vdd(vdd), .A(_11749_), .B(_11750_), .C(_11752_), .Y(_11965_) );
NAND2X1 NAND2X1_1560 ( .gnd(gnd), .vdd(vdd), .A(_11964_), .B(_11965_), .Y(_11966_) );
NOR2X1 NOR2X1_1942 ( .gnd(gnd), .vdd(vdd), .A(_11964_), .B(_11965_), .Y(_11967_) );
NOR2X1 NOR2X1_1943 ( .gnd(gnd), .vdd(vdd), .A(_9287__bF_buf2), .B(_11967_), .Y(_11968_) );
AOI22X1 AOI22X1_85 ( .gnd(gnd), .vdd(vdd), .A(_11966_), .B(_11968_), .C(_11958_), .D(_11963_), .Y(_11969_) );
NAND2X1 NAND2X1_1561 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_230_), .B(_11791__bF_buf2), .Y(_11970_) );
INVX1 INVX1_835 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_230_), .Y(_11971_) );
OAI21X1 OAI21X1_3345 ( .gnd(gnd), .vdd(vdd), .A(_11790_), .B(_11788_), .C(_11971_), .Y(_11972_) );
AND2X2 AND2X2_747 ( .gnd(gnd), .vdd(vdd), .A(_11970_), .B(_11972_), .Y(_11973_) );
AOI21X1 AOI21X1_2027 ( .gnd(gnd), .vdd(vdd), .A(_11761_), .B(_11759_), .C(_11762_), .Y(_11974_) );
XNOR2X1 XNOR2X1_519 ( .gnd(gnd), .vdd(vdd), .A(_11974_), .B(_11973_), .Y(_11975_) );
AOI21X1 AOI21X1_2028 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe64_bF_buf2), .B(_11975_), .C(micro_hash_ucr_3_pipe66_bF_buf3), .Y(_11976_) );
OAI21X1 OAI21X1_3346 ( .gnd(gnd), .vdd(vdd), .A(_11969_), .B(micro_hash_ucr_3_pipe64_bF_buf1), .C(_11976_), .Y(_11977_) );
XOR2X1 XOR2X1_212 ( .gnd(gnd), .vdd(vdd), .A(_11791__bF_buf1), .B(micro_hash_ucr_3_Wx_238_), .Y(_11978_) );
OAI21X1 OAI21X1_3347 ( .gnd(gnd), .vdd(vdd), .A(_11527_), .B(_11538_), .C(_11540_), .Y(_11979_) );
NOR2X1 NOR2X1_1944 ( .gnd(gnd), .vdd(vdd), .A(_11978_), .B(_11979_), .Y(_11980_) );
AND2X2 AND2X2_748 ( .gnd(gnd), .vdd(vdd), .A(_11979_), .B(_11978_), .Y(_11981_) );
OAI21X1 OAI21X1_3348 ( .gnd(gnd), .vdd(vdd), .A(_11981_), .B(_11980_), .C(micro_hash_ucr_3_pipe66_bF_buf2), .Y(_11982_) );
AND2X2 AND2X2_749 ( .gnd(gnd), .vdd(vdd), .A(_11977_), .B(_11982_), .Y(_11983_) );
XNOR2X1 XNOR2X1_520 ( .gnd(gnd), .vdd(vdd), .A(_11791__bF_buf0), .B(micro_hash_ucr_3_Wx_246_), .Y(_11984_) );
INVX1 INVX1_836 ( .gnd(gnd), .vdd(vdd), .A(_11773_), .Y(_11985_) );
OAI21X1 OAI21X1_3349 ( .gnd(gnd), .vdd(vdd), .A(_11769_), .B(_11772_), .C(_11985_), .Y(_11986_) );
INVX1 INVX1_837 ( .gnd(gnd), .vdd(vdd), .A(_11986_), .Y(_11987_) );
AND2X2 AND2X2_750 ( .gnd(gnd), .vdd(vdd), .A(_11987_), .B(_11984_), .Y(_11988_) );
NOR2X1 NOR2X1_1945 ( .gnd(gnd), .vdd(vdd), .A(_11984_), .B(_11987_), .Y(_11989_) );
OAI21X1 OAI21X1_3350 ( .gnd(gnd), .vdd(vdd), .A(_11988_), .B(_11989_), .C(micro_hash_ucr_3_pipe68_bF_buf1), .Y(_11990_) );
OAI21X1 OAI21X1_3351 ( .gnd(gnd), .vdd(vdd), .A(_11983_), .B(micro_hash_ucr_3_pipe68_bF_buf0), .C(_11990_), .Y(_11991_) );
XNOR2X1 XNOR2X1_521 ( .gnd(gnd), .vdd(vdd), .A(_11791__bF_buf5), .B(micro_hash_ucr_3_Wx_254_), .Y(_11992_) );
AOI21X1 AOI21X1_2029 ( .gnd(gnd), .vdd(vdd), .A(_11781_), .B(_11779_), .C(_11782_), .Y(_11993_) );
AND2X2 AND2X2_751 ( .gnd(gnd), .vdd(vdd), .A(_11992_), .B(_11993_), .Y(_11994_) );
NOR2X1 NOR2X1_1946 ( .gnd(gnd), .vdd(vdd), .A(_8800__bF_buf2), .B(_11994_), .Y(_11995_) );
OAI21X1 OAI21X1_3352 ( .gnd(gnd), .vdd(vdd), .A(_11992_), .B(_11993_), .C(_11995_), .Y(_11996_) );
AOI22X1 AOI22X1_86 ( .gnd(gnd), .vdd(vdd), .A(_10381_), .B(_11996_), .C(_11991_), .D(_9283__bF_buf1), .Y(_8702__6_) );
OAI21X1 OAI21X1_3353 ( .gnd(gnd), .vdd(vdd), .A(_8855_), .B(_11852__bF_buf1), .C(_11966_), .Y(_11997_) );
NAND2X1 NAND2X1_1562 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_k_6_), .B(micro_hash_ucr_3_x_6_), .Y(_11998_) );
NAND2X1 NAND2X1_1563 ( .gnd(gnd), .vdd(vdd), .A(_11998_), .B(_11789_), .Y(_11999_) );
XOR2X1 XOR2X1_213 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_k_7_), .B(micro_hash_ucr_3_x_7_), .Y(_12000_) );
XOR2X1 XOR2X1_214 ( .gnd(gnd), .vdd(vdd), .A(_11999_), .B(_12000_), .Y(_12001_) );
XNOR2X1 XNOR2X1_522 ( .gnd(gnd), .vdd(vdd), .A(_12001__bF_buf4), .B(micro_hash_ucr_3_Wx_223_), .Y(_12002_) );
AND2X2 AND2X2_752 ( .gnd(gnd), .vdd(vdd), .A(_11997_), .B(_12002_), .Y(_12003_) );
OAI21X1 OAI21X1_3354 ( .gnd(gnd), .vdd(vdd), .A(_8956_), .B(_11852__bF_buf0), .C(_11950_), .Y(_12004_) );
XNOR2X1 XNOR2X1_523 ( .gnd(gnd), .vdd(vdd), .A(_12001__bF_buf3), .B(micro_hash_ucr_3_Wx_199_), .Y(_12005_) );
XNOR2X1 XNOR2X1_524 ( .gnd(gnd), .vdd(vdd), .A(_12004_), .B(_12005_), .Y(_12006_) );
OAI21X1 OAI21X1_3355 ( .gnd(gnd), .vdd(vdd), .A(_8955_), .B(_11852__bF_buf3), .C(_11915_), .Y(_12007_) );
XNOR2X1 XNOR2X1_525 ( .gnd(gnd), .vdd(vdd), .A(_12001__bF_buf2), .B(micro_hash_ucr_3_Wx_151_), .Y(_12008_) );
XNOR2X1 XNOR2X1_526 ( .gnd(gnd), .vdd(vdd), .A(_12007_), .B(_12008_), .Y(_12009_) );
NAND2X1 NAND2X1_1564 ( .gnd(gnd), .vdd(vdd), .A(_11889_), .B(_11891_), .Y(_12010_) );
OAI21X1 OAI21X1_3356 ( .gnd(gnd), .vdd(vdd), .A(_9132_), .B(_11852__bF_buf2), .C(_12010_), .Y(_12011_) );
XNOR2X1 XNOR2X1_527 ( .gnd(gnd), .vdd(vdd), .A(_12001__bF_buf1), .B(micro_hash_ucr_3_Wx_119_), .Y(_12012_) );
AND2X2 AND2X2_753 ( .gnd(gnd), .vdd(vdd), .A(_12011_), .B(_12012_), .Y(_12013_) );
OAI21X1 OAI21X1_3357 ( .gnd(gnd), .vdd(vdd), .A(_9232_), .B(_11852__bF_buf1), .C(_11865_), .Y(_12014_) );
XNOR2X1 XNOR2X1_528 ( .gnd(gnd), .vdd(vdd), .A(_12001__bF_buf0), .B(micro_hash_ucr_3_Wx_87_), .Y(_12015_) );
XNOR2X1 XNOR2X1_529 ( .gnd(gnd), .vdd(vdd), .A(_12014_), .B(_12015_), .Y(_12016_) );
NAND2X1 NAND2X1_1565 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_70_), .B(_11791__bF_buf4), .Y(_12017_) );
OAI21X1 OAI21X1_3358 ( .gnd(gnd), .vdd(vdd), .A(_11848_), .B(_11846_), .C(_12017_), .Y(_12018_) );
XNOR2X1 XNOR2X1_530 ( .gnd(gnd), .vdd(vdd), .A(_12001__bF_buf4), .B(_9257_), .Y(_12019_) );
XNOR2X1 XNOR2X1_531 ( .gnd(gnd), .vdd(vdd), .A(_12018_), .B(_12019_), .Y(_12020_) );
OAI21X1 OAI21X1_3359 ( .gnd(gnd), .vdd(vdd), .A(_9278_), .B(_11852__bF_buf0), .C(_11842_), .Y(_12021_) );
XNOR2X1 XNOR2X1_532 ( .gnd(gnd), .vdd(vdd), .A(_12001__bF_buf3), .B(micro_hash_ucr_3_Wx_63_), .Y(_12022_) );
XNOR2X1 XNOR2X1_533 ( .gnd(gnd), .vdd(vdd), .A(_12021_), .B(_12022_), .Y(_12023_) );
AOI21X1 AOI21X1_2030 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_6_), .B(_11791__bF_buf3), .C(_11800_), .Y(_12024_) );
XOR2X1 XOR2X1_215 ( .gnd(gnd), .vdd(vdd), .A(_12001__bF_buf2), .B(micro_hash_ucr_3_Wx_7_), .Y(_12025_) );
AOI21X1 AOI21X1_2031 ( .gnd(gnd), .vdd(vdd), .A(_12025_), .B(_12024_), .C(_9341_), .Y(_12026_) );
OAI21X1 OAI21X1_3360 ( .gnd(gnd), .vdd(vdd), .A(_12024_), .B(_12025_), .C(_12026_), .Y(_12027_) );
AND2X2 AND2X2_754 ( .gnd(gnd), .vdd(vdd), .A(H_3_23_), .B(micro_hash_ucr_3_pipe6_bF_buf1), .Y(_12028_) );
INVX1 INVX1_838 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_7_), .Y(_12029_) );
OAI21X1 OAI21X1_3361 ( .gnd(gnd), .vdd(vdd), .A(_12029_), .B(micro_hash_ucr_3_pipe6_bF_buf0), .C(_9341_), .Y(_12030_) );
OAI21X1 OAI21X1_3362 ( .gnd(gnd), .vdd(vdd), .A(_12028_), .B(_12030_), .C(_12027_), .Y(_12031_) );
INVX1 INVX1_839 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_14_), .Y(_12032_) );
NAND2X1 NAND2X1_1566 ( .gnd(gnd), .vdd(vdd), .A(_11792_), .B(_11793_), .Y(_12033_) );
OAI21X1 OAI21X1_3363 ( .gnd(gnd), .vdd(vdd), .A(_12032_), .B(_11852__bF_buf3), .C(_12033_), .Y(_12034_) );
XNOR2X1 XNOR2X1_534 ( .gnd(gnd), .vdd(vdd), .A(_12001__bF_buf1), .B(micro_hash_ucr_3_Wx_15_), .Y(_12035_) );
XNOR2X1 XNOR2X1_535 ( .gnd(gnd), .vdd(vdd), .A(_12034_), .B(_12035_), .Y(_12036_) );
AOI21X1 AOI21X1_2032 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe10_bF_buf0), .B(_12036_), .C(micro_hash_ucr_3_pipe12), .Y(_12037_) );
OAI21X1 OAI21X1_3364 ( .gnd(gnd), .vdd(vdd), .A(_12031_), .B(micro_hash_ucr_3_pipe10_bF_buf3), .C(_12037_), .Y(_12038_) );
OAI21X1 OAI21X1_3365 ( .gnd(gnd), .vdd(vdd), .A(_11804_), .B(_11852__bF_buf2), .C(_11808_), .Y(_12039_) );
XNOR2X1 XNOR2X1_536 ( .gnd(gnd), .vdd(vdd), .A(_12001__bF_buf0), .B(micro_hash_ucr_3_Wx_23_), .Y(_12040_) );
AOI21X1 AOI21X1_2033 ( .gnd(gnd), .vdd(vdd), .A(_12040_), .B(_12039_), .C(_9340_), .Y(_12041_) );
OAI21X1 OAI21X1_3366 ( .gnd(gnd), .vdd(vdd), .A(_12039_), .B(_12040_), .C(_12041_), .Y(_12042_) );
NAND3X1 NAND3X1_599 ( .gnd(gnd), .vdd(vdd), .A(_9335__bF_buf2), .B(_12042_), .C(_12038_), .Y(_12043_) );
NAND2X1 NAND2X1_1567 ( .gnd(gnd), .vdd(vdd), .A(_11814_), .B(_11815_), .Y(_12044_) );
OAI21X1 OAI21X1_3367 ( .gnd(gnd), .vdd(vdd), .A(_11813_), .B(_11852__bF_buf1), .C(_12044_), .Y(_12045_) );
XNOR2X1 XNOR2X1_537 ( .gnd(gnd), .vdd(vdd), .A(_12001__bF_buf4), .B(micro_hash_ucr_3_Wx_31_), .Y(_12046_) );
XNOR2X1 XNOR2X1_538 ( .gnd(gnd), .vdd(vdd), .A(_12045_), .B(_12046_), .Y(_12047_) );
AOI21X1 AOI21X1_2034 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe14_bF_buf2), .B(_12047_), .C(micro_hash_ucr_3_pipe16_bF_buf2), .Y(_12048_) );
INVX1 INVX1_840 ( .gnd(gnd), .vdd(vdd), .A(_11821_), .Y(_12049_) );
OAI21X1 OAI21X1_3368 ( .gnd(gnd), .vdd(vdd), .A(_11822_), .B(_12049_), .C(_11818_), .Y(_12050_) );
XNOR2X1 XNOR2X1_539 ( .gnd(gnd), .vdd(vdd), .A(_12001__bF_buf3), .B(micro_hash_ucr_3_Wx_39_), .Y(_12051_) );
OAI21X1 OAI21X1_3369 ( .gnd(gnd), .vdd(vdd), .A(_12050_), .B(_12051_), .C(micro_hash_ucr_3_pipe16_bF_buf1), .Y(_12052_) );
AOI21X1 AOI21X1_2035 ( .gnd(gnd), .vdd(vdd), .A(_12050_), .B(_12051_), .C(_12052_), .Y(_12053_) );
AOI21X1 AOI21X1_2036 ( .gnd(gnd), .vdd(vdd), .A(_12048_), .B(_12043_), .C(_12053_), .Y(_12054_) );
OAI21X1 OAI21X1_3370 ( .gnd(gnd), .vdd(vdd), .A(_11825_), .B(_11852__bF_buf0), .C(_11829_), .Y(_12055_) );
XOR2X1 XOR2X1_216 ( .gnd(gnd), .vdd(vdd), .A(_12001__bF_buf2), .B(micro_hash_ucr_3_Wx_47_), .Y(_12056_) );
XNOR2X1 XNOR2X1_540 ( .gnd(gnd), .vdd(vdd), .A(_12055_), .B(_12056_), .Y(_12057_) );
OAI21X1 OAI21X1_3371 ( .gnd(gnd), .vdd(vdd), .A(_12057_), .B(_9334__bF_buf2), .C(_9329__bF_buf4), .Y(_12058_) );
AOI21X1 AOI21X1_2037 ( .gnd(gnd), .vdd(vdd), .A(_9334__bF_buf1), .B(_12054_), .C(_12058_), .Y(_12059_) );
NAND2X1 NAND2X1_1568 ( .gnd(gnd), .vdd(vdd), .A(_11833_), .B(_11834_), .Y(_12060_) );
OAI21X1 OAI21X1_3372 ( .gnd(gnd), .vdd(vdd), .A(_11832_), .B(_11852__bF_buf3), .C(_12060_), .Y(_12061_) );
XNOR2X1 XNOR2X1_541 ( .gnd(gnd), .vdd(vdd), .A(_12001__bF_buf1), .B(micro_hash_ucr_3_Wx_55_), .Y(_12062_) );
OAI21X1 OAI21X1_3373 ( .gnd(gnd), .vdd(vdd), .A(_12061_), .B(_12062_), .C(micro_hash_ucr_3_pipe20_bF_buf1), .Y(_12063_) );
AOI21X1 AOI21X1_2038 ( .gnd(gnd), .vdd(vdd), .A(_12061_), .B(_12062_), .C(_12063_), .Y(_12064_) );
OAI21X1 OAI21X1_3374 ( .gnd(gnd), .vdd(vdd), .A(_12059_), .B(_12064_), .C(_9330__bF_buf4), .Y(_12065_) );
OAI21X1 OAI21X1_3375 ( .gnd(gnd), .vdd(vdd), .A(_9330__bF_buf3), .B(_12023_), .C(_12065_), .Y(_12066_) );
MUX2X1 MUX2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_12066_), .B(_12020_), .S(_9328__bF_buf1), .Y(_12067_) );
AOI21X1 AOI21X1_2039 ( .gnd(gnd), .vdd(vdd), .A(_11855_), .B(_11858_), .C(_11853_), .Y(_12068_) );
XNOR2X1 XNOR2X1_542 ( .gnd(gnd), .vdd(vdd), .A(_12001__bF_buf0), .B(_9135_), .Y(_12069_) );
AOI21X1 AOI21X1_2040 ( .gnd(gnd), .vdd(vdd), .A(_12069_), .B(_12068_), .C(_9323__bF_buf3), .Y(_12070_) );
OAI21X1 OAI21X1_3376 ( .gnd(gnd), .vdd(vdd), .A(_12068_), .B(_12069_), .C(_12070_), .Y(_12071_) );
OAI21X1 OAI21X1_3377 ( .gnd(gnd), .vdd(vdd), .A(_12067_), .B(micro_hash_ucr_3_pipe26_bF_buf3), .C(_12071_), .Y(_12072_) );
NAND2X1 NAND2X1_1569 ( .gnd(gnd), .vdd(vdd), .A(_9324__bF_buf3), .B(_12072_), .Y(_12073_) );
OAI21X1 OAI21X1_3378 ( .gnd(gnd), .vdd(vdd), .A(_9324__bF_buf2), .B(_12016_), .C(_12073_), .Y(_12074_) );
NAND2X1 NAND2X1_1570 ( .gnd(gnd), .vdd(vdd), .A(_11870_), .B(_11872_), .Y(_12075_) );
OAI21X1 OAI21X1_3379 ( .gnd(gnd), .vdd(vdd), .A(_9206_), .B(_11852__bF_buf2), .C(_12075_), .Y(_12076_) );
XNOR2X1 XNOR2X1_543 ( .gnd(gnd), .vdd(vdd), .A(_12001__bF_buf4), .B(micro_hash_ucr_3_Wx_95_), .Y(_12077_) );
XNOR2X1 XNOR2X1_544 ( .gnd(gnd), .vdd(vdd), .A(_12076_), .B(_12077_), .Y(_12078_) );
OAI21X1 OAI21X1_3380 ( .gnd(gnd), .vdd(vdd), .A(_12078_), .B(_9322__bF_buf0), .C(_9317__bF_buf2), .Y(_12079_) );
AOI21X1 AOI21X1_2041 ( .gnd(gnd), .vdd(vdd), .A(_9322__bF_buf3), .B(_12074_), .C(_12079_), .Y(_12080_) );
NAND2X1 NAND2X1_1571 ( .gnd(gnd), .vdd(vdd), .A(_11875_), .B(_11877_), .Y(_12081_) );
OAI21X1 OAI21X1_3381 ( .gnd(gnd), .vdd(vdd), .A(_9061_), .B(_11852__bF_buf1), .C(_12081_), .Y(_12082_) );
XNOR2X1 XNOR2X1_545 ( .gnd(gnd), .vdd(vdd), .A(_12001__bF_buf3), .B(_9065_), .Y(_12083_) );
XNOR2X1 XNOR2X1_546 ( .gnd(gnd), .vdd(vdd), .A(_12082_), .B(_12083_), .Y(_12084_) );
OAI21X1 OAI21X1_3382 ( .gnd(gnd), .vdd(vdd), .A(_12084_), .B(_9317__bF_buf1), .C(_9318__bF_buf4), .Y(_12085_) );
AOI21X1 AOI21X1_2042 ( .gnd(gnd), .vdd(vdd), .A(_11883_), .B(_11886_), .C(_11881_), .Y(_12086_) );
XNOR2X1 XNOR2X1_547 ( .gnd(gnd), .vdd(vdd), .A(_12001__bF_buf2), .B(_8959_), .Y(_12087_) );
AOI21X1 AOI21X1_2043 ( .gnd(gnd), .vdd(vdd), .A(_12087_), .B(_12086_), .C(_9318__bF_buf3), .Y(_12088_) );
OAI21X1 OAI21X1_3383 ( .gnd(gnd), .vdd(vdd), .A(_12086_), .B(_12087_), .C(_12088_), .Y(_12089_) );
OAI21X1 OAI21X1_3384 ( .gnd(gnd), .vdd(vdd), .A(_12080_), .B(_12085_), .C(_12089_), .Y(_12090_) );
NAND2X1 NAND2X1_1572 ( .gnd(gnd), .vdd(vdd), .A(_9316__bF_buf0), .B(_12090_), .Y(_12091_) );
OAI21X1 OAI21X1_3385 ( .gnd(gnd), .vdd(vdd), .A(_12011_), .B(_12012_), .C(micro_hash_ucr_3_pipe36_bF_buf3), .Y(_12092_) );
OAI21X1 OAI21X1_3386 ( .gnd(gnd), .vdd(vdd), .A(_12013_), .B(_12092_), .C(_12091_), .Y(_12093_) );
NAND2X1 NAND2X1_1573 ( .gnd(gnd), .vdd(vdd), .A(_11896_), .B(_11898_), .Y(_12094_) );
OAI21X1 OAI21X1_3387 ( .gnd(gnd), .vdd(vdd), .A(_8985_), .B(_11852__bF_buf0), .C(_12094_), .Y(_12095_) );
XNOR2X1 XNOR2X1_548 ( .gnd(gnd), .vdd(vdd), .A(_12001__bF_buf1), .B(micro_hash_ucr_3_Wx_127_), .Y(_12096_) );
OAI21X1 OAI21X1_3388 ( .gnd(gnd), .vdd(vdd), .A(_12095_), .B(_12096_), .C(micro_hash_ucr_3_pipe38_bF_buf2), .Y(_12097_) );
AOI21X1 AOI21X1_2044 ( .gnd(gnd), .vdd(vdd), .A(_12095_), .B(_12096_), .C(_12097_), .Y(_12098_) );
AOI21X1 AOI21X1_2045 ( .gnd(gnd), .vdd(vdd), .A(_9311__bF_buf0), .B(_12093_), .C(_12098_), .Y(_12099_) );
NAND2X1 NAND2X1_1574 ( .gnd(gnd), .vdd(vdd), .A(_11901_), .B(_11903_), .Y(_12100_) );
OAI21X1 OAI21X1_3389 ( .gnd(gnd), .vdd(vdd), .A(_9092_), .B(_11852__bF_buf3), .C(_12100_), .Y(_12101_) );
XOR2X1 XOR2X1_217 ( .gnd(gnd), .vdd(vdd), .A(_12001__bF_buf0), .B(micro_hash_ucr_3_Wx_135_), .Y(_12102_) );
XNOR2X1 XNOR2X1_549 ( .gnd(gnd), .vdd(vdd), .A(_12101_), .B(_12102_), .Y(_12103_) );
OAI21X1 OAI21X1_3390 ( .gnd(gnd), .vdd(vdd), .A(_12103_), .B(_9312__bF_buf1), .C(_9310__bF_buf2), .Y(_12104_) );
AOI21X1 AOI21X1_2046 ( .gnd(gnd), .vdd(vdd), .A(_9312__bF_buf0), .B(_12099_), .C(_12104_), .Y(_12105_) );
NAND2X1 NAND2X1_1575 ( .gnd(gnd), .vdd(vdd), .A(_11907_), .B(_11909_), .Y(_12106_) );
OAI21X1 OAI21X1_3391 ( .gnd(gnd), .vdd(vdd), .A(_9207_), .B(_11852__bF_buf2), .C(_12106_), .Y(_12107_) );
XNOR2X1 XNOR2X1_550 ( .gnd(gnd), .vdd(vdd), .A(_12001__bF_buf4), .B(micro_hash_ucr_3_Wx_143_), .Y(_12108_) );
OAI21X1 OAI21X1_3392 ( .gnd(gnd), .vdd(vdd), .A(_12107_), .B(_12108_), .C(micro_hash_ucr_3_pipe42_bF_buf0), .Y(_12109_) );
AOI21X1 AOI21X1_2047 ( .gnd(gnd), .vdd(vdd), .A(_12107_), .B(_12108_), .C(_12109_), .Y(_12110_) );
OAI21X1 OAI21X1_3393 ( .gnd(gnd), .vdd(vdd), .A(_12105_), .B(_12110_), .C(_9305__bF_buf1), .Y(_12111_) );
OAI21X1 OAI21X1_3394 ( .gnd(gnd), .vdd(vdd), .A(_9305__bF_buf0), .B(_12009_), .C(_12111_), .Y(_12112_) );
INVX1 INVX1_841 ( .gnd(gnd), .vdd(vdd), .A(_11921_), .Y(_12113_) );
OAI21X1 OAI21X1_3395 ( .gnd(gnd), .vdd(vdd), .A(_11922_), .B(_12113_), .C(_11919_), .Y(_12114_) );
XNOR2X1 XNOR2X1_551 ( .gnd(gnd), .vdd(vdd), .A(_12001__bF_buf3), .B(_9015_), .Y(_12115_) );
XNOR2X1 XNOR2X1_552 ( .gnd(gnd), .vdd(vdd), .A(_12114_), .B(_12115_), .Y(_12116_) );
MUX2X1 MUX2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_12112_), .B(_12116_), .S(_9306__bF_buf0), .Y(_12117_) );
NOR2X1 NOR2X1_1947 ( .gnd(gnd), .vdd(vdd), .A(_11926_), .B(_11927_), .Y(_12118_) );
AOI21X1 AOI21X1_2048 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_166_), .B(_11791__bF_buf2), .C(_12118_), .Y(_12119_) );
XNOR2X1 XNOR2X1_553 ( .gnd(gnd), .vdd(vdd), .A(_12001__bF_buf2), .B(_8988_), .Y(_12120_) );
AOI21X1 AOI21X1_2049 ( .gnd(gnd), .vdd(vdd), .A(_12120_), .B(_12119_), .C(_9304__bF_buf3), .Y(_12121_) );
OAI21X1 OAI21X1_3396 ( .gnd(gnd), .vdd(vdd), .A(_12119_), .B(_12120_), .C(_12121_), .Y(_12122_) );
OAI21X1 OAI21X1_3397 ( .gnd(gnd), .vdd(vdd), .A(_12117_), .B(micro_hash_ucr_3_pipe48_bF_buf3), .C(_12122_), .Y(_12123_) );
OAI21X1 OAI21X1_3398 ( .gnd(gnd), .vdd(vdd), .A(_8854_), .B(_11852__bF_buf1), .C(_11933_), .Y(_12124_) );
XNOR2X1 XNOR2X1_554 ( .gnd(gnd), .vdd(vdd), .A(_12001__bF_buf1), .B(micro_hash_ucr_3_Wx_175_), .Y(_12125_) );
OAI21X1 OAI21X1_3399 ( .gnd(gnd), .vdd(vdd), .A(_12124_), .B(_12125_), .C(micro_hash_ucr_3_pipe50_bF_buf3), .Y(_12126_) );
AOI21X1 AOI21X1_2050 ( .gnd(gnd), .vdd(vdd), .A(_12124_), .B(_12125_), .C(_12126_), .Y(_12127_) );
AOI21X1 AOI21X1_2051 ( .gnd(gnd), .vdd(vdd), .A(_9299__bF_buf3), .B(_12123_), .C(_12127_), .Y(_12128_) );
NAND2X1 NAND2X1_1576 ( .gnd(gnd), .vdd(vdd), .A(_11937_), .B(_11939_), .Y(_12129_) );
OAI21X1 OAI21X1_3400 ( .gnd(gnd), .vdd(vdd), .A(_9093_), .B(_11852__bF_buf0), .C(_12129_), .Y(_12130_) );
XNOR2X1 XNOR2X1_555 ( .gnd(gnd), .vdd(vdd), .A(_12001__bF_buf0), .B(_9096_), .Y(_12131_) );
XNOR2X1 XNOR2X1_556 ( .gnd(gnd), .vdd(vdd), .A(_12130_), .B(_12131_), .Y(_12132_) );
OAI21X1 OAI21X1_3401 ( .gnd(gnd), .vdd(vdd), .A(_12132_), .B(_9300__bF_buf1), .C(_9298__bF_buf0), .Y(_12133_) );
AOI21X1 AOI21X1_2052 ( .gnd(gnd), .vdd(vdd), .A(_9300__bF_buf0), .B(_12128_), .C(_12133_), .Y(_12134_) );
NAND2X1 NAND2X1_1577 ( .gnd(gnd), .vdd(vdd), .A(_11943_), .B(_11944_), .Y(_12135_) );
OAI21X1 OAI21X1_3402 ( .gnd(gnd), .vdd(vdd), .A(_9062_), .B(_11852__bF_buf3), .C(_12135_), .Y(_12136_) );
XNOR2X1 XNOR2X1_557 ( .gnd(gnd), .vdd(vdd), .A(_12001__bF_buf4), .B(micro_hash_ucr_3_Wx_191_), .Y(_12137_) );
OAI21X1 OAI21X1_3403 ( .gnd(gnd), .vdd(vdd), .A(_12136_), .B(_12137_), .C(micro_hash_ucr_3_pipe54_bF_buf2), .Y(_12138_) );
AOI21X1 AOI21X1_2053 ( .gnd(gnd), .vdd(vdd), .A(_12136_), .B(_12137_), .C(_12138_), .Y(_12139_) );
OAI21X1 OAI21X1_3404 ( .gnd(gnd), .vdd(vdd), .A(_12134_), .B(_12139_), .C(_9293__bF_buf3), .Y(_12140_) );
OAI21X1 OAI21X1_3405 ( .gnd(gnd), .vdd(vdd), .A(_9293__bF_buf2), .B(_12006_), .C(_12140_), .Y(_12141_) );
NAND2X1 NAND2X1_1578 ( .gnd(gnd), .vdd(vdd), .A(_11954_), .B(_11955_), .Y(_12142_) );
OAI21X1 OAI21X1_3406 ( .gnd(gnd), .vdd(vdd), .A(_9012_), .B(_11852__bF_buf2), .C(_12142_), .Y(_12143_) );
XOR2X1 XOR2X1_218 ( .gnd(gnd), .vdd(vdd), .A(_12001__bF_buf3), .B(micro_hash_ucr_3_Wx_207_), .Y(_12144_) );
XNOR2X1 XNOR2X1_558 ( .gnd(gnd), .vdd(vdd), .A(_12143_), .B(_12144_), .Y(_12145_) );
MUX2X1 MUX2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_12141_), .B(_12145_), .S(_9294__bF_buf4), .Y(_12146_) );
INVX1 INVX1_842 ( .gnd(gnd), .vdd(vdd), .A(_11961_), .Y(_12147_) );
NOR2X1 NOR2X1_1948 ( .gnd(gnd), .vdd(vdd), .A(_11959_), .B(_12147_), .Y(_12148_) );
AOI21X1 AOI21X1_2054 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_214_), .B(_11791__bF_buf1), .C(_12148_), .Y(_12149_) );
XOR2X1 XOR2X1_219 ( .gnd(gnd), .vdd(vdd), .A(_12001__bF_buf2), .B(micro_hash_ucr_3_Wx_215_), .Y(_12150_) );
AOI21X1 AOI21X1_2055 ( .gnd(gnd), .vdd(vdd), .A(_12150_), .B(_12149_), .C(_9292__bF_buf2), .Y(_12151_) );
OAI21X1 OAI21X1_3407 ( .gnd(gnd), .vdd(vdd), .A(_12149_), .B(_12150_), .C(_12151_), .Y(_12152_) );
OAI21X1 OAI21X1_3408 ( .gnd(gnd), .vdd(vdd), .A(_12146_), .B(micro_hash_ucr_3_pipe60_bF_buf0), .C(_12152_), .Y(_12153_) );
NAND2X1 NAND2X1_1579 ( .gnd(gnd), .vdd(vdd), .A(_9287__bF_buf1), .B(_12153_), .Y(_12154_) );
OAI21X1 OAI21X1_3409 ( .gnd(gnd), .vdd(vdd), .A(_11997_), .B(_12002_), .C(micro_hash_ucr_3_pipe62_bF_buf1), .Y(_12155_) );
OAI21X1 OAI21X1_3410 ( .gnd(gnd), .vdd(vdd), .A(_12003_), .B(_12155_), .C(_12154_), .Y(_12156_) );
INVX1 INVX1_843 ( .gnd(gnd), .vdd(vdd), .A(_11973_), .Y(_12157_) );
OAI21X1 OAI21X1_3411 ( .gnd(gnd), .vdd(vdd), .A(_11974_), .B(_12157_), .C(_11970_), .Y(_12158_) );
XNOR2X1 XNOR2X1_559 ( .gnd(gnd), .vdd(vdd), .A(_12001__bF_buf1), .B(micro_hash_ucr_3_Wx_231_), .Y(_12159_) );
AND2X2 AND2X2_755 ( .gnd(gnd), .vdd(vdd), .A(_12158_), .B(_12159_), .Y(_12160_) );
OAI21X1 OAI21X1_3412 ( .gnd(gnd), .vdd(vdd), .A(_12158_), .B(_12159_), .C(micro_hash_ucr_3_pipe64_bF_buf0), .Y(_12161_) );
OAI21X1 OAI21X1_3413 ( .gnd(gnd), .vdd(vdd), .A(_12160_), .B(_12161_), .C(_9286__bF_buf1), .Y(_12162_) );
AOI21X1 AOI21X1_2056 ( .gnd(gnd), .vdd(vdd), .A(_9288__bF_buf2), .B(_12156_), .C(_12162_), .Y(_12163_) );
AOI21X1 AOI21X1_2057 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_238_), .B(_11791__bF_buf0), .C(_11981_), .Y(_12164_) );
XNOR2X1 XNOR2X1_560 ( .gnd(gnd), .vdd(vdd), .A(_12001__bF_buf0), .B(micro_hash_ucr_3_Wx_239_), .Y(_12165_) );
AND2X2 AND2X2_756 ( .gnd(gnd), .vdd(vdd), .A(_12164_), .B(_12165_), .Y(_12166_) );
OAI21X1 OAI21X1_3414 ( .gnd(gnd), .vdd(vdd), .A(_12164_), .B(_12165_), .C(micro_hash_ucr_3_pipe66_bF_buf1), .Y(_12167_) );
OAI21X1 OAI21X1_3415 ( .gnd(gnd), .vdd(vdd), .A(_12166_), .B(_12167_), .C(_9282__bF_buf3), .Y(_12168_) );
AOI21X1 AOI21X1_2058 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_246_), .B(_11791__bF_buf5), .C(_11989_), .Y(_12169_) );
XOR2X1 XOR2X1_220 ( .gnd(gnd), .vdd(vdd), .A(_12001__bF_buf4), .B(micro_hash_ucr_3_Wx_247_), .Y(_12170_) );
AOI21X1 AOI21X1_2059 ( .gnd(gnd), .vdd(vdd), .A(_12170_), .B(_12169_), .C(_9282__bF_buf2), .Y(_12171_) );
OAI21X1 OAI21X1_3416 ( .gnd(gnd), .vdd(vdd), .A(_12169_), .B(_12170_), .C(_12171_), .Y(_12172_) );
OAI21X1 OAI21X1_3417 ( .gnd(gnd), .vdd(vdd), .A(_12163_), .B(_12168_), .C(_12172_), .Y(_12173_) );
NAND2X1 NAND2X1_1580 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_254_), .B(_11791__bF_buf4), .Y(_12174_) );
OAI21X1 OAI21X1_3418 ( .gnd(gnd), .vdd(vdd), .A(_11992_), .B(_11993_), .C(_12174_), .Y(_12175_) );
XNOR2X1 XNOR2X1_561 ( .gnd(gnd), .vdd(vdd), .A(_12001__bF_buf3), .B(micro_hash_ucr_3_Wx_255_), .Y(_12176_) );
AND2X2 AND2X2_757 ( .gnd(gnd), .vdd(vdd), .A(_12175_), .B(_12176_), .Y(_12177_) );
OAI21X1 OAI21X1_3419 ( .gnd(gnd), .vdd(vdd), .A(_12175_), .B(_12176_), .C(micro_hash_ucr_3_pipe69), .Y(_12178_) );
OAI21X1 OAI21X1_3420 ( .gnd(gnd), .vdd(vdd), .A(_12177_), .B(_12178_), .C(_8705__bF_buf2), .Y(_12179_) );
AOI21X1 AOI21X1_2060 ( .gnd(gnd), .vdd(vdd), .A(_9283__bF_buf0), .B(_12173_), .C(_12179_), .Y(_8702__7_) );
INVX2 INVX2_392 ( .gnd(gnd), .vdd(vdd), .A(_9371_), .Y(_12180_) );
OAI21X1 OAI21X1_3421 ( .gnd(gnd), .vdd(vdd), .A(_12899_), .B(_9372_), .C(_12180_), .Y(_12181_) );
OAI21X1 OAI21X1_3422 ( .gnd(gnd), .vdd(vdd), .A(_9340_), .B(micro_hash_ucr_3_pipe13), .C(_9335__bF_buf1), .Y(_12182_) );
AOI21X1 AOI21X1_2061 ( .gnd(gnd), .vdd(vdd), .A(_9366_), .B(_12181_), .C(_12182_), .Y(_12183_) );
NAND3X1 NAND3X1_600 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe6_bF_buf3), .B(_9335__bF_buf0), .C(_9340_), .Y(_12184_) );
NOR2X1 NOR2X1_1949 ( .gnd(gnd), .vdd(vdd), .A(_9374_), .B(_12184_), .Y(_12185_) );
OAI21X1 OAI21X1_3423 ( .gnd(gnd), .vdd(vdd), .A(_12185_), .B(micro_hash_ucr_3_b_0_bF_buf3_), .C(_9337_), .Y(_12186_) );
OAI21X1 OAI21X1_3424 ( .gnd(gnd), .vdd(vdd), .A(_12183_), .B(_12186_), .C(_9336__bF_buf3), .Y(_12187_) );
AOI21X1 AOI21X1_2062 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe16_bF_buf0), .B(_12902_), .C(micro_hash_ucr_3_pipe17_bF_buf0), .Y(_12188_) );
AOI21X1 AOI21X1_2063 ( .gnd(gnd), .vdd(vdd), .A(_12188_), .B(_12187_), .C(micro_hash_ucr_3_pipe18_bF_buf4), .Y(_12189_) );
OAI21X1 OAI21X1_3425 ( .gnd(gnd), .vdd(vdd), .A(_9334__bF_buf0), .B(micro_hash_ucr_3_b_0_bF_buf2_), .C(_9333__bF_buf3), .Y(_12190_) );
OAI21X1 OAI21X1_3426 ( .gnd(gnd), .vdd(vdd), .A(_12189_), .B(_12190_), .C(_9329__bF_buf3), .Y(_12191_) );
AOI21X1 AOI21X1_2064 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe20_bF_buf0), .B(_12902_), .C(micro_hash_ucr_3_pipe21_bF_buf3), .Y(_12192_) );
AOI21X1 AOI21X1_2065 ( .gnd(gnd), .vdd(vdd), .A(_12192_), .B(_12191_), .C(micro_hash_ucr_3_pipe22_bF_buf1), .Y(_12193_) );
OAI21X1 OAI21X1_3427 ( .gnd(gnd), .vdd(vdd), .A(_9330__bF_buf2), .B(micro_hash_ucr_3_b_0_bF_buf1_), .C(_9326__bF_buf0), .Y(_12194_) );
OAI21X1 OAI21X1_3428 ( .gnd(gnd), .vdd(vdd), .A(_12193_), .B(_12194_), .C(_9328__bF_buf0), .Y(_12195_) );
AOI21X1 AOI21X1_2066 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe24_bF_buf0), .B(_12902_), .C(micro_hash_ucr_3_pipe25_bF_buf0), .Y(_12196_) );
AOI21X1 AOI21X1_2067 ( .gnd(gnd), .vdd(vdd), .A(_12196_), .B(_12195_), .C(micro_hash_ucr_3_pipe26_bF_buf2), .Y(_12197_) );
OAI21X1 OAI21X1_3429 ( .gnd(gnd), .vdd(vdd), .A(_9323__bF_buf2), .B(micro_hash_ucr_3_b_0_bF_buf0_), .C(_9325__bF_buf0), .Y(_12198_) );
OAI21X1 OAI21X1_3430 ( .gnd(gnd), .vdd(vdd), .A(_12197_), .B(_12198_), .C(_9324__bF_buf1), .Y(_12199_) );
AOI21X1 AOI21X1_2068 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe28_bF_buf3), .B(_12902_), .C(micro_hash_ucr_3_pipe29_bF_buf3), .Y(_12200_) );
AOI21X1 AOI21X1_2069 ( .gnd(gnd), .vdd(vdd), .A(_12200_), .B(_12199_), .C(micro_hash_ucr_3_pipe30_bF_buf3), .Y(_12201_) );
OAI21X1 OAI21X1_3431 ( .gnd(gnd), .vdd(vdd), .A(_9322__bF_buf2), .B(micro_hash_ucr_3_b_0_bF_buf3_), .C(_9321__bF_buf1), .Y(_12202_) );
OAI21X1 OAI21X1_3432 ( .gnd(gnd), .vdd(vdd), .A(_12201_), .B(_12202_), .C(_9317__bF_buf0), .Y(_12203_) );
AOI21X1 AOI21X1_2070 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe32_bF_buf1), .B(_12902_), .C(micro_hash_ucr_3_pipe33_bF_buf2), .Y(_12204_) );
AOI21X1 AOI21X1_2071 ( .gnd(gnd), .vdd(vdd), .A(_12204_), .B(_12203_), .C(micro_hash_ucr_3_pipe34_bF_buf2), .Y(_12205_) );
OAI21X1 OAI21X1_3433 ( .gnd(gnd), .vdd(vdd), .A(_9318__bF_buf2), .B(micro_hash_ucr_3_b_0_bF_buf2_), .C(_9314_), .Y(_12206_) );
OAI21X1 OAI21X1_3434 ( .gnd(gnd), .vdd(vdd), .A(_12205_), .B(_12206_), .C(_9316__bF_buf3), .Y(_12207_) );
AOI21X1 AOI21X1_2072 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe36_bF_buf2), .B(_12902_), .C(micro_hash_ucr_3_pipe37_bF_buf2), .Y(_12208_) );
AOI21X1 AOI21X1_2073 ( .gnd(gnd), .vdd(vdd), .A(_12208_), .B(_12207_), .C(micro_hash_ucr_3_pipe38_bF_buf1), .Y(_12209_) );
OAI21X1 OAI21X1_3435 ( .gnd(gnd), .vdd(vdd), .A(_9311__bF_buf4), .B(micro_hash_ucr_3_b_0_bF_buf1_), .C(_9313_), .Y(_12210_) );
OAI21X1 OAI21X1_3436 ( .gnd(gnd), .vdd(vdd), .A(_12209_), .B(_12210_), .C(_9312__bF_buf3), .Y(_12211_) );
AOI21X1 AOI21X1_2074 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe40_bF_buf2), .B(_12902_), .C(micro_hash_ucr_3_pipe41_bF_buf2), .Y(_12212_) );
AOI21X1 AOI21X1_2075 ( .gnd(gnd), .vdd(vdd), .A(_12212_), .B(_12211_), .C(micro_hash_ucr_3_pipe42_bF_buf3), .Y(_12213_) );
OAI21X1 OAI21X1_3437 ( .gnd(gnd), .vdd(vdd), .A(_9310__bF_buf1), .B(micro_hash_ucr_3_b_0_bF_buf0_), .C(_9309__bF_buf2), .Y(_12214_) );
OAI21X1 OAI21X1_3438 ( .gnd(gnd), .vdd(vdd), .A(_12213_), .B(_12214_), .C(_9305__bF_buf4), .Y(_12215_) );
AOI21X1 AOI21X1_2076 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe44_bF_buf1), .B(_12902_), .C(micro_hash_ucr_3_pipe45_bF_buf1), .Y(_12216_) );
AOI21X1 AOI21X1_2077 ( .gnd(gnd), .vdd(vdd), .A(_12216_), .B(_12215_), .C(micro_hash_ucr_3_pipe46_bF_buf2), .Y(_12217_) );
OAI21X1 OAI21X1_3439 ( .gnd(gnd), .vdd(vdd), .A(_9306__bF_buf3), .B(micro_hash_ucr_3_b_0_bF_buf3_), .C(_9302_), .Y(_12218_) );
OAI21X1 OAI21X1_3440 ( .gnd(gnd), .vdd(vdd), .A(_12217_), .B(_12218_), .C(_9304__bF_buf2), .Y(_12219_) );
AOI21X1 AOI21X1_2078 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe48_bF_buf2), .B(_12902_), .C(micro_hash_ucr_3_pipe49_bF_buf1), .Y(_12220_) );
AOI21X1 AOI21X1_2079 ( .gnd(gnd), .vdd(vdd), .A(_12220_), .B(_12219_), .C(micro_hash_ucr_3_pipe50_bF_buf2), .Y(_12221_) );
OAI21X1 OAI21X1_3441 ( .gnd(gnd), .vdd(vdd), .A(_9299__bF_buf2), .B(micro_hash_ucr_3_b_0_bF_buf2_), .C(_9301__bF_buf1), .Y(_12222_) );
OAI21X1 OAI21X1_3442 ( .gnd(gnd), .vdd(vdd), .A(_12221_), .B(_12222_), .C(_9300__bF_buf3), .Y(_12223_) );
AOI21X1 AOI21X1_2080 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe52_bF_buf1), .B(_12902_), .C(micro_hash_ucr_3_pipe53), .Y(_12224_) );
AOI21X1 AOI21X1_2081 ( .gnd(gnd), .vdd(vdd), .A(_12224_), .B(_12223_), .C(micro_hash_ucr_3_pipe54_bF_buf1), .Y(_12225_) );
OAI21X1 OAI21X1_3443 ( .gnd(gnd), .vdd(vdd), .A(_9298__bF_buf4), .B(micro_hash_ucr_3_b_0_bF_buf1_), .C(_9297_), .Y(_12226_) );
OAI21X1 OAI21X1_3444 ( .gnd(gnd), .vdd(vdd), .A(_12225_), .B(_12226_), .C(_9293__bF_buf1), .Y(_12227_) );
AOI21X1 AOI21X1_2082 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe56_bF_buf3), .B(_12902_), .C(micro_hash_ucr_3_pipe57_bF_buf0), .Y(_12228_) );
AOI21X1 AOI21X1_2083 ( .gnd(gnd), .vdd(vdd), .A(_12228_), .B(_12227_), .C(micro_hash_ucr_3_pipe58_bF_buf2), .Y(_12229_) );
OAI21X1 OAI21X1_3445 ( .gnd(gnd), .vdd(vdd), .A(_9294__bF_buf3), .B(micro_hash_ucr_3_b_0_bF_buf0_), .C(_9290__bF_buf2), .Y(_12230_) );
OAI21X1 OAI21X1_3446 ( .gnd(gnd), .vdd(vdd), .A(_12229_), .B(_12230_), .C(_9292__bF_buf1), .Y(_12231_) );
AOI21X1 AOI21X1_2084 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe60_bF_buf4), .B(_12902_), .C(micro_hash_ucr_3_pipe61_bF_buf2), .Y(_12232_) );
AOI21X1 AOI21X1_2085 ( .gnd(gnd), .vdd(vdd), .A(_12232_), .B(_12231_), .C(micro_hash_ucr_3_pipe62_bF_buf0), .Y(_12233_) );
OAI21X1 OAI21X1_3447 ( .gnd(gnd), .vdd(vdd), .A(_9287__bF_buf0), .B(micro_hash_ucr_3_b_0_bF_buf3_), .C(_9289__bF_buf1), .Y(_12234_) );
OAI21X1 OAI21X1_3448 ( .gnd(gnd), .vdd(vdd), .A(_12233_), .B(_12234_), .C(_9288__bF_buf1), .Y(_12235_) );
AOI21X1 AOI21X1_2086 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe64_bF_buf4), .B(_12902_), .C(micro_hash_ucr_3_pipe65_bF_buf0), .Y(_12236_) );
AOI21X1 AOI21X1_2087 ( .gnd(gnd), .vdd(vdd), .A(_12236_), .B(_12235_), .C(micro_hash_ucr_3_pipe66_bF_buf0), .Y(_12237_) );
OAI21X1 OAI21X1_3449 ( .gnd(gnd), .vdd(vdd), .A(_9286__bF_buf0), .B(micro_hash_ucr_3_b_0_bF_buf2_), .C(_9285__bF_buf3), .Y(_12238_) );
OAI21X1 OAI21X1_3450 ( .gnd(gnd), .vdd(vdd), .A(_12237_), .B(_12238_), .C(_9282__bF_buf1), .Y(_12239_) );
OAI21X1 OAI21X1_3451 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_0_bF_buf1_), .B(_9282__bF_buf0), .C(_12239_), .Y(_12240_) );
NOR2X1 NOR2X1_1950 ( .gnd(gnd), .vdd(vdd), .A(_10381_), .B(_12240_), .Y(_8701__0_) );
OAI21X1 OAI21X1_3452 ( .gnd(gnd), .vdd(vdd), .A(_12906_), .B(_9372_), .C(_12180_), .Y(_12241_) );
AOI21X1 AOI21X1_2088 ( .gnd(gnd), .vdd(vdd), .A(_9366_), .B(_12241_), .C(_12182_), .Y(_12242_) );
OAI21X1 OAI21X1_3453 ( .gnd(gnd), .vdd(vdd), .A(_12185_), .B(micro_hash_ucr_3_b_1_bF_buf0_), .C(_9337_), .Y(_12243_) );
OAI21X1 OAI21X1_3454 ( .gnd(gnd), .vdd(vdd), .A(_12242_), .B(_12243_), .C(_9336__bF_buf2), .Y(_12244_) );
AOI21X1 AOI21X1_2089 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe16_bF_buf4), .B(_12908__bF_buf3), .C(micro_hash_ucr_3_pipe17_bF_buf3), .Y(_12245_) );
AOI21X1 AOI21X1_2090 ( .gnd(gnd), .vdd(vdd), .A(_12245_), .B(_12244_), .C(micro_hash_ucr_3_pipe18_bF_buf3), .Y(_12246_) );
OAI21X1 OAI21X1_3455 ( .gnd(gnd), .vdd(vdd), .A(_9334__bF_buf3), .B(micro_hash_ucr_3_b_1_bF_buf3_), .C(_9333__bF_buf2), .Y(_12247_) );
OAI21X1 OAI21X1_3456 ( .gnd(gnd), .vdd(vdd), .A(_12246_), .B(_12247_), .C(_9329__bF_buf2), .Y(_12248_) );
AOI21X1 AOI21X1_2091 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe20_bF_buf4), .B(_12908__bF_buf2), .C(micro_hash_ucr_3_pipe21_bF_buf2), .Y(_12249_) );
AOI21X1 AOI21X1_2092 ( .gnd(gnd), .vdd(vdd), .A(_12249_), .B(_12248_), .C(micro_hash_ucr_3_pipe22_bF_buf0), .Y(_12250_) );
OAI21X1 OAI21X1_3457 ( .gnd(gnd), .vdd(vdd), .A(_9330__bF_buf1), .B(micro_hash_ucr_3_b_1_bF_buf2_), .C(_9326__bF_buf3), .Y(_12251_) );
OAI21X1 OAI21X1_3458 ( .gnd(gnd), .vdd(vdd), .A(_12250_), .B(_12251_), .C(_9328__bF_buf3), .Y(_12252_) );
AOI21X1 AOI21X1_2093 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe24_bF_buf4), .B(_12908__bF_buf1), .C(micro_hash_ucr_3_pipe25_bF_buf3), .Y(_12253_) );
AOI21X1 AOI21X1_2094 ( .gnd(gnd), .vdd(vdd), .A(_12253_), .B(_12252_), .C(micro_hash_ucr_3_pipe26_bF_buf1), .Y(_12254_) );
OAI21X1 OAI21X1_3459 ( .gnd(gnd), .vdd(vdd), .A(_9323__bF_buf1), .B(micro_hash_ucr_3_b_1_bF_buf1_), .C(_9325__bF_buf3), .Y(_12255_) );
OAI21X1 OAI21X1_3460 ( .gnd(gnd), .vdd(vdd), .A(_12254_), .B(_12255_), .C(_9324__bF_buf0), .Y(_12256_) );
AOI21X1 AOI21X1_2095 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe28_bF_buf2), .B(_12908__bF_buf0), .C(micro_hash_ucr_3_pipe29_bF_buf2), .Y(_12257_) );
AOI21X1 AOI21X1_2096 ( .gnd(gnd), .vdd(vdd), .A(_12257_), .B(_12256_), .C(micro_hash_ucr_3_pipe30_bF_buf2), .Y(_12258_) );
OAI21X1 OAI21X1_3461 ( .gnd(gnd), .vdd(vdd), .A(_9322__bF_buf1), .B(micro_hash_ucr_3_b_1_bF_buf0_), .C(_9321__bF_buf0), .Y(_12259_) );
OAI21X1 OAI21X1_3462 ( .gnd(gnd), .vdd(vdd), .A(_12258_), .B(_12259_), .C(_9317__bF_buf4), .Y(_12260_) );
AOI21X1 AOI21X1_2097 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe32_bF_buf0), .B(_12908__bF_buf3), .C(micro_hash_ucr_3_pipe33_bF_buf1), .Y(_12261_) );
AOI21X1 AOI21X1_2098 ( .gnd(gnd), .vdd(vdd), .A(_12261_), .B(_12260_), .C(micro_hash_ucr_3_pipe34_bF_buf1), .Y(_12262_) );
OAI21X1 OAI21X1_3463 ( .gnd(gnd), .vdd(vdd), .A(_9318__bF_buf1), .B(micro_hash_ucr_3_b_1_bF_buf3_), .C(_9314_), .Y(_12263_) );
OAI21X1 OAI21X1_3464 ( .gnd(gnd), .vdd(vdd), .A(_12262_), .B(_12263_), .C(_9316__bF_buf2), .Y(_12264_) );
AOI21X1 AOI21X1_2099 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe36_bF_buf1), .B(_12908__bF_buf2), .C(micro_hash_ucr_3_pipe37_bF_buf1), .Y(_12265_) );
AOI21X1 AOI21X1_2100 ( .gnd(gnd), .vdd(vdd), .A(_12265_), .B(_12264_), .C(micro_hash_ucr_3_pipe38_bF_buf0), .Y(_12266_) );
OAI21X1 OAI21X1_3465 ( .gnd(gnd), .vdd(vdd), .A(_9311__bF_buf3), .B(micro_hash_ucr_3_b_1_bF_buf2_), .C(_9313_), .Y(_12267_) );
OAI21X1 OAI21X1_3466 ( .gnd(gnd), .vdd(vdd), .A(_12266_), .B(_12267_), .C(_9312__bF_buf2), .Y(_12268_) );
AOI21X1 AOI21X1_2101 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe40_bF_buf1), .B(_12908__bF_buf1), .C(micro_hash_ucr_3_pipe41_bF_buf1), .Y(_12269_) );
AOI21X1 AOI21X1_2102 ( .gnd(gnd), .vdd(vdd), .A(_12269_), .B(_12268_), .C(micro_hash_ucr_3_pipe42_bF_buf2), .Y(_12270_) );
OAI21X1 OAI21X1_3467 ( .gnd(gnd), .vdd(vdd), .A(_9310__bF_buf0), .B(micro_hash_ucr_3_b_1_bF_buf1_), .C(_9309__bF_buf1), .Y(_12271_) );
OAI21X1 OAI21X1_3468 ( .gnd(gnd), .vdd(vdd), .A(_12270_), .B(_12271_), .C(_9305__bF_buf3), .Y(_12272_) );
AOI21X1 AOI21X1_2103 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe44_bF_buf0), .B(_12908__bF_buf0), .C(micro_hash_ucr_3_pipe45_bF_buf0), .Y(_12273_) );
AOI21X1 AOI21X1_2104 ( .gnd(gnd), .vdd(vdd), .A(_12273_), .B(_12272_), .C(micro_hash_ucr_3_pipe46_bF_buf1), .Y(_12274_) );
OAI21X1 OAI21X1_3469 ( .gnd(gnd), .vdd(vdd), .A(_9306__bF_buf2), .B(micro_hash_ucr_3_b_1_bF_buf0_), .C(_9302_), .Y(_12275_) );
OAI21X1 OAI21X1_3470 ( .gnd(gnd), .vdd(vdd), .A(_12274_), .B(_12275_), .C(_9304__bF_buf1), .Y(_12276_) );
AOI21X1 AOI21X1_2105 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe48_bF_buf1), .B(_12908__bF_buf3), .C(micro_hash_ucr_3_pipe49_bF_buf0), .Y(_12277_) );
AOI21X1 AOI21X1_2106 ( .gnd(gnd), .vdd(vdd), .A(_12277_), .B(_12276_), .C(micro_hash_ucr_3_pipe50_bF_buf1), .Y(_12278_) );
OAI21X1 OAI21X1_3471 ( .gnd(gnd), .vdd(vdd), .A(_9299__bF_buf1), .B(micro_hash_ucr_3_b_1_bF_buf3_), .C(_9301__bF_buf0), .Y(_12279_) );
OAI21X1 OAI21X1_3472 ( .gnd(gnd), .vdd(vdd), .A(_12278_), .B(_12279_), .C(_9300__bF_buf2), .Y(_12280_) );
AOI21X1 AOI21X1_2107 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe52_bF_buf0), .B(_12908__bF_buf2), .C(micro_hash_ucr_3_pipe53), .Y(_12281_) );
AOI21X1 AOI21X1_2108 ( .gnd(gnd), .vdd(vdd), .A(_12281_), .B(_12280_), .C(micro_hash_ucr_3_pipe54_bF_buf0), .Y(_12282_) );
OAI21X1 OAI21X1_3473 ( .gnd(gnd), .vdd(vdd), .A(_9298__bF_buf3), .B(micro_hash_ucr_3_b_1_bF_buf2_), .C(_9297_), .Y(_12283_) );
OAI21X1 OAI21X1_3474 ( .gnd(gnd), .vdd(vdd), .A(_12282_), .B(_12283_), .C(_9293__bF_buf0), .Y(_12284_) );
AOI21X1 AOI21X1_2109 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe56_bF_buf2), .B(_12908__bF_buf1), .C(micro_hash_ucr_3_pipe57_bF_buf3), .Y(_12285_) );
AOI21X1 AOI21X1_2110 ( .gnd(gnd), .vdd(vdd), .A(_12285_), .B(_12284_), .C(micro_hash_ucr_3_pipe58_bF_buf1), .Y(_12286_) );
OAI21X1 OAI21X1_3475 ( .gnd(gnd), .vdd(vdd), .A(_9294__bF_buf2), .B(micro_hash_ucr_3_b_1_bF_buf1_), .C(_9290__bF_buf1), .Y(_12287_) );
OAI21X1 OAI21X1_3476 ( .gnd(gnd), .vdd(vdd), .A(_12286_), .B(_12287_), .C(_9292__bF_buf0), .Y(_12288_) );
AOI21X1 AOI21X1_2111 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe60_bF_buf3), .B(_12908__bF_buf0), .C(micro_hash_ucr_3_pipe61_bF_buf1), .Y(_12289_) );
AOI21X1 AOI21X1_2112 ( .gnd(gnd), .vdd(vdd), .A(_12289_), .B(_12288_), .C(micro_hash_ucr_3_pipe62_bF_buf3), .Y(_12290_) );
OAI21X1 OAI21X1_3477 ( .gnd(gnd), .vdd(vdd), .A(_9287__bF_buf4), .B(micro_hash_ucr_3_b_1_bF_buf0_), .C(_9289__bF_buf0), .Y(_12291_) );
OAI21X1 OAI21X1_3478 ( .gnd(gnd), .vdd(vdd), .A(_12290_), .B(_12291_), .C(_9288__bF_buf0), .Y(_12292_) );
AOI21X1 AOI21X1_2113 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe64_bF_buf3), .B(_12908__bF_buf3), .C(micro_hash_ucr_3_pipe65_bF_buf3), .Y(_12293_) );
AOI21X1 AOI21X1_2114 ( .gnd(gnd), .vdd(vdd), .A(_12293_), .B(_12292_), .C(micro_hash_ucr_3_pipe66_bF_buf4), .Y(_12294_) );
OAI21X1 OAI21X1_3479 ( .gnd(gnd), .vdd(vdd), .A(_9286__bF_buf3), .B(micro_hash_ucr_3_b_1_bF_buf3_), .C(_9285__bF_buf2), .Y(_12295_) );
OAI21X1 OAI21X1_3480 ( .gnd(gnd), .vdd(vdd), .A(_12294_), .B(_12295_), .C(_9282__bF_buf4), .Y(_12296_) );
OAI21X1 OAI21X1_3481 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_1_bF_buf2_), .B(_9282__bF_buf3), .C(_12296_), .Y(_12297_) );
NOR2X1 NOR2X1_1951 ( .gnd(gnd), .vdd(vdd), .A(_10381_), .B(_12297_), .Y(_8701__1_) );
OAI21X1 OAI21X1_3482 ( .gnd(gnd), .vdd(vdd), .A(_8779_), .B(_9372_), .C(_12180_), .Y(_12298_) );
AOI21X1 AOI21X1_2115 ( .gnd(gnd), .vdd(vdd), .A(_9366_), .B(_12298_), .C(_12182_), .Y(_12299_) );
OAI21X1 OAI21X1_3483 ( .gnd(gnd), .vdd(vdd), .A(_12185_), .B(micro_hash_ucr_3_b_2_bF_buf0_), .C(_9337_), .Y(_12300_) );
OAI21X1 OAI21X1_3484 ( .gnd(gnd), .vdd(vdd), .A(_12299_), .B(_12300_), .C(_9336__bF_buf1), .Y(_12301_) );
AOI21X1 AOI21X1_2116 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe16_bF_buf3), .B(_8789__bF_buf3), .C(micro_hash_ucr_3_pipe17_bF_buf2), .Y(_12302_) );
AOI21X1 AOI21X1_2117 ( .gnd(gnd), .vdd(vdd), .A(_12302_), .B(_12301_), .C(micro_hash_ucr_3_pipe18_bF_buf2), .Y(_12303_) );
OAI21X1 OAI21X1_3485 ( .gnd(gnd), .vdd(vdd), .A(_9334__bF_buf2), .B(micro_hash_ucr_3_b_2_bF_buf3_), .C(_9333__bF_buf1), .Y(_12304_) );
OAI21X1 OAI21X1_3486 ( .gnd(gnd), .vdd(vdd), .A(_12303_), .B(_12304_), .C(_9329__bF_buf1), .Y(_12305_) );
AOI21X1 AOI21X1_2118 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe20_bF_buf3), .B(_8789__bF_buf2), .C(micro_hash_ucr_3_pipe21_bF_buf1), .Y(_12306_) );
AOI21X1 AOI21X1_2119 ( .gnd(gnd), .vdd(vdd), .A(_12306_), .B(_12305_), .C(micro_hash_ucr_3_pipe22_bF_buf4), .Y(_12307_) );
OAI21X1 OAI21X1_3487 ( .gnd(gnd), .vdd(vdd), .A(_9330__bF_buf0), .B(micro_hash_ucr_3_b_2_bF_buf2_), .C(_9326__bF_buf2), .Y(_12308_) );
OAI21X1 OAI21X1_3488 ( .gnd(gnd), .vdd(vdd), .A(_12307_), .B(_12308_), .C(_9328__bF_buf2), .Y(_12309_) );
AOI21X1 AOI21X1_2120 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe24_bF_buf3), .B(_8789__bF_buf1), .C(micro_hash_ucr_3_pipe25_bF_buf2), .Y(_12310_) );
AOI21X1 AOI21X1_2121 ( .gnd(gnd), .vdd(vdd), .A(_12310_), .B(_12309_), .C(micro_hash_ucr_3_pipe26_bF_buf0), .Y(_12311_) );
OAI21X1 OAI21X1_3489 ( .gnd(gnd), .vdd(vdd), .A(_9323__bF_buf0), .B(micro_hash_ucr_3_b_2_bF_buf1_), .C(_9325__bF_buf2), .Y(_12312_) );
OAI21X1 OAI21X1_3490 ( .gnd(gnd), .vdd(vdd), .A(_12311_), .B(_12312_), .C(_9324__bF_buf4), .Y(_12313_) );
AOI21X1 AOI21X1_2122 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe28_bF_buf1), .B(_8789__bF_buf0), .C(micro_hash_ucr_3_pipe29_bF_buf1), .Y(_12314_) );
AOI21X1 AOI21X1_2123 ( .gnd(gnd), .vdd(vdd), .A(_12314_), .B(_12313_), .C(micro_hash_ucr_3_pipe30_bF_buf1), .Y(_12315_) );
OAI21X1 OAI21X1_3491 ( .gnd(gnd), .vdd(vdd), .A(_9322__bF_buf0), .B(micro_hash_ucr_3_b_2_bF_buf0_), .C(_9321__bF_buf3), .Y(_12316_) );
OAI21X1 OAI21X1_3492 ( .gnd(gnd), .vdd(vdd), .A(_12315_), .B(_12316_), .C(_9317__bF_buf3), .Y(_12317_) );
AOI21X1 AOI21X1_2124 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe32_bF_buf3), .B(_8789__bF_buf3), .C(micro_hash_ucr_3_pipe33_bF_buf0), .Y(_12318_) );
AOI21X1 AOI21X1_2125 ( .gnd(gnd), .vdd(vdd), .A(_12318_), .B(_12317_), .C(micro_hash_ucr_3_pipe34_bF_buf0), .Y(_12319_) );
OAI21X1 OAI21X1_3493 ( .gnd(gnd), .vdd(vdd), .A(_9318__bF_buf0), .B(micro_hash_ucr_3_b_2_bF_buf3_), .C(_9314_), .Y(_12320_) );
OAI21X1 OAI21X1_3494 ( .gnd(gnd), .vdd(vdd), .A(_12319_), .B(_12320_), .C(_9316__bF_buf1), .Y(_12321_) );
AOI21X1 AOI21X1_2126 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe36_bF_buf0), .B(_8789__bF_buf2), .C(micro_hash_ucr_3_pipe37_bF_buf0), .Y(_12322_) );
AOI21X1 AOI21X1_2127 ( .gnd(gnd), .vdd(vdd), .A(_12322_), .B(_12321_), .C(micro_hash_ucr_3_pipe38_bF_buf3), .Y(_12323_) );
OAI21X1 OAI21X1_3495 ( .gnd(gnd), .vdd(vdd), .A(_9311__bF_buf2), .B(micro_hash_ucr_3_b_2_bF_buf2_), .C(_9313_), .Y(_12324_) );
OAI21X1 OAI21X1_3496 ( .gnd(gnd), .vdd(vdd), .A(_12323_), .B(_12324_), .C(_9312__bF_buf1), .Y(_12325_) );
AOI21X1 AOI21X1_2128 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe40_bF_buf0), .B(_8789__bF_buf1), .C(micro_hash_ucr_3_pipe41_bF_buf0), .Y(_12326_) );
AOI21X1 AOI21X1_2129 ( .gnd(gnd), .vdd(vdd), .A(_12326_), .B(_12325_), .C(micro_hash_ucr_3_pipe42_bF_buf1), .Y(_12327_) );
OAI21X1 OAI21X1_3497 ( .gnd(gnd), .vdd(vdd), .A(_9310__bF_buf4), .B(micro_hash_ucr_3_b_2_bF_buf1_), .C(_9309__bF_buf0), .Y(_12328_) );
OAI21X1 OAI21X1_3498 ( .gnd(gnd), .vdd(vdd), .A(_12327_), .B(_12328_), .C(_9305__bF_buf2), .Y(_12329_) );
AOI21X1 AOI21X1_2130 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe44_bF_buf3), .B(_8789__bF_buf0), .C(micro_hash_ucr_3_pipe45_bF_buf3), .Y(_12330_) );
AOI21X1 AOI21X1_2131 ( .gnd(gnd), .vdd(vdd), .A(_12330_), .B(_12329_), .C(micro_hash_ucr_3_pipe46_bF_buf0), .Y(_12331_) );
OAI21X1 OAI21X1_3499 ( .gnd(gnd), .vdd(vdd), .A(_9306__bF_buf1), .B(micro_hash_ucr_3_b_2_bF_buf0_), .C(_9302_), .Y(_12332_) );
OAI21X1 OAI21X1_3500 ( .gnd(gnd), .vdd(vdd), .A(_12331_), .B(_12332_), .C(_9304__bF_buf0), .Y(_12333_) );
AOI21X1 AOI21X1_2132 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe48_bF_buf0), .B(_8789__bF_buf3), .C(micro_hash_ucr_3_pipe49_bF_buf3), .Y(_12334_) );
AOI21X1 AOI21X1_2133 ( .gnd(gnd), .vdd(vdd), .A(_12334_), .B(_12333_), .C(micro_hash_ucr_3_pipe50_bF_buf0), .Y(_12335_) );
OAI21X1 OAI21X1_3501 ( .gnd(gnd), .vdd(vdd), .A(_9299__bF_buf0), .B(micro_hash_ucr_3_b_2_bF_buf3_), .C(_9301__bF_buf3), .Y(_12336_) );
OAI21X1 OAI21X1_3502 ( .gnd(gnd), .vdd(vdd), .A(_12335_), .B(_12336_), .C(_9300__bF_buf1), .Y(_12337_) );
AOI21X1 AOI21X1_2134 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe52_bF_buf4), .B(_8789__bF_buf2), .C(micro_hash_ucr_3_pipe53), .Y(_12338_) );
AOI21X1 AOI21X1_2135 ( .gnd(gnd), .vdd(vdd), .A(_12338_), .B(_12337_), .C(micro_hash_ucr_3_pipe54_bF_buf3), .Y(_12339_) );
OAI21X1 OAI21X1_3503 ( .gnd(gnd), .vdd(vdd), .A(_9298__bF_buf2), .B(micro_hash_ucr_3_b_2_bF_buf2_), .C(_9297_), .Y(_12340_) );
OAI21X1 OAI21X1_3504 ( .gnd(gnd), .vdd(vdd), .A(_12339_), .B(_12340_), .C(_9293__bF_buf3), .Y(_12341_) );
AOI21X1 AOI21X1_2136 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe56_bF_buf1), .B(_8789__bF_buf1), .C(micro_hash_ucr_3_pipe57_bF_buf2), .Y(_12342_) );
AOI21X1 AOI21X1_2137 ( .gnd(gnd), .vdd(vdd), .A(_12342_), .B(_12341_), .C(micro_hash_ucr_3_pipe58_bF_buf0), .Y(_12343_) );
OAI21X1 OAI21X1_3505 ( .gnd(gnd), .vdd(vdd), .A(_9294__bF_buf1), .B(micro_hash_ucr_3_b_2_bF_buf1_), .C(_9290__bF_buf0), .Y(_12344_) );
OAI21X1 OAI21X1_3506 ( .gnd(gnd), .vdd(vdd), .A(_12343_), .B(_12344_), .C(_9292__bF_buf3), .Y(_12345_) );
AOI21X1 AOI21X1_2138 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe60_bF_buf2), .B(_8789__bF_buf0), .C(micro_hash_ucr_3_pipe61_bF_buf0), .Y(_12346_) );
AOI21X1 AOI21X1_2139 ( .gnd(gnd), .vdd(vdd), .A(_12346_), .B(_12345_), .C(micro_hash_ucr_3_pipe62_bF_buf2), .Y(_12347_) );
OAI21X1 OAI21X1_3507 ( .gnd(gnd), .vdd(vdd), .A(_9287__bF_buf3), .B(micro_hash_ucr_3_b_2_bF_buf0_), .C(_9289__bF_buf3), .Y(_12348_) );
OAI21X1 OAI21X1_3508 ( .gnd(gnd), .vdd(vdd), .A(_12347_), .B(_12348_), .C(_9288__bF_buf3), .Y(_12349_) );
AOI21X1 AOI21X1_2140 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe64_bF_buf2), .B(_8789__bF_buf3), .C(micro_hash_ucr_3_pipe65_bF_buf2), .Y(_12350_) );
AOI21X1 AOI21X1_2141 ( .gnd(gnd), .vdd(vdd), .A(_12350_), .B(_12349_), .C(micro_hash_ucr_3_pipe66_bF_buf3), .Y(_12351_) );
OAI21X1 OAI21X1_3509 ( .gnd(gnd), .vdd(vdd), .A(_9286__bF_buf2), .B(micro_hash_ucr_3_b_2_bF_buf3_), .C(_9285__bF_buf1), .Y(_12352_) );
OAI21X1 OAI21X1_3510 ( .gnd(gnd), .vdd(vdd), .A(_12351_), .B(_12352_), .C(_9282__bF_buf2), .Y(_12353_) );
OAI21X1 OAI21X1_3511 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_2_bF_buf2_), .B(_9282__bF_buf1), .C(_12353_), .Y(_12354_) );
NOR2X1 NOR2X1_1952 ( .gnd(gnd), .vdd(vdd), .A(_10381_), .B(_12354_), .Y(_8701__2_) );
OAI21X1 OAI21X1_3512 ( .gnd(gnd), .vdd(vdd), .A(_8793_), .B(_9372_), .C(_12180_), .Y(_12355_) );
AOI21X1 AOI21X1_2142 ( .gnd(gnd), .vdd(vdd), .A(_9366_), .B(_12355_), .C(_12182_), .Y(_12356_) );
OAI21X1 OAI21X1_3513 ( .gnd(gnd), .vdd(vdd), .A(_12185_), .B(micro_hash_ucr_3_b_3_bF_buf3_), .C(_9337_), .Y(_12357_) );
OAI21X1 OAI21X1_3514 ( .gnd(gnd), .vdd(vdd), .A(_12356_), .B(_12357_), .C(_9336__bF_buf0), .Y(_12358_) );
AOI21X1 AOI21X1_2143 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe16_bF_buf2), .B(_8794_), .C(micro_hash_ucr_3_pipe17_bF_buf1), .Y(_12359_) );
AOI21X1 AOI21X1_2144 ( .gnd(gnd), .vdd(vdd), .A(_12359_), .B(_12358_), .C(micro_hash_ucr_3_pipe18_bF_buf1), .Y(_12360_) );
OAI21X1 OAI21X1_3515 ( .gnd(gnd), .vdd(vdd), .A(_9334__bF_buf1), .B(micro_hash_ucr_3_b_3_bF_buf2_), .C(_9333__bF_buf0), .Y(_12361_) );
OAI21X1 OAI21X1_3516 ( .gnd(gnd), .vdd(vdd), .A(_12360_), .B(_12361_), .C(_9329__bF_buf0), .Y(_12362_) );
AOI21X1 AOI21X1_2145 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe20_bF_buf2), .B(_8794_), .C(micro_hash_ucr_3_pipe21_bF_buf0), .Y(_12363_) );
AOI21X1 AOI21X1_2146 ( .gnd(gnd), .vdd(vdd), .A(_12363_), .B(_12362_), .C(micro_hash_ucr_3_pipe22_bF_buf3), .Y(_12364_) );
OAI21X1 OAI21X1_3517 ( .gnd(gnd), .vdd(vdd), .A(_9330__bF_buf4), .B(micro_hash_ucr_3_b_3_bF_buf1_), .C(_9326__bF_buf1), .Y(_12365_) );
OAI21X1 OAI21X1_3518 ( .gnd(gnd), .vdd(vdd), .A(_12364_), .B(_12365_), .C(_9328__bF_buf1), .Y(_12366_) );
AOI21X1 AOI21X1_2147 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe24_bF_buf2), .B(_8794_), .C(micro_hash_ucr_3_pipe25_bF_buf1), .Y(_12367_) );
AOI21X1 AOI21X1_2148 ( .gnd(gnd), .vdd(vdd), .A(_12367_), .B(_12366_), .C(micro_hash_ucr_3_pipe26_bF_buf4), .Y(_12368_) );
OAI21X1 OAI21X1_3519 ( .gnd(gnd), .vdd(vdd), .A(_9323__bF_buf3), .B(micro_hash_ucr_3_b_3_bF_buf0_), .C(_9325__bF_buf1), .Y(_12369_) );
OAI21X1 OAI21X1_3520 ( .gnd(gnd), .vdd(vdd), .A(_12368_), .B(_12369_), .C(_9324__bF_buf3), .Y(_12370_) );
AOI21X1 AOI21X1_2149 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe28_bF_buf0), .B(_8794_), .C(micro_hash_ucr_3_pipe29_bF_buf0), .Y(_12371_) );
AOI21X1 AOI21X1_2150 ( .gnd(gnd), .vdd(vdd), .A(_12371_), .B(_12370_), .C(micro_hash_ucr_3_pipe30_bF_buf0), .Y(_12372_) );
OAI21X1 OAI21X1_3521 ( .gnd(gnd), .vdd(vdd), .A(_9322__bF_buf3), .B(micro_hash_ucr_3_b_3_bF_buf3_), .C(_9321__bF_buf2), .Y(_12373_) );
OAI21X1 OAI21X1_3522 ( .gnd(gnd), .vdd(vdd), .A(_12372_), .B(_12373_), .C(_9317__bF_buf2), .Y(_12374_) );
AOI21X1 AOI21X1_2151 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe32_bF_buf2), .B(_8794_), .C(micro_hash_ucr_3_pipe33_bF_buf3), .Y(_12375_) );
AOI21X1 AOI21X1_2152 ( .gnd(gnd), .vdd(vdd), .A(_12375_), .B(_12374_), .C(micro_hash_ucr_3_pipe34_bF_buf4), .Y(_12376_) );
OAI21X1 OAI21X1_3523 ( .gnd(gnd), .vdd(vdd), .A(_9318__bF_buf4), .B(micro_hash_ucr_3_b_3_bF_buf2_), .C(_9314_), .Y(_12377_) );
OAI21X1 OAI21X1_3524 ( .gnd(gnd), .vdd(vdd), .A(_12376_), .B(_12377_), .C(_9316__bF_buf0), .Y(_12378_) );
AOI21X1 AOI21X1_2153 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe36_bF_buf4), .B(_8794_), .C(micro_hash_ucr_3_pipe37_bF_buf3), .Y(_12379_) );
AOI21X1 AOI21X1_2154 ( .gnd(gnd), .vdd(vdd), .A(_12379_), .B(_12378_), .C(micro_hash_ucr_3_pipe38_bF_buf2), .Y(_12380_) );
OAI21X1 OAI21X1_3525 ( .gnd(gnd), .vdd(vdd), .A(_9311__bF_buf1), .B(micro_hash_ucr_3_b_3_bF_buf1_), .C(_9313_), .Y(_12381_) );
OAI21X1 OAI21X1_3526 ( .gnd(gnd), .vdd(vdd), .A(_12380_), .B(_12381_), .C(_9312__bF_buf0), .Y(_12382_) );
AOI21X1 AOI21X1_2155 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe40_bF_buf4), .B(_8794_), .C(micro_hash_ucr_3_pipe41_bF_buf3), .Y(_12383_) );
AOI21X1 AOI21X1_2156 ( .gnd(gnd), .vdd(vdd), .A(_12383_), .B(_12382_), .C(micro_hash_ucr_3_pipe42_bF_buf0), .Y(_12384_) );
OAI21X1 OAI21X1_3527 ( .gnd(gnd), .vdd(vdd), .A(_9310__bF_buf3), .B(micro_hash_ucr_3_b_3_bF_buf0_), .C(_9309__bF_buf3), .Y(_12385_) );
OAI21X1 OAI21X1_3528 ( .gnd(gnd), .vdd(vdd), .A(_12384_), .B(_12385_), .C(_9305__bF_buf1), .Y(_12386_) );
AOI21X1 AOI21X1_2157 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe44_bF_buf2), .B(_8794_), .C(micro_hash_ucr_3_pipe45_bF_buf2), .Y(_12387_) );
AOI21X1 AOI21X1_2158 ( .gnd(gnd), .vdd(vdd), .A(_12387_), .B(_12386_), .C(micro_hash_ucr_3_pipe46_bF_buf4), .Y(_12388_) );
OAI21X1 OAI21X1_3529 ( .gnd(gnd), .vdd(vdd), .A(_9306__bF_buf0), .B(micro_hash_ucr_3_b_3_bF_buf3_), .C(_9302_), .Y(_12389_) );
OAI21X1 OAI21X1_3530 ( .gnd(gnd), .vdd(vdd), .A(_12388_), .B(_12389_), .C(_9304__bF_buf3), .Y(_12390_) );
AOI21X1 AOI21X1_2159 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe48_bF_buf4), .B(_8794_), .C(micro_hash_ucr_3_pipe49_bF_buf2), .Y(_12391_) );
AOI21X1 AOI21X1_2160 ( .gnd(gnd), .vdd(vdd), .A(_12391_), .B(_12390_), .C(micro_hash_ucr_3_pipe50_bF_buf4), .Y(_12392_) );
OAI21X1 OAI21X1_3531 ( .gnd(gnd), .vdd(vdd), .A(_9299__bF_buf3), .B(micro_hash_ucr_3_b_3_bF_buf2_), .C(_9301__bF_buf2), .Y(_12393_) );
OAI21X1 OAI21X1_3532 ( .gnd(gnd), .vdd(vdd), .A(_12392_), .B(_12393_), .C(_9300__bF_buf0), .Y(_12394_) );
AOI21X1 AOI21X1_2161 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe52_bF_buf3), .B(_8794_), .C(micro_hash_ucr_3_pipe53), .Y(_12395_) );
AOI21X1 AOI21X1_2162 ( .gnd(gnd), .vdd(vdd), .A(_12395_), .B(_12394_), .C(micro_hash_ucr_3_pipe54_bF_buf2), .Y(_12396_) );
OAI21X1 OAI21X1_3533 ( .gnd(gnd), .vdd(vdd), .A(_9298__bF_buf1), .B(micro_hash_ucr_3_b_3_bF_buf1_), .C(_9297_), .Y(_12397_) );
OAI21X1 OAI21X1_3534 ( .gnd(gnd), .vdd(vdd), .A(_12396_), .B(_12397_), .C(_9293__bF_buf2), .Y(_12398_) );
AOI21X1 AOI21X1_2163 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe56_bF_buf0), .B(_8794_), .C(micro_hash_ucr_3_pipe57_bF_buf1), .Y(_12399_) );
AOI21X1 AOI21X1_2164 ( .gnd(gnd), .vdd(vdd), .A(_12399_), .B(_12398_), .C(micro_hash_ucr_3_pipe58_bF_buf3), .Y(_12400_) );
OAI21X1 OAI21X1_3535 ( .gnd(gnd), .vdd(vdd), .A(_9294__bF_buf0), .B(micro_hash_ucr_3_b_3_bF_buf0_), .C(_9290__bF_buf3), .Y(_12401_) );
OAI21X1 OAI21X1_3536 ( .gnd(gnd), .vdd(vdd), .A(_12400_), .B(_12401_), .C(_9292__bF_buf2), .Y(_12402_) );
AOI21X1 AOI21X1_2165 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe60_bF_buf1), .B(_8794_), .C(micro_hash_ucr_3_pipe61_bF_buf3), .Y(_12403_) );
AOI21X1 AOI21X1_2166 ( .gnd(gnd), .vdd(vdd), .A(_12403_), .B(_12402_), .C(micro_hash_ucr_3_pipe62_bF_buf1), .Y(_12404_) );
OAI21X1 OAI21X1_3537 ( .gnd(gnd), .vdd(vdd), .A(_9287__bF_buf2), .B(micro_hash_ucr_3_b_3_bF_buf3_), .C(_9289__bF_buf2), .Y(_12405_) );
OAI21X1 OAI21X1_3538 ( .gnd(gnd), .vdd(vdd), .A(_12404_), .B(_12405_), .C(_9288__bF_buf2), .Y(_12406_) );
AOI21X1 AOI21X1_2167 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe64_bF_buf1), .B(_8794_), .C(micro_hash_ucr_3_pipe65_bF_buf1), .Y(_12407_) );
AOI21X1 AOI21X1_2168 ( .gnd(gnd), .vdd(vdd), .A(_12407_), .B(_12406_), .C(micro_hash_ucr_3_pipe66_bF_buf2), .Y(_12408_) );
OAI21X1 OAI21X1_3539 ( .gnd(gnd), .vdd(vdd), .A(_9286__bF_buf1), .B(micro_hash_ucr_3_b_3_bF_buf2_), .C(_9285__bF_buf0), .Y(_12409_) );
OAI21X1 OAI21X1_3540 ( .gnd(gnd), .vdd(vdd), .A(_12408_), .B(_12409_), .C(_9282__bF_buf0), .Y(_12410_) );
OAI21X1 OAI21X1_3541 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_3_bF_buf1_), .B(_9282__bF_buf4), .C(_12410_), .Y(_12411_) );
NOR2X1 NOR2X1_1953 ( .gnd(gnd), .vdd(vdd), .A(_10381_), .B(_12411_), .Y(_8701__3_) );
NAND2X1 NAND2X1_1581 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_4_bF_buf4_), .B(micro_hash_ucr_3_pipe66_bF_buf1), .Y(_12412_) );
NAND2X1 NAND2X1_1582 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_4_bF_buf3_), .B(micro_hash_ucr_3_pipe64_bF_buf0), .Y(_12413_) );
NAND2X1 NAND2X1_1583 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe63), .B(_12848__bF_buf0), .Y(_12414_) );
NAND2X1 NAND2X1_1584 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_4_bF_buf2_), .B(micro_hash_ucr_3_pipe62_bF_buf0), .Y(_12415_) );
NAND2X1 NAND2X1_1585 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe61_bF_buf2), .B(_12848__bF_buf3), .Y(_12416_) );
NAND2X1 NAND2X1_1586 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_4_bF_buf1_), .B(micro_hash_ucr_3_pipe60_bF_buf0), .Y(_12417_) );
NAND2X1 NAND2X1_1587 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe59), .B(_12848__bF_buf2), .Y(_12418_) );
NAND2X1 NAND2X1_1588 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_4_bF_buf0_), .B(micro_hash_ucr_3_pipe58_bF_buf2), .Y(_12419_) );
NAND2X1 NAND2X1_1589 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe57_bF_buf0), .B(_12848__bF_buf1), .Y(_12420_) );
NAND2X1 NAND2X1_1590 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_0_), .B(micro_hash_ucr_3_pipe53), .Y(_12421_) );
NAND2X1 NAND2X1_1591 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe49_bF_buf1), .B(_12848__bF_buf0), .Y(_12422_) );
NAND2X1 NAND2X1_1592 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_4_bF_buf4_), .B(micro_hash_ucr_3_pipe42_bF_buf3), .Y(_12423_) );
NAND2X1 NAND2X1_1593 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe41_bF_buf2), .B(_12848__bF_buf3), .Y(_12424_) );
NAND2X1 NAND2X1_1594 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_4_bF_buf3_), .B(micro_hash_ucr_3_pipe40_bF_buf3), .Y(_12425_) );
NAND2X1 NAND2X1_1595 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe39_bF_buf1), .B(_12848__bF_buf2), .Y(_12426_) );
NAND2X1 NAND2X1_1596 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_4_bF_buf2_), .B(micro_hash_ucr_3_pipe38_bF_buf1), .Y(_12427_) );
NAND2X1 NAND2X1_1597 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe37_bF_buf2), .B(_12848__bF_buf1), .Y(_12428_) );
NAND2X1 NAND2X1_1598 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_4_bF_buf1_), .B(micro_hash_ucr_3_pipe36_bF_buf3), .Y(_12429_) );
NAND2X1 NAND2X1_1599 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe35_bF_buf3), .B(_12848__bF_buf0), .Y(_12430_) );
NAND2X1 NAND2X1_1600 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_4_bF_buf0_), .B(micro_hash_ucr_3_pipe34_bF_buf3), .Y(_12431_) );
NAND2X1 NAND2X1_1601 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe33_bF_buf2), .B(_12848__bF_buf3), .Y(_12432_) );
NAND2X1 NAND2X1_1602 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_4_bF_buf4_), .B(micro_hash_ucr_3_pipe32_bF_buf1), .Y(_12433_) );
NOR2X1 NOR2X1_1954 ( .gnd(gnd), .vdd(vdd), .A(_12848__bF_buf2), .B(_9321__bF_buf1), .Y(_12434_) );
NAND2X1 NAND2X1_1603 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_4_bF_buf3_), .B(micro_hash_ucr_3_pipe30_bF_buf4), .Y(_12435_) );
NOR2X1 NOR2X1_1955 ( .gnd(gnd), .vdd(vdd), .A(_12848__bF_buf1), .B(_9320_), .Y(_12436_) );
NAND2X1 NAND2X1_1604 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_0_), .B(micro_hash_ucr_3_pipe25_bF_buf0), .Y(_12437_) );
NAND2X1 NAND2X1_1605 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe21_bF_buf3), .B(_12848__bF_buf0), .Y(_12438_) );
NAND2X1 NAND2X1_1606 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_4_bF_buf2_), .B(micro_hash_ucr_3_pipe18_bF_buf0), .Y(_12439_) );
NOR2X1 NOR2X1_1956 ( .gnd(gnd), .vdd(vdd), .A(H_3_12_), .B(micro_hash_ucr_3_pipe14_bF_buf1), .Y(_12440_) );
NOR2X1 NOR2X1_1957 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe15_bF_buf1), .B(micro_hash_ucr_3_pipe11), .Y(_12441_) );
NAND3X1 NAND3X1_601 ( .gnd(gnd), .vdd(vdd), .A(_9495_), .B(_12440_), .C(_12441_), .Y(_12442_) );
NAND2X1 NAND2X1_1607 ( .gnd(gnd), .vdd(vdd), .A(_9829_), .B(_10155_), .Y(_12443_) );
OAI22X1 OAI22X1_145 ( .gnd(gnd), .vdd(vdd), .A(_12442_), .B(_12443_), .C(_9600_), .D(micro_hash_ucr_3_c_0_), .Y(_12444_) );
NAND2X1 NAND2X1_1608 ( .gnd(gnd), .vdd(vdd), .A(_9336__bF_buf3), .B(_12444_), .Y(_12445_) );
NOR2X1 NOR2X1_1958 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_4_bF_buf1_), .B(_9627_), .Y(_12446_) );
NOR2X1 NOR2X1_1959 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe17_bF_buf0), .B(_12446_), .Y(_12447_) );
AOI22X1 AOI22X1_87 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_0_), .B(micro_hash_ucr_3_pipe17_bF_buf3), .C(_12447_), .D(_12445_), .Y(_12448_) );
OAI21X1 OAI21X1_3542 ( .gnd(gnd), .vdd(vdd), .A(_12448_), .B(micro_hash_ucr_3_pipe18_bF_buf4), .C(_12439_), .Y(_12449_) );
NAND2X1 NAND2X1_1609 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe19), .B(_12848__bF_buf3), .Y(_12450_) );
OAI21X1 OAI21X1_3543 ( .gnd(gnd), .vdd(vdd), .A(_12449_), .B(micro_hash_ucr_3_pipe19), .C(_12450_), .Y(_12451_) );
AOI21X1 AOI21X1_2169 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_4_bF_buf0_), .B(micro_hash_ucr_3_pipe20_bF_buf1), .C(micro_hash_ucr_3_pipe21_bF_buf2), .Y(_12452_) );
OAI21X1 OAI21X1_3544 ( .gnd(gnd), .vdd(vdd), .A(_12451_), .B(micro_hash_ucr_3_pipe20_bF_buf0), .C(_12452_), .Y(_12453_) );
AOI21X1 AOI21X1_2170 ( .gnd(gnd), .vdd(vdd), .A(_12438_), .B(_12453_), .C(micro_hash_ucr_3_pipe22_bF_buf2), .Y(_12454_) );
OAI21X1 OAI21X1_3545 ( .gnd(gnd), .vdd(vdd), .A(_9330__bF_buf3), .B(micro_hash_ucr_3_b_4_bF_buf4_), .C(_9326__bF_buf0), .Y(_12455_) );
AOI21X1 AOI21X1_2171 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_0_), .B(micro_hash_ucr_3_pipe23), .C(micro_hash_ucr_3_pipe24_bF_buf1), .Y(_12456_) );
OAI21X1 OAI21X1_3546 ( .gnd(gnd), .vdd(vdd), .A(_12454_), .B(_12455_), .C(_12456_), .Y(_12457_) );
NAND2X1 NAND2X1_1610 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe24_bF_buf0), .B(_10333_), .Y(_12458_) );
NAND3X1 NAND3X1_602 ( .gnd(gnd), .vdd(vdd), .A(_9327_), .B(_12458_), .C(_12457_), .Y(_12459_) );
AOI21X1 AOI21X1_2172 ( .gnd(gnd), .vdd(vdd), .A(_12437_), .B(_12459_), .C(micro_hash_ucr_3_pipe26_bF_buf3), .Y(_12460_) );
OAI21X1 OAI21X1_3547 ( .gnd(gnd), .vdd(vdd), .A(_10333_), .B(_9323__bF_buf2), .C(_9325__bF_buf0), .Y(_12461_) );
AOI21X1 AOI21X1_2173 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe27), .B(_12848__bF_buf2), .C(micro_hash_ucr_3_pipe28_bF_buf4), .Y(_12462_) );
OAI21X1 OAI21X1_3548 ( .gnd(gnd), .vdd(vdd), .A(_12460_), .B(_12461_), .C(_12462_), .Y(_12463_) );
NAND2X1 NAND2X1_1611 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_4_bF_buf3_), .B(micro_hash_ucr_3_pipe28_bF_buf3), .Y(_12464_) );
AOI21X1 AOI21X1_2174 ( .gnd(gnd), .vdd(vdd), .A(_12464_), .B(_12463_), .C(micro_hash_ucr_3_pipe29_bF_buf3), .Y(_12465_) );
OAI21X1 OAI21X1_3549 ( .gnd(gnd), .vdd(vdd), .A(_12465_), .B(_12436_), .C(_9322__bF_buf2), .Y(_12466_) );
AOI21X1 AOI21X1_2175 ( .gnd(gnd), .vdd(vdd), .A(_12435_), .B(_12466_), .C(micro_hash_ucr_3_pipe31), .Y(_12467_) );
OAI21X1 OAI21X1_3550 ( .gnd(gnd), .vdd(vdd), .A(_12467_), .B(_12434_), .C(_9317__bF_buf1), .Y(_12468_) );
NAND3X1 NAND3X1_603 ( .gnd(gnd), .vdd(vdd), .A(_9319_), .B(_12433_), .C(_12468_), .Y(_12469_) );
NAND3X1 NAND3X1_604 ( .gnd(gnd), .vdd(vdd), .A(_9318__bF_buf3), .B(_12432_), .C(_12469_), .Y(_12470_) );
NAND3X1 NAND3X1_605 ( .gnd(gnd), .vdd(vdd), .A(_9314_), .B(_12431_), .C(_12470_), .Y(_12471_) );
NAND3X1 NAND3X1_606 ( .gnd(gnd), .vdd(vdd), .A(_9316__bF_buf3), .B(_12430_), .C(_12471_), .Y(_12472_) );
NAND3X1 NAND3X1_607 ( .gnd(gnd), .vdd(vdd), .A(_9315_), .B(_12429_), .C(_12472_), .Y(_12473_) );
NAND3X1 NAND3X1_608 ( .gnd(gnd), .vdd(vdd), .A(_9311__bF_buf0), .B(_12428_), .C(_12473_), .Y(_12474_) );
NAND3X1 NAND3X1_609 ( .gnd(gnd), .vdd(vdd), .A(_9313_), .B(_12427_), .C(_12474_), .Y(_12475_) );
NAND3X1 NAND3X1_610 ( .gnd(gnd), .vdd(vdd), .A(_9312__bF_buf3), .B(_12426_), .C(_12475_), .Y(_12476_) );
NAND3X1 NAND3X1_611 ( .gnd(gnd), .vdd(vdd), .A(_9308_), .B(_12425_), .C(_12476_), .Y(_12477_) );
NAND3X1 NAND3X1_612 ( .gnd(gnd), .vdd(vdd), .A(_9310__bF_buf2), .B(_12424_), .C(_12477_), .Y(_12478_) );
AOI21X1 AOI21X1_2176 ( .gnd(gnd), .vdd(vdd), .A(_12423_), .B(_12478_), .C(micro_hash_ucr_3_pipe43), .Y(_12479_) );
OAI21X1 OAI21X1_3551 ( .gnd(gnd), .vdd(vdd), .A(_12848__bF_buf1), .B(_9309__bF_buf2), .C(_9305__bF_buf0), .Y(_12480_) );
AOI21X1 AOI21X1_2177 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe44_bF_buf1), .B(_10333_), .C(micro_hash_ucr_3_pipe45_bF_buf1), .Y(_12481_) );
OAI21X1 OAI21X1_3552 ( .gnd(gnd), .vdd(vdd), .A(_12479_), .B(_12480_), .C(_12481_), .Y(_12482_) );
AOI21X1 AOI21X1_2178 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_0_), .B(micro_hash_ucr_3_pipe45_bF_buf0), .C(micro_hash_ucr_3_pipe46_bF_buf3), .Y(_12483_) );
AOI22X1 AOI22X1_88 ( .gnd(gnd), .vdd(vdd), .A(_10333_), .B(micro_hash_ucr_3_pipe46_bF_buf2), .C(_12482_), .D(_12483_), .Y(_12484_) );
NAND2X1 NAND2X1_1612 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe47), .B(_12848__bF_buf0), .Y(_12485_) );
OAI21X1 OAI21X1_3553 ( .gnd(gnd), .vdd(vdd), .A(_12484_), .B(micro_hash_ucr_3_pipe47), .C(_12485_), .Y(_12486_) );
AOI21X1 AOI21X1_2179 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_4_bF_buf2_), .B(micro_hash_ucr_3_pipe48_bF_buf3), .C(micro_hash_ucr_3_pipe49_bF_buf0), .Y(_12487_) );
OAI21X1 OAI21X1_3554 ( .gnd(gnd), .vdd(vdd), .A(_12486_), .B(micro_hash_ucr_3_pipe48_bF_buf2), .C(_12487_), .Y(_12488_) );
AOI21X1 AOI21X1_2180 ( .gnd(gnd), .vdd(vdd), .A(_12422_), .B(_12488_), .C(micro_hash_ucr_3_pipe50_bF_buf3), .Y(_12489_) );
OAI21X1 OAI21X1_3555 ( .gnd(gnd), .vdd(vdd), .A(_9299__bF_buf2), .B(micro_hash_ucr_3_b_4_bF_buf1_), .C(_9301__bF_buf1), .Y(_12490_) );
AOI21X1 AOI21X1_2181 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_0_), .B(micro_hash_ucr_3_pipe51), .C(micro_hash_ucr_3_pipe52_bF_buf2), .Y(_12491_) );
OAI21X1 OAI21X1_3556 ( .gnd(gnd), .vdd(vdd), .A(_12489_), .B(_12490_), .C(_12491_), .Y(_12492_) );
NAND2X1 NAND2X1_1613 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe52_bF_buf1), .B(_10333_), .Y(_12493_) );
NAND3X1 NAND3X1_613 ( .gnd(gnd), .vdd(vdd), .A(_9296_), .B(_12493_), .C(_12492_), .Y(_12494_) );
AOI21X1 AOI21X1_2182 ( .gnd(gnd), .vdd(vdd), .A(_12421_), .B(_12494_), .C(micro_hash_ucr_3_pipe54_bF_buf1), .Y(_12495_) );
OAI21X1 OAI21X1_3557 ( .gnd(gnd), .vdd(vdd), .A(_10333_), .B(_9298__bF_buf0), .C(_9297_), .Y(_12496_) );
AOI21X1 AOI21X1_2183 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe55), .B(_12848__bF_buf3), .C(micro_hash_ucr_3_pipe56_bF_buf4), .Y(_12497_) );
OAI21X1 OAI21X1_3558 ( .gnd(gnd), .vdd(vdd), .A(_12495_), .B(_12496_), .C(_12497_), .Y(_12498_) );
NAND2X1 NAND2X1_1614 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_4_bF_buf0_), .B(micro_hash_ucr_3_pipe56_bF_buf3), .Y(_12499_) );
NAND3X1 NAND3X1_614 ( .gnd(gnd), .vdd(vdd), .A(_9295_), .B(_12499_), .C(_12498_), .Y(_12500_) );
NAND3X1 NAND3X1_615 ( .gnd(gnd), .vdd(vdd), .A(_9294__bF_buf4), .B(_12420_), .C(_12500_), .Y(_12501_) );
NAND3X1 NAND3X1_616 ( .gnd(gnd), .vdd(vdd), .A(_9290__bF_buf2), .B(_12419_), .C(_12501_), .Y(_12502_) );
NAND3X1 NAND3X1_617 ( .gnd(gnd), .vdd(vdd), .A(_9292__bF_buf1), .B(_12418_), .C(_12502_), .Y(_12503_) );
NAND3X1 NAND3X1_618 ( .gnd(gnd), .vdd(vdd), .A(_9291_), .B(_12417_), .C(_12503_), .Y(_12504_) );
NAND3X1 NAND3X1_619 ( .gnd(gnd), .vdd(vdd), .A(_9287__bF_buf1), .B(_12416_), .C(_12504_), .Y(_12505_) );
NAND3X1 NAND3X1_620 ( .gnd(gnd), .vdd(vdd), .A(_9289__bF_buf1), .B(_12415_), .C(_12505_), .Y(_12506_) );
NAND3X1 NAND3X1_621 ( .gnd(gnd), .vdd(vdd), .A(_9288__bF_buf1), .B(_12414_), .C(_12506_), .Y(_12507_) );
NAND3X1 NAND3X1_622 ( .gnd(gnd), .vdd(vdd), .A(_9284_), .B(_12413_), .C(_12507_), .Y(_12508_) );
OAI21X1 OAI21X1_3559 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_0_), .B(_9284_), .C(_12508_), .Y(_12509_) );
OAI21X1 OAI21X1_3560 ( .gnd(gnd), .vdd(vdd), .A(_12509_), .B(micro_hash_ucr_3_pipe66_bF_buf0), .C(_12412_), .Y(_12510_) );
OAI21X1 OAI21X1_3561 ( .gnd(gnd), .vdd(vdd), .A(_12848__bF_buf2), .B(_9285__bF_buf3), .C(_9282__bF_buf3), .Y(_12511_) );
AOI21X1 AOI21X1_2184 ( .gnd(gnd), .vdd(vdd), .A(_9285__bF_buf2), .B(_12510_), .C(_12511_), .Y(_12512_) );
OAI21X1 OAI21X1_3562 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_4_bF_buf4_), .B(_9282__bF_buf2), .C(_10380_), .Y(_12513_) );
OAI22X1 OAI22X1_146 ( .gnd(gnd), .vdd(vdd), .A(_12848__bF_buf1), .B(_11524_), .C(_12512_), .D(_12513_), .Y(_8701__4_) );
NAND2X1 NAND2X1_1615 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe66_bF_buf4), .B(_8814__bF_buf0), .Y(_12514_) );
NAND2X1 NAND2X1_1616 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_1_bF_buf3_), .B(micro_hash_ucr_3_pipe65_bF_buf0), .Y(_12515_) );
NAND2X1 NAND2X1_1617 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe64_bF_buf4), .B(_8814__bF_buf3), .Y(_12516_) );
NAND2X1 NAND2X1_1618 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_1_bF_buf2_), .B(micro_hash_ucr_3_pipe63), .Y(_12517_) );
NAND2X1 NAND2X1_1619 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe62_bF_buf3), .B(_8814__bF_buf2), .Y(_12518_) );
NAND2X1 NAND2X1_1620 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_1_bF_buf1_), .B(micro_hash_ucr_3_pipe61_bF_buf1), .Y(_12519_) );
NAND2X1 NAND2X1_1621 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe60_bF_buf4), .B(_8814__bF_buf1), .Y(_12520_) );
NAND2X1 NAND2X1_1622 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_1_bF_buf0_), .B(micro_hash_ucr_3_pipe59), .Y(_12521_) );
NAND2X1 NAND2X1_1623 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe55), .B(_9483_), .Y(_12522_) );
NOR2X1 NOR2X1_1960 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_5_bF_buf2_), .B(_9298__bF_buf4), .Y(_12523_) );
NAND2X1 NAND2X1_1624 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe53), .B(_9483_), .Y(_12524_) );
NAND2X1 NAND2X1_1625 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_1_bF_buf3_), .B(micro_hash_ucr_3_pipe47), .Y(_12525_) );
NAND2X1 NAND2X1_1626 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_1_bF_buf2_), .B(micro_hash_ucr_3_pipe45_bF_buf3), .Y(_12526_) );
NOR2X1 NOR2X1_1961 ( .gnd(gnd), .vdd(vdd), .A(_8814__bF_buf0), .B(_9312__bF_buf2), .Y(_12527_) );
NAND2X1 NAND2X1_1627 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_1_bF_buf1_), .B(micro_hash_ucr_3_pipe39_bF_buf0), .Y(_12528_) );
NOR2X1 NOR2X1_1962 ( .gnd(gnd), .vdd(vdd), .A(_8814__bF_buf3), .B(_9311__bF_buf4), .Y(_12529_) );
NAND2X1 NAND2X1_1628 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_1_bF_buf0_), .B(micro_hash_ucr_3_pipe37_bF_buf1), .Y(_12530_) );
NOR2X1 NOR2X1_1963 ( .gnd(gnd), .vdd(vdd), .A(_8814__bF_buf2), .B(_9316__bF_buf2), .Y(_12531_) );
NAND2X1 NAND2X1_1629 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_1_bF_buf3_), .B(micro_hash_ucr_3_pipe35_bF_buf2), .Y(_12532_) );
NOR2X1 NOR2X1_1964 ( .gnd(gnd), .vdd(vdd), .A(_9483_), .B(_9321__bF_buf0), .Y(_12533_) );
NAND2X1 NAND2X1_1630 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_5_bF_buf1_), .B(micro_hash_ucr_3_pipe30_bF_buf3), .Y(_12534_) );
NOR2X1 NOR2X1_1965 ( .gnd(gnd), .vdd(vdd), .A(_9483_), .B(_9320_), .Y(_12535_) );
NAND2X1 NAND2X1_1631 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_1_bF_buf2_), .B(micro_hash_ucr_3_pipe25_bF_buf3), .Y(_12536_) );
NAND2X1 NAND2X1_1632 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_5_bF_buf0_), .B(micro_hash_ucr_3_pipe20_bF_buf4), .Y(_12537_) );
NAND2X1 NAND2X1_1633 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_5_bF_buf3_), .B(micro_hash_ucr_3_pipe18_bF_buf3), .Y(_12538_) );
NAND2X1 NAND2X1_1634 ( .gnd(gnd), .vdd(vdd), .A(_8814__bF_buf1), .B(_9626_), .Y(_12539_) );
NAND2X1 NAND2X1_1635 ( .gnd(gnd), .vdd(vdd), .A(_9335__bF_buf3), .B(_9495_), .Y(_12540_) );
NOR2X1 NOR2X1_1966 ( .gnd(gnd), .vdd(vdd), .A(_12540_), .B(_9716_), .Y(_12541_) );
NOR2X1 NOR2X1_1967 ( .gnd(gnd), .vdd(vdd), .A(H_3_13_), .B(micro_hash_ucr_3_pipe10_bF_buf2), .Y(_12542_) );
NAND3X1 NAND3X1_623 ( .gnd(gnd), .vdd(vdd), .A(_10042_), .B(_12542_), .C(_12541_), .Y(_12543_) );
AOI21X1 AOI21X1_2185 ( .gnd(gnd), .vdd(vdd), .A(_12543_), .B(_12539_), .C(micro_hash_ucr_3_pipe15_bF_buf0), .Y(_12544_) );
OAI21X1 OAI21X1_3563 ( .gnd(gnd), .vdd(vdd), .A(_9600_), .B(micro_hash_ucr_3_c_1_bF_buf1_), .C(_9336__bF_buf2), .Y(_12545_) );
OAI22X1 OAI22X1_147 ( .gnd(gnd), .vdd(vdd), .A(_8814__bF_buf0), .B(_9336__bF_buf1), .C(_12544_), .D(_12545_), .Y(_12546_) );
NAND2X1 NAND2X1_1636 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe17_bF_buf2), .B(_9483_), .Y(_12547_) );
OAI21X1 OAI21X1_3564 ( .gnd(gnd), .vdd(vdd), .A(_12546_), .B(micro_hash_ucr_3_pipe17_bF_buf1), .C(_12547_), .Y(_12548_) );
OAI21X1 OAI21X1_3565 ( .gnd(gnd), .vdd(vdd), .A(_12548_), .B(micro_hash_ucr_3_pipe18_bF_buf2), .C(_12538_), .Y(_12549_) );
NAND2X1 NAND2X1_1637 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe19), .B(_9483_), .Y(_12550_) );
OAI21X1 OAI21X1_3566 ( .gnd(gnd), .vdd(vdd), .A(_12549_), .B(micro_hash_ucr_3_pipe19), .C(_12550_), .Y(_12551_) );
OAI21X1 OAI21X1_3567 ( .gnd(gnd), .vdd(vdd), .A(_12551_), .B(micro_hash_ucr_3_pipe20_bF_buf3), .C(_12537_), .Y(_12552_) );
OAI21X1 OAI21X1_3568 ( .gnd(gnd), .vdd(vdd), .A(_9483_), .B(_9331_), .C(_9330__bF_buf2), .Y(_12553_) );
AOI21X1 AOI21X1_2186 ( .gnd(gnd), .vdd(vdd), .A(_9331_), .B(_12552_), .C(_12553_), .Y(_12554_) );
OAI21X1 OAI21X1_3569 ( .gnd(gnd), .vdd(vdd), .A(_9330__bF_buf1), .B(micro_hash_ucr_3_b_5_bF_buf2_), .C(_9326__bF_buf3), .Y(_12555_) );
AOI21X1 AOI21X1_2187 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_1_bF_buf0_), .B(micro_hash_ucr_3_pipe23), .C(micro_hash_ucr_3_pipe24_bF_buf4), .Y(_12556_) );
OAI21X1 OAI21X1_3570 ( .gnd(gnd), .vdd(vdd), .A(_12554_), .B(_12555_), .C(_12556_), .Y(_12557_) );
NAND2X1 NAND2X1_1638 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe24_bF_buf3), .B(_8814__bF_buf3), .Y(_12558_) );
NAND3X1 NAND3X1_624 ( .gnd(gnd), .vdd(vdd), .A(_9327_), .B(_12558_), .C(_12557_), .Y(_12559_) );
AOI21X1 AOI21X1_2188 ( .gnd(gnd), .vdd(vdd), .A(_12536_), .B(_12559_), .C(micro_hash_ucr_3_pipe26_bF_buf2), .Y(_12560_) );
OAI21X1 OAI21X1_3571 ( .gnd(gnd), .vdd(vdd), .A(_8814__bF_buf2), .B(_9323__bF_buf1), .C(_9325__bF_buf3), .Y(_12561_) );
AOI21X1 AOI21X1_2189 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe27), .B(_9483_), .C(micro_hash_ucr_3_pipe28_bF_buf2), .Y(_12562_) );
OAI21X1 OAI21X1_3572 ( .gnd(gnd), .vdd(vdd), .A(_12560_), .B(_12561_), .C(_12562_), .Y(_12563_) );
NAND2X1 NAND2X1_1639 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_5_bF_buf1_), .B(micro_hash_ucr_3_pipe28_bF_buf1), .Y(_12564_) );
AOI21X1 AOI21X1_2190 ( .gnd(gnd), .vdd(vdd), .A(_12564_), .B(_12563_), .C(micro_hash_ucr_3_pipe29_bF_buf2), .Y(_12565_) );
OAI21X1 OAI21X1_3573 ( .gnd(gnd), .vdd(vdd), .A(_12565_), .B(_12535_), .C(_9322__bF_buf1), .Y(_12566_) );
AOI21X1 AOI21X1_2191 ( .gnd(gnd), .vdd(vdd), .A(_12534_), .B(_12566_), .C(micro_hash_ucr_3_pipe31), .Y(_12567_) );
OAI21X1 OAI21X1_3574 ( .gnd(gnd), .vdd(vdd), .A(_12567_), .B(_12533_), .C(_9317__bF_buf0), .Y(_12568_) );
AOI21X1 AOI21X1_2192 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_5_bF_buf0_), .B(micro_hash_ucr_3_pipe32_bF_buf0), .C(micro_hash_ucr_3_pipe33_bF_buf1), .Y(_12569_) );
OAI21X1 OAI21X1_3575 ( .gnd(gnd), .vdd(vdd), .A(_9319_), .B(micro_hash_ucr_3_c_1_bF_buf3_), .C(_9318__bF_buf2), .Y(_12570_) );
AOI21X1 AOI21X1_2193 ( .gnd(gnd), .vdd(vdd), .A(_12569_), .B(_12568_), .C(_12570_), .Y(_12571_) );
NOR2X1 NOR2X1_1968 ( .gnd(gnd), .vdd(vdd), .A(_8814__bF_buf1), .B(_9318__bF_buf1), .Y(_12572_) );
OAI21X1 OAI21X1_3576 ( .gnd(gnd), .vdd(vdd), .A(_12571_), .B(_12572_), .C(_9314_), .Y(_12573_) );
AOI21X1 AOI21X1_2194 ( .gnd(gnd), .vdd(vdd), .A(_12532_), .B(_12573_), .C(micro_hash_ucr_3_pipe36_bF_buf2), .Y(_12574_) );
OAI21X1 OAI21X1_3577 ( .gnd(gnd), .vdd(vdd), .A(_12574_), .B(_12531_), .C(_9315_), .Y(_12575_) );
AOI21X1 AOI21X1_2195 ( .gnd(gnd), .vdd(vdd), .A(_12530_), .B(_12575_), .C(micro_hash_ucr_3_pipe38_bF_buf0), .Y(_12576_) );
OAI21X1 OAI21X1_3578 ( .gnd(gnd), .vdd(vdd), .A(_12576_), .B(_12529_), .C(_9313_), .Y(_12577_) );
AOI21X1 AOI21X1_2196 ( .gnd(gnd), .vdd(vdd), .A(_12528_), .B(_12577_), .C(micro_hash_ucr_3_pipe40_bF_buf2), .Y(_12578_) );
OAI21X1 OAI21X1_3579 ( .gnd(gnd), .vdd(vdd), .A(_12578_), .B(_12527_), .C(_9308_), .Y(_12579_) );
AOI21X1 AOI21X1_2197 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_1_bF_buf2_), .B(micro_hash_ucr_3_pipe41_bF_buf1), .C(micro_hash_ucr_3_pipe42_bF_buf2), .Y(_12580_) );
OAI21X1 OAI21X1_3580 ( .gnd(gnd), .vdd(vdd), .A(_9310__bF_buf1), .B(micro_hash_ucr_3_b_5_bF_buf3_), .C(_9309__bF_buf1), .Y(_12581_) );
AOI21X1 AOI21X1_2198 ( .gnd(gnd), .vdd(vdd), .A(_12580_), .B(_12579_), .C(_12581_), .Y(_12582_) );
OAI21X1 OAI21X1_3581 ( .gnd(gnd), .vdd(vdd), .A(_9483_), .B(_9309__bF_buf0), .C(_9305__bF_buf4), .Y(_12583_) );
OAI22X1 OAI22X1_148 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_5_bF_buf2_), .B(_9305__bF_buf3), .C(_12582_), .D(_12583_), .Y(_12584_) );
OAI21X1 OAI21X1_3582 ( .gnd(gnd), .vdd(vdd), .A(_12584_), .B(micro_hash_ucr_3_pipe45_bF_buf2), .C(_12526_), .Y(_12585_) );
NAND2X1 NAND2X1_1640 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe46_bF_buf1), .B(_8814__bF_buf0), .Y(_12586_) );
OAI21X1 OAI21X1_3583 ( .gnd(gnd), .vdd(vdd), .A(_12585_), .B(micro_hash_ucr_3_pipe46_bF_buf0), .C(_12586_), .Y(_12587_) );
OAI21X1 OAI21X1_3584 ( .gnd(gnd), .vdd(vdd), .A(_12587_), .B(micro_hash_ucr_3_pipe47), .C(_12525_), .Y(_12588_) );
NAND2X1 NAND2X1_1641 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe48_bF_buf1), .B(_8814__bF_buf3), .Y(_12589_) );
OAI21X1 OAI21X1_3585 ( .gnd(gnd), .vdd(vdd), .A(_12588_), .B(micro_hash_ucr_3_pipe48_bF_buf0), .C(_12589_), .Y(_12590_) );
AOI21X1 AOI21X1_2199 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_1_bF_buf1_), .B(micro_hash_ucr_3_pipe49_bF_buf3), .C(micro_hash_ucr_3_pipe50_bF_buf2), .Y(_12591_) );
OAI21X1 OAI21X1_3586 ( .gnd(gnd), .vdd(vdd), .A(_12590_), .B(micro_hash_ucr_3_pipe49_bF_buf2), .C(_12591_), .Y(_12592_) );
AOI21X1 AOI21X1_2200 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe50_bF_buf1), .B(_8814__bF_buf2), .C(micro_hash_ucr_3_pipe51), .Y(_12593_) );
OAI21X1 OAI21X1_3587 ( .gnd(gnd), .vdd(vdd), .A(_9483_), .B(_9301__bF_buf0), .C(_9300__bF_buf3), .Y(_12594_) );
AOI21X1 AOI21X1_2201 ( .gnd(gnd), .vdd(vdd), .A(_12593_), .B(_12592_), .C(_12594_), .Y(_12595_) );
NOR2X1 NOR2X1_1969 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_5_bF_buf1_), .B(_9300__bF_buf2), .Y(_12596_) );
OAI21X1 OAI21X1_3588 ( .gnd(gnd), .vdd(vdd), .A(_12595_), .B(_12596_), .C(_9296_), .Y(_12597_) );
AOI21X1 AOI21X1_2202 ( .gnd(gnd), .vdd(vdd), .A(_12524_), .B(_12597_), .C(micro_hash_ucr_3_pipe54_bF_buf0), .Y(_12598_) );
OAI21X1 OAI21X1_3589 ( .gnd(gnd), .vdd(vdd), .A(_12598_), .B(_12523_), .C(_9297_), .Y(_12599_) );
NAND3X1 NAND3X1_625 ( .gnd(gnd), .vdd(vdd), .A(_9293__bF_buf1), .B(_12522_), .C(_12599_), .Y(_12600_) );
AOI21X1 AOI21X1_2203 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_5_bF_buf0_), .B(micro_hash_ucr_3_pipe56_bF_buf2), .C(micro_hash_ucr_3_pipe57_bF_buf3), .Y(_12601_) );
OAI21X1 OAI21X1_3590 ( .gnd(gnd), .vdd(vdd), .A(_9295_), .B(micro_hash_ucr_3_c_1_bF_buf0_), .C(_9294__bF_buf3), .Y(_12602_) );
AOI21X1 AOI21X1_2204 ( .gnd(gnd), .vdd(vdd), .A(_12601_), .B(_12600_), .C(_12602_), .Y(_12603_) );
NOR2X1 NOR2X1_1970 ( .gnd(gnd), .vdd(vdd), .A(_8814__bF_buf1), .B(_9294__bF_buf2), .Y(_12604_) );
OAI21X1 OAI21X1_3591 ( .gnd(gnd), .vdd(vdd), .A(_12603_), .B(_12604_), .C(_9290__bF_buf1), .Y(_12605_) );
NAND3X1 NAND3X1_626 ( .gnd(gnd), .vdd(vdd), .A(_9292__bF_buf0), .B(_12521_), .C(_12605_), .Y(_12606_) );
NAND3X1 NAND3X1_627 ( .gnd(gnd), .vdd(vdd), .A(_9291_), .B(_12520_), .C(_12606_), .Y(_12607_) );
NAND3X1 NAND3X1_628 ( .gnd(gnd), .vdd(vdd), .A(_9287__bF_buf0), .B(_12519_), .C(_12607_), .Y(_12608_) );
NAND3X1 NAND3X1_629 ( .gnd(gnd), .vdd(vdd), .A(_9289__bF_buf0), .B(_12518_), .C(_12608_), .Y(_12609_) );
NAND3X1 NAND3X1_630 ( .gnd(gnd), .vdd(vdd), .A(_9288__bF_buf0), .B(_12517_), .C(_12609_), .Y(_12610_) );
NAND3X1 NAND3X1_631 ( .gnd(gnd), .vdd(vdd), .A(_9284_), .B(_12516_), .C(_12610_), .Y(_12611_) );
NAND3X1 NAND3X1_632 ( .gnd(gnd), .vdd(vdd), .A(_9286__bF_buf0), .B(_12515_), .C(_12611_), .Y(_12612_) );
NAND3X1 NAND3X1_633 ( .gnd(gnd), .vdd(vdd), .A(_9285__bF_buf1), .B(_12514_), .C(_12612_), .Y(_12613_) );
AOI21X1 AOI21X1_2205 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_1_bF_buf3_), .B(micro_hash_ucr_3_pipe67), .C(micro_hash_ucr_3_pipe68_bF_buf3), .Y(_12614_) );
AND2X2 AND2X2_758 ( .gnd(gnd), .vdd(vdd), .A(_12613_), .B(_12614_), .Y(_12615_) );
OAI21X1 OAI21X1_3592 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_5_bF_buf3_), .B(_9282__bF_buf1), .C(_10380_), .Y(_12616_) );
OAI22X1 OAI22X1_149 ( .gnd(gnd), .vdd(vdd), .A(_9483_), .B(_11524_), .C(_12615_), .D(_12616_), .Y(_8701__5_) );
NAND2X1 NAND2X1_1642 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_2_), .B(micro_hash_ucr_3_pipe63), .Y(_12617_) );
NAND2X1 NAND2X1_1643 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_6_bF_buf2_), .B(micro_hash_ucr_3_pipe60_bF_buf3), .Y(_12618_) );
NAND2X1 NAND2X1_1644 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe59), .B(_9593__bF_buf1), .Y(_12619_) );
NAND2X1 NAND2X1_1645 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_6_bF_buf1_), .B(micro_hash_ucr_3_pipe58_bF_buf1), .Y(_12620_) );
NAND2X1 NAND2X1_1646 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe57_bF_buf2), .B(_9593__bF_buf0), .Y(_12621_) );
NAND2X1 NAND2X1_1647 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_6_bF_buf0_), .B(micro_hash_ucr_3_pipe56_bF_buf1), .Y(_12622_) );
NAND2X1 NAND2X1_1648 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe55), .B(_9593__bF_buf3), .Y(_12623_) );
NAND2X1 NAND2X1_1649 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_6_bF_buf3_), .B(micro_hash_ucr_3_pipe54_bF_buf3), .Y(_12624_) );
NAND2X1 NAND2X1_1650 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe53), .B(_9593__bF_buf2), .Y(_12625_) );
NAND2X1 NAND2X1_1651 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_6_bF_buf2_), .B(micro_hash_ucr_3_pipe52_bF_buf0), .Y(_12626_) );
NAND2X1 NAND2X1_1652 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe51), .B(_9593__bF_buf1), .Y(_12627_) );
NAND2X1 NAND2X1_1653 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_2_), .B(micro_hash_ucr_3_pipe47), .Y(_12628_) );
NAND2X1 NAND2X1_1654 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe46_bF_buf4), .B(_8828_), .Y(_12629_) );
NAND2X1 NAND2X1_1655 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_2_), .B(micro_hash_ucr_3_pipe45_bF_buf1), .Y(_12630_) );
NAND2X1 NAND2X1_1656 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_6_bF_buf1_), .B(micro_hash_ucr_3_pipe36_bF_buf1), .Y(_12631_) );
NAND2X1 NAND2X1_1657 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe35_bF_buf1), .B(_9593__bF_buf0), .Y(_12632_) );
NAND2X1 NAND2X1_1658 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_6_bF_buf0_), .B(micro_hash_ucr_3_pipe34_bF_buf2), .Y(_12633_) );
NAND2X1 NAND2X1_1659 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe33_bF_buf0), .B(_9593__bF_buf3), .Y(_12634_) );
NAND2X1 NAND2X1_1660 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_6_bF_buf3_), .B(micro_hash_ucr_3_pipe32_bF_buf3), .Y(_12635_) );
NAND2X1 NAND2X1_1661 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe31), .B(_9593__bF_buf2), .Y(_12636_) );
NAND2X1 NAND2X1_1662 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_6_bF_buf2_), .B(micro_hash_ucr_3_pipe30_bF_buf2), .Y(_12637_) );
NOR2X1 NOR2X1_1971 ( .gnd(gnd), .vdd(vdd), .A(_9593__bF_buf1), .B(_9320_), .Y(_12638_) );
NAND2X1 NAND2X1_1663 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_6_bF_buf1_), .B(micro_hash_ucr_3_pipe28_bF_buf0), .Y(_12639_) );
NOR2X1 NOR2X1_1972 ( .gnd(gnd), .vdd(vdd), .A(_9593__bF_buf0), .B(_9325__bF_buf2), .Y(_12640_) );
NAND2X1 NAND2X1_1664 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_6_bF_buf0_), .B(micro_hash_ucr_3_pipe26_bF_buf1), .Y(_12641_) );
NOR2X1 NOR2X1_1973 ( .gnd(gnd), .vdd(vdd), .A(_9593__bF_buf3), .B(_9327_), .Y(_12642_) );
NAND2X1 NAND2X1_1665 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_6_bF_buf3_), .B(micro_hash_ucr_3_pipe24_bF_buf2), .Y(_12643_) );
NOR2X1 NOR2X1_1974 ( .gnd(gnd), .vdd(vdd), .A(_9593__bF_buf2), .B(_9326__bF_buf2), .Y(_12644_) );
NAND2X1 NAND2X1_1666 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_6_bF_buf2_), .B(micro_hash_ucr_3_pipe22_bF_buf1), .Y(_12645_) );
NOR2X1 NOR2X1_1975 ( .gnd(gnd), .vdd(vdd), .A(_9593__bF_buf1), .B(_9331_), .Y(_12646_) );
NAND2X1 NAND2X1_1667 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_6_bF_buf1_), .B(micro_hash_ucr_3_pipe20_bF_buf2), .Y(_12647_) );
NAND2X1 NAND2X1_1668 ( .gnd(gnd), .vdd(vdd), .A(_8828_), .B(_9626_), .Y(_12648_) );
NOR2X1 NOR2X1_1976 ( .gnd(gnd), .vdd(vdd), .A(H_3_14_), .B(micro_hash_ucr_3_pipe10_bF_buf1), .Y(_12649_) );
NAND3X1 NAND3X1_634 ( .gnd(gnd), .vdd(vdd), .A(_10042_), .B(_12649_), .C(_12541_), .Y(_12650_) );
AOI21X1 AOI21X1_2206 ( .gnd(gnd), .vdd(vdd), .A(_12650_), .B(_12648_), .C(micro_hash_ucr_3_pipe15_bF_buf3), .Y(_12651_) );
OAI21X1 OAI21X1_3593 ( .gnd(gnd), .vdd(vdd), .A(_9600_), .B(micro_hash_ucr_3_c_2_), .C(_9336__bF_buf0), .Y(_12652_) );
OAI22X1 OAI22X1_150 ( .gnd(gnd), .vdd(vdd), .A(_8828_), .B(_9336__bF_buf3), .C(_12651_), .D(_12652_), .Y(_12653_) );
NAND2X1 NAND2X1_1669 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe17_bF_buf0), .B(_9593__bF_buf0), .Y(_12654_) );
OAI21X1 OAI21X1_3594 ( .gnd(gnd), .vdd(vdd), .A(_12653_), .B(micro_hash_ucr_3_pipe17_bF_buf3), .C(_12654_), .Y(_12655_) );
NOR2X1 NOR2X1_1977 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe18_bF_buf1), .B(_12655_), .Y(_12656_) );
OAI21X1 OAI21X1_3595 ( .gnd(gnd), .vdd(vdd), .A(_8828_), .B(_9334__bF_buf0), .C(_9333__bF_buf3), .Y(_12657_) );
AOI21X1 AOI21X1_2207 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe19), .B(_9593__bF_buf3), .C(micro_hash_ucr_3_pipe20_bF_buf1), .Y(_12658_) );
OAI21X1 OAI21X1_3596 ( .gnd(gnd), .vdd(vdd), .A(_12656_), .B(_12657_), .C(_12658_), .Y(_12659_) );
AOI21X1 AOI21X1_2208 ( .gnd(gnd), .vdd(vdd), .A(_12647_), .B(_12659_), .C(micro_hash_ucr_3_pipe21_bF_buf1), .Y(_12660_) );
OAI21X1 OAI21X1_3597 ( .gnd(gnd), .vdd(vdd), .A(_12660_), .B(_12646_), .C(_9330__bF_buf0), .Y(_12661_) );
AOI21X1 AOI21X1_2209 ( .gnd(gnd), .vdd(vdd), .A(_12645_), .B(_12661_), .C(micro_hash_ucr_3_pipe23), .Y(_12662_) );
OAI21X1 OAI21X1_3598 ( .gnd(gnd), .vdd(vdd), .A(_12662_), .B(_12644_), .C(_9328__bF_buf0), .Y(_12663_) );
AOI21X1 AOI21X1_2210 ( .gnd(gnd), .vdd(vdd), .A(_12643_), .B(_12663_), .C(micro_hash_ucr_3_pipe25_bF_buf2), .Y(_12664_) );
OAI21X1 OAI21X1_3599 ( .gnd(gnd), .vdd(vdd), .A(_12664_), .B(_12642_), .C(_9323__bF_buf0), .Y(_12665_) );
AOI21X1 AOI21X1_2211 ( .gnd(gnd), .vdd(vdd), .A(_12641_), .B(_12665_), .C(micro_hash_ucr_3_pipe27), .Y(_12666_) );
OAI21X1 OAI21X1_3600 ( .gnd(gnd), .vdd(vdd), .A(_12666_), .B(_12640_), .C(_9324__bF_buf2), .Y(_12667_) );
AOI21X1 AOI21X1_2212 ( .gnd(gnd), .vdd(vdd), .A(_12639_), .B(_12667_), .C(micro_hash_ucr_3_pipe29_bF_buf1), .Y(_12668_) );
OAI21X1 OAI21X1_3601 ( .gnd(gnd), .vdd(vdd), .A(_12668_), .B(_12638_), .C(_9322__bF_buf0), .Y(_12669_) );
NAND3X1 NAND3X1_635 ( .gnd(gnd), .vdd(vdd), .A(_9321__bF_buf3), .B(_12637_), .C(_12669_), .Y(_12670_) );
NAND3X1 NAND3X1_636 ( .gnd(gnd), .vdd(vdd), .A(_9317__bF_buf4), .B(_12636_), .C(_12670_), .Y(_12671_) );
NAND3X1 NAND3X1_637 ( .gnd(gnd), .vdd(vdd), .A(_9319_), .B(_12635_), .C(_12671_), .Y(_12672_) );
NAND3X1 NAND3X1_638 ( .gnd(gnd), .vdd(vdd), .A(_9318__bF_buf0), .B(_12634_), .C(_12672_), .Y(_12673_) );
NAND3X1 NAND3X1_639 ( .gnd(gnd), .vdd(vdd), .A(_9314_), .B(_12633_), .C(_12673_), .Y(_12674_) );
NAND3X1 NAND3X1_640 ( .gnd(gnd), .vdd(vdd), .A(_9316__bF_buf1), .B(_12632_), .C(_12674_), .Y(_12675_) );
AOI21X1 AOI21X1_2213 ( .gnd(gnd), .vdd(vdd), .A(_12631_), .B(_12675_), .C(micro_hash_ucr_3_pipe37_bF_buf0), .Y(_12676_) );
OAI21X1 OAI21X1_3602 ( .gnd(gnd), .vdd(vdd), .A(_9593__bF_buf2), .B(_9315_), .C(_9311__bF_buf3), .Y(_12677_) );
AOI21X1 AOI21X1_2214 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe38_bF_buf3), .B(_8828_), .C(micro_hash_ucr_3_pipe39_bF_buf3), .Y(_12678_) );
OAI21X1 OAI21X1_3603 ( .gnd(gnd), .vdd(vdd), .A(_12676_), .B(_12677_), .C(_12678_), .Y(_12679_) );
AOI21X1 AOI21X1_2215 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_2_), .B(micro_hash_ucr_3_pipe39_bF_buf2), .C(micro_hash_ucr_3_pipe40_bF_buf1), .Y(_12680_) );
AOI22X1 AOI22X1_89 ( .gnd(gnd), .vdd(vdd), .A(_8828_), .B(micro_hash_ucr_3_pipe40_bF_buf0), .C(_12679_), .D(_12680_), .Y(_12681_) );
OAI21X1 OAI21X1_3604 ( .gnd(gnd), .vdd(vdd), .A(_9593__bF_buf1), .B(_9308_), .C(_9310__bF_buf0), .Y(_12682_) );
AOI21X1 AOI21X1_2216 ( .gnd(gnd), .vdd(vdd), .A(_9308_), .B(_12681_), .C(_12682_), .Y(_12683_) );
OAI21X1 OAI21X1_3605 ( .gnd(gnd), .vdd(vdd), .A(_9310__bF_buf4), .B(micro_hash_ucr_3_b_6_bF_buf0_), .C(_9309__bF_buf3), .Y(_12684_) );
AOI21X1 AOI21X1_2217 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_2_), .B(micro_hash_ucr_3_pipe43), .C(micro_hash_ucr_3_pipe44_bF_buf0), .Y(_12685_) );
OAI21X1 OAI21X1_3606 ( .gnd(gnd), .vdd(vdd), .A(_12683_), .B(_12684_), .C(_12685_), .Y(_12686_) );
NAND2X1 NAND2X1_1670 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe44_bF_buf3), .B(_8828_), .Y(_12687_) );
NAND3X1 NAND3X1_641 ( .gnd(gnd), .vdd(vdd), .A(_9307_), .B(_12687_), .C(_12686_), .Y(_12688_) );
NAND3X1 NAND3X1_642 ( .gnd(gnd), .vdd(vdd), .A(_9306__bF_buf3), .B(_12630_), .C(_12688_), .Y(_12689_) );
NAND3X1 NAND3X1_643 ( .gnd(gnd), .vdd(vdd), .A(_9302_), .B(_12629_), .C(_12689_), .Y(_12690_) );
AOI21X1 AOI21X1_2218 ( .gnd(gnd), .vdd(vdd), .A(_12628_), .B(_12690_), .C(micro_hash_ucr_3_pipe48_bF_buf4), .Y(_12691_) );
OAI21X1 OAI21X1_3607 ( .gnd(gnd), .vdd(vdd), .A(_8828_), .B(_9304__bF_buf2), .C(_9303_), .Y(_12692_) );
AOI21X1 AOI21X1_2219 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe49_bF_buf1), .B(_9593__bF_buf0), .C(micro_hash_ucr_3_pipe50_bF_buf0), .Y(_12693_) );
OAI21X1 OAI21X1_3608 ( .gnd(gnd), .vdd(vdd), .A(_12691_), .B(_12692_), .C(_12693_), .Y(_12694_) );
NAND2X1 NAND2X1_1671 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_6_bF_buf3_), .B(micro_hash_ucr_3_pipe50_bF_buf4), .Y(_12695_) );
NAND3X1 NAND3X1_644 ( .gnd(gnd), .vdd(vdd), .A(_9301__bF_buf3), .B(_12695_), .C(_12694_), .Y(_12696_) );
NAND3X1 NAND3X1_645 ( .gnd(gnd), .vdd(vdd), .A(_9300__bF_buf1), .B(_12627_), .C(_12696_), .Y(_12697_) );
NAND3X1 NAND3X1_646 ( .gnd(gnd), .vdd(vdd), .A(_9296_), .B(_12626_), .C(_12697_), .Y(_12698_) );
NAND3X1 NAND3X1_647 ( .gnd(gnd), .vdd(vdd), .A(_9298__bF_buf3), .B(_12625_), .C(_12698_), .Y(_12699_) );
NAND3X1 NAND3X1_648 ( .gnd(gnd), .vdd(vdd), .A(_9297_), .B(_12624_), .C(_12699_), .Y(_12700_) );
NAND3X1 NAND3X1_649 ( .gnd(gnd), .vdd(vdd), .A(_9293__bF_buf0), .B(_12623_), .C(_12700_), .Y(_12701_) );
NAND3X1 NAND3X1_650 ( .gnd(gnd), .vdd(vdd), .A(_9295_), .B(_12622_), .C(_12701_), .Y(_12702_) );
NAND3X1 NAND3X1_651 ( .gnd(gnd), .vdd(vdd), .A(_9294__bF_buf1), .B(_12621_), .C(_12702_), .Y(_12703_) );
NAND3X1 NAND3X1_652 ( .gnd(gnd), .vdd(vdd), .A(_9290__bF_buf0), .B(_12620_), .C(_12703_), .Y(_12704_) );
NAND3X1 NAND3X1_653 ( .gnd(gnd), .vdd(vdd), .A(_9292__bF_buf3), .B(_12619_), .C(_12704_), .Y(_12705_) );
AOI21X1 AOI21X1_2220 ( .gnd(gnd), .vdd(vdd), .A(_12618_), .B(_12705_), .C(micro_hash_ucr_3_pipe61_bF_buf0), .Y(_12706_) );
OAI21X1 OAI21X1_3609 ( .gnd(gnd), .vdd(vdd), .A(_9593__bF_buf3), .B(_9291_), .C(_9287__bF_buf4), .Y(_12707_) );
AOI21X1 AOI21X1_2221 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe62_bF_buf2), .B(_8828_), .C(micro_hash_ucr_3_pipe63), .Y(_12708_) );
OAI21X1 OAI21X1_3610 ( .gnd(gnd), .vdd(vdd), .A(_12706_), .B(_12707_), .C(_12708_), .Y(_12709_) );
NAND2X1 NAND2X1_1672 ( .gnd(gnd), .vdd(vdd), .A(_12617_), .B(_12709_), .Y(_12710_) );
OAI21X1 OAI21X1_3611 ( .gnd(gnd), .vdd(vdd), .A(_8828_), .B(_9288__bF_buf3), .C(_9284_), .Y(_12711_) );
AOI21X1 AOI21X1_2222 ( .gnd(gnd), .vdd(vdd), .A(_9288__bF_buf2), .B(_12710_), .C(_12711_), .Y(_12712_) );
OAI21X1 OAI21X1_3612 ( .gnd(gnd), .vdd(vdd), .A(_9284_), .B(micro_hash_ucr_3_c_2_), .C(_9286__bF_buf3), .Y(_12713_) );
NAND2X1 NAND2X1_1673 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_6_bF_buf2_), .B(micro_hash_ucr_3_pipe66_bF_buf3), .Y(_12714_) );
OAI21X1 OAI21X1_3613 ( .gnd(gnd), .vdd(vdd), .A(_12712_), .B(_12713_), .C(_12714_), .Y(_12715_) );
OAI21X1 OAI21X1_3614 ( .gnd(gnd), .vdd(vdd), .A(_9593__bF_buf2), .B(_9285__bF_buf0), .C(_9282__bF_buf0), .Y(_12716_) );
AOI21X1 AOI21X1_2223 ( .gnd(gnd), .vdd(vdd), .A(_9285__bF_buf3), .B(_12715_), .C(_12716_), .Y(_12717_) );
OAI21X1 OAI21X1_3615 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_6_bF_buf1_), .B(_9282__bF_buf4), .C(_10380_), .Y(_12718_) );
OAI22X1 OAI22X1_151 ( .gnd(gnd), .vdd(vdd), .A(_9593__bF_buf1), .B(_11524_), .C(_12717_), .D(_12718_), .Y(_8701__6_) );
NAND2X1 NAND2X1_1674 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe63), .B(_9701__bF_buf1), .Y(_12719_) );
NAND2X1 NAND2X1_1675 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_7_bF_buf2_), .B(micro_hash_ucr_3_pipe62_bF_buf1), .Y(_12720_) );
NAND2X1 NAND2X1_1676 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe61_bF_buf3), .B(_9701__bF_buf0), .Y(_12721_) );
NAND2X1 NAND2X1_1677 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_3_bF_buf3_), .B(micro_hash_ucr_3_pipe57_bF_buf1), .Y(_12722_) );
NAND2X1 NAND2X1_1678 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_7_bF_buf1_), .B(micro_hash_ucr_3_pipe52_bF_buf4), .Y(_12723_) );
NAND2X1 NAND2X1_1679 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_7_bF_buf0_), .B(micro_hash_ucr_3_pipe50_bF_buf3), .Y(_12724_) );
INVX8 INVX8_286 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_7_bF_buf3_), .Y(_12725_) );
NOR2X1 NOR2X1_1978 ( .gnd(gnd), .vdd(vdd), .A(_9701__bF_buf3), .B(_9309__bF_buf2), .Y(_12726_) );
NAND2X1 NAND2X1_1680 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_7_bF_buf2_), .B(micro_hash_ucr_3_pipe42_bF_buf1), .Y(_12727_) );
NOR2X1 NOR2X1_1979 ( .gnd(gnd), .vdd(vdd), .A(_9701__bF_buf2), .B(_9308_), .Y(_12728_) );
NAND2X1 NAND2X1_1681 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_3_bF_buf2_), .B(micro_hash_ucr_3_pipe33_bF_buf3), .Y(_12729_) );
NAND2X1 NAND2X1_1682 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe29_bF_buf0), .B(_9701__bF_buf1), .Y(_12730_) );
NAND2X1 NAND2X1_1683 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_3_bF_buf1_), .B(micro_hash_ucr_3_pipe27), .Y(_12731_) );
NAND2X1 NAND2X1_1684 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_3_bF_buf0_), .B(micro_hash_ucr_3_pipe25_bF_buf1), .Y(_12732_) );
NOR2X1 NOR2X1_1980 ( .gnd(gnd), .vdd(vdd), .A(_12725_), .B(_9329__bF_buf4), .Y(_12733_) );
NAND2X1 NAND2X1_1685 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_3_bF_buf3_), .B(micro_hash_ucr_3_pipe19), .Y(_12734_) );
NOR2X1 NOR2X1_1981 ( .gnd(gnd), .vdd(vdd), .A(_12725_), .B(_9334__bF_buf3), .Y(_12735_) );
NAND2X1 NAND2X1_1686 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_3_bF_buf2_), .B(micro_hash_ucr_3_pipe17_bF_buf2), .Y(_12736_) );
NOR2X1 NOR2X1_1982 ( .gnd(gnd), .vdd(vdd), .A(_12725_), .B(_9336__bF_buf2), .Y(_12737_) );
NAND2X1 NAND2X1_1687 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_7_bF_buf1_), .B(micro_hash_ucr_3_pipe14_bF_buf0), .Y(_12738_) );
INVX1 INVX1_844 ( .gnd(gnd), .vdd(vdd), .A(_9495_), .Y(_12739_) );
NOR2X1 NOR2X1_1983 ( .gnd(gnd), .vdd(vdd), .A(_9489_), .B(_9374_), .Y(_12740_) );
NOR2X1 NOR2X1_1984 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_7_bF_buf0_), .B(micro_hash_ucr_3_pipe11), .Y(_12741_) );
OAI21X1 OAI21X1_3616 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe10_bF_buf0), .B(_9343_), .C(_12741_), .Y(_12742_) );
NOR2X1 NOR2X1_1985 ( .gnd(gnd), .vdd(vdd), .A(H_3_15_), .B(micro_hash_ucr_3_pipe10_bF_buf3), .Y(_12743_) );
NAND3X1 NAND3X1_654 ( .gnd(gnd), .vdd(vdd), .A(_9343_), .B(_10042_), .C(_12743_), .Y(_12744_) );
OAI22X1 OAI22X1_152 ( .gnd(gnd), .vdd(vdd), .A(_9488_), .B(_12744_), .C(_12740_), .D(_12742_), .Y(_12745_) );
AOI22X1 AOI22X1_90 ( .gnd(gnd), .vdd(vdd), .A(_9701__bF_buf0), .B(_9838_), .C(_12745_), .D(_9337_), .Y(_12746_) );
NOR2X1 NOR2X1_1986 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_7_bF_buf3_), .B(_9379_), .Y(_12747_) );
OAI21X1 OAI21X1_3617 ( .gnd(gnd), .vdd(vdd), .A(_9339_), .B(micro_hash_ucr_3_c_3_bF_buf1_), .C(_9335__bF_buf2), .Y(_12748_) );
OAI21X1 OAI21X1_3618 ( .gnd(gnd), .vdd(vdd), .A(_12747_), .B(_12748_), .C(_9337_), .Y(_12749_) );
OAI21X1 OAI21X1_3619 ( .gnd(gnd), .vdd(vdd), .A(_12746_), .B(_12739_), .C(_12749_), .Y(_12750_) );
OAI21X1 OAI21X1_3620 ( .gnd(gnd), .vdd(vdd), .A(_9337_), .B(micro_hash_ucr_3_c_3_bF_buf0_), .C(_9336__bF_buf1), .Y(_12751_) );
AOI21X1 AOI21X1_2224 ( .gnd(gnd), .vdd(vdd), .A(_12738_), .B(_12750_), .C(_12751_), .Y(_12752_) );
OAI21X1 OAI21X1_3621 ( .gnd(gnd), .vdd(vdd), .A(_12752_), .B(_12737_), .C(_9332_), .Y(_12753_) );
AOI21X1 AOI21X1_2225 ( .gnd(gnd), .vdd(vdd), .A(_12736_), .B(_12753_), .C(micro_hash_ucr_3_pipe18_bF_buf0), .Y(_12754_) );
OAI21X1 OAI21X1_3622 ( .gnd(gnd), .vdd(vdd), .A(_12754_), .B(_12735_), .C(_9333__bF_buf2), .Y(_12755_) );
AOI21X1 AOI21X1_2226 ( .gnd(gnd), .vdd(vdd), .A(_12734_), .B(_12755_), .C(micro_hash_ucr_3_pipe20_bF_buf0), .Y(_12756_) );
OAI21X1 OAI21X1_3623 ( .gnd(gnd), .vdd(vdd), .A(_12756_), .B(_12733_), .C(_9331_), .Y(_12757_) );
AOI21X1 AOI21X1_2227 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_3_bF_buf3_), .B(micro_hash_ucr_3_pipe21_bF_buf0), .C(micro_hash_ucr_3_pipe22_bF_buf0), .Y(_12758_) );
OAI21X1 OAI21X1_3624 ( .gnd(gnd), .vdd(vdd), .A(_9330__bF_buf4), .B(micro_hash_ucr_3_b_7_bF_buf2_), .C(_9326__bF_buf1), .Y(_12759_) );
AOI21X1 AOI21X1_2228 ( .gnd(gnd), .vdd(vdd), .A(_12758_), .B(_12757_), .C(_12759_), .Y(_12760_) );
OAI21X1 OAI21X1_3625 ( .gnd(gnd), .vdd(vdd), .A(_9701__bF_buf3), .B(_9326__bF_buf0), .C(_9328__bF_buf3), .Y(_12761_) );
OAI22X1 OAI22X1_153 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_7_bF_buf1_), .B(_9328__bF_buf2), .C(_12760_), .D(_12761_), .Y(_12762_) );
OAI21X1 OAI21X1_3626 ( .gnd(gnd), .vdd(vdd), .A(_12762_), .B(micro_hash_ucr_3_pipe25_bF_buf0), .C(_12732_), .Y(_12763_) );
NAND2X1 NAND2X1_1688 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe26_bF_buf0), .B(_12725_), .Y(_12764_) );
OAI21X1 OAI21X1_3627 ( .gnd(gnd), .vdd(vdd), .A(_12763_), .B(micro_hash_ucr_3_pipe26_bF_buf4), .C(_12764_), .Y(_12765_) );
OAI21X1 OAI21X1_3628 ( .gnd(gnd), .vdd(vdd), .A(_12765_), .B(micro_hash_ucr_3_pipe27), .C(_12731_), .Y(_12766_) );
NAND2X1 NAND2X1_1689 ( .gnd(gnd), .vdd(vdd), .A(_9324__bF_buf1), .B(_12766_), .Y(_12767_) );
OAI21X1 OAI21X1_3629 ( .gnd(gnd), .vdd(vdd), .A(_12725_), .B(_9324__bF_buf0), .C(_12767_), .Y(_12768_) );
OAI21X1 OAI21X1_3630 ( .gnd(gnd), .vdd(vdd), .A(_12768_), .B(micro_hash_ucr_3_pipe29_bF_buf3), .C(_12730_), .Y(_12769_) );
OAI21X1 OAI21X1_3631 ( .gnd(gnd), .vdd(vdd), .A(_9322__bF_buf3), .B(micro_hash_ucr_3_b_7_bF_buf0_), .C(_9321__bF_buf2), .Y(_12770_) );
AOI21X1 AOI21X1_2229 ( .gnd(gnd), .vdd(vdd), .A(_9322__bF_buf2), .B(_12769_), .C(_12770_), .Y(_12771_) );
OAI21X1 OAI21X1_3632 ( .gnd(gnd), .vdd(vdd), .A(_9701__bF_buf2), .B(_9321__bF_buf1), .C(_9317__bF_buf3), .Y(_12772_) );
OAI22X1 OAI22X1_154 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_7_bF_buf3_), .B(_9317__bF_buf2), .C(_12771_), .D(_12772_), .Y(_12773_) );
OAI21X1 OAI21X1_3633 ( .gnd(gnd), .vdd(vdd), .A(_12773_), .B(micro_hash_ucr_3_pipe33_bF_buf2), .C(_12729_), .Y(_12774_) );
NAND2X1 NAND2X1_1690 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe34_bF_buf1), .B(_12725_), .Y(_12775_) );
OAI21X1 OAI21X1_3634 ( .gnd(gnd), .vdd(vdd), .A(_12774_), .B(micro_hash_ucr_3_pipe34_bF_buf0), .C(_12775_), .Y(_12776_) );
NAND2X1 NAND2X1_1691 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_3_bF_buf2_), .B(micro_hash_ucr_3_pipe35_bF_buf0), .Y(_12777_) );
OAI21X1 OAI21X1_3635 ( .gnd(gnd), .vdd(vdd), .A(_12776_), .B(micro_hash_ucr_3_pipe35_bF_buf3), .C(_12777_), .Y(_12778_) );
AOI21X1 AOI21X1_2230 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe36_bF_buf0), .B(_12725_), .C(micro_hash_ucr_3_pipe37_bF_buf3), .Y(_12779_) );
OAI21X1 OAI21X1_3636 ( .gnd(gnd), .vdd(vdd), .A(_12778_), .B(micro_hash_ucr_3_pipe36_bF_buf4), .C(_12779_), .Y(_12780_) );
AOI21X1 AOI21X1_2231 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_3_bF_buf1_), .B(micro_hash_ucr_3_pipe37_bF_buf2), .C(micro_hash_ucr_3_pipe38_bF_buf2), .Y(_12781_) );
AOI22X1 AOI22X1_91 ( .gnd(gnd), .vdd(vdd), .A(_12725_), .B(micro_hash_ucr_3_pipe38_bF_buf1), .C(_12780_), .D(_12781_), .Y(_12782_) );
AOI21X1 AOI21X1_2232 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe39_bF_buf1), .B(_9701__bF_buf1), .C(micro_hash_ucr_3_pipe40_bF_buf4), .Y(_12783_) );
OAI21X1 OAI21X1_3637 ( .gnd(gnd), .vdd(vdd), .A(_12782_), .B(micro_hash_ucr_3_pipe39_bF_buf0), .C(_12783_), .Y(_12784_) );
NAND2X1 NAND2X1_1692 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_7_bF_buf2_), .B(micro_hash_ucr_3_pipe40_bF_buf3), .Y(_12785_) );
AOI21X1 AOI21X1_2233 ( .gnd(gnd), .vdd(vdd), .A(_12785_), .B(_12784_), .C(micro_hash_ucr_3_pipe41_bF_buf0), .Y(_12786_) );
OAI21X1 OAI21X1_3638 ( .gnd(gnd), .vdd(vdd), .A(_12786_), .B(_12728_), .C(_9310__bF_buf3), .Y(_12787_) );
AOI21X1 AOI21X1_2234 ( .gnd(gnd), .vdd(vdd), .A(_12727_), .B(_12787_), .C(micro_hash_ucr_3_pipe43), .Y(_12788_) );
OAI21X1 OAI21X1_3639 ( .gnd(gnd), .vdd(vdd), .A(_12788_), .B(_12726_), .C(_9305__bF_buf2), .Y(_12789_) );
OAI21X1 OAI21X1_3640 ( .gnd(gnd), .vdd(vdd), .A(_12725_), .B(_9305__bF_buf1), .C(_12789_), .Y(_12790_) );
AND2X2 AND2X2_759 ( .gnd(gnd), .vdd(vdd), .A(_12790_), .B(_9307_), .Y(_12791_) );
OAI21X1 OAI21X1_3641 ( .gnd(gnd), .vdd(vdd), .A(_9701__bF_buf0), .B(_9307_), .C(_9306__bF_buf2), .Y(_12792_) );
AOI21X1 AOI21X1_2235 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe46_bF_buf3), .B(_12725_), .C(micro_hash_ucr_3_pipe47), .Y(_12793_) );
OAI21X1 OAI21X1_3642 ( .gnd(gnd), .vdd(vdd), .A(_12791_), .B(_12792_), .C(_12793_), .Y(_12794_) );
AOI21X1 AOI21X1_2236 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_3_bF_buf0_), .B(micro_hash_ucr_3_pipe47), .C(micro_hash_ucr_3_pipe48_bF_buf3), .Y(_12795_) );
AOI22X1 AOI22X1_92 ( .gnd(gnd), .vdd(vdd), .A(_12725_), .B(micro_hash_ucr_3_pipe48_bF_buf2), .C(_12794_), .D(_12795_), .Y(_12796_) );
NAND2X1 NAND2X1_1693 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe49_bF_buf0), .B(_9701__bF_buf3), .Y(_12797_) );
OAI21X1 OAI21X1_3643 ( .gnd(gnd), .vdd(vdd), .A(_12796_), .B(micro_hash_ucr_3_pipe49_bF_buf3), .C(_12797_), .Y(_12798_) );
OAI21X1 OAI21X1_3644 ( .gnd(gnd), .vdd(vdd), .A(_12798_), .B(micro_hash_ucr_3_pipe50_bF_buf2), .C(_12724_), .Y(_12799_) );
NAND2X1 NAND2X1_1694 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe51), .B(_9701__bF_buf2), .Y(_12800_) );
OAI21X1 OAI21X1_3645 ( .gnd(gnd), .vdd(vdd), .A(_12799_), .B(micro_hash_ucr_3_pipe51), .C(_12800_), .Y(_12801_) );
OAI21X1 OAI21X1_3646 ( .gnd(gnd), .vdd(vdd), .A(_12801_), .B(micro_hash_ucr_3_pipe52_bF_buf3), .C(_12723_), .Y(_12802_) );
OAI21X1 OAI21X1_3647 ( .gnd(gnd), .vdd(vdd), .A(_9701__bF_buf1), .B(_9296_), .C(_9298__bF_buf2), .Y(_12803_) );
AOI21X1 AOI21X1_2237 ( .gnd(gnd), .vdd(vdd), .A(_9296_), .B(_12802_), .C(_12803_), .Y(_12804_) );
OAI21X1 OAI21X1_3648 ( .gnd(gnd), .vdd(vdd), .A(_9298__bF_buf1), .B(micro_hash_ucr_3_b_7_bF_buf1_), .C(_9297_), .Y(_12805_) );
AOI21X1 AOI21X1_2238 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_3_bF_buf3_), .B(micro_hash_ucr_3_pipe55), .C(micro_hash_ucr_3_pipe56_bF_buf0), .Y(_12806_) );
OAI21X1 OAI21X1_3649 ( .gnd(gnd), .vdd(vdd), .A(_12804_), .B(_12805_), .C(_12806_), .Y(_12807_) );
NAND2X1 NAND2X1_1695 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe56_bF_buf4), .B(_12725_), .Y(_12808_) );
NAND3X1 NAND3X1_655 ( .gnd(gnd), .vdd(vdd), .A(_9295_), .B(_12808_), .C(_12807_), .Y(_12809_) );
AOI21X1 AOI21X1_2239 ( .gnd(gnd), .vdd(vdd), .A(_12722_), .B(_12809_), .C(micro_hash_ucr_3_pipe58_bF_buf0), .Y(_12810_) );
OAI21X1 OAI21X1_3650 ( .gnd(gnd), .vdd(vdd), .A(_12725_), .B(_9294__bF_buf0), .C(_9290__bF_buf3), .Y(_12811_) );
AOI21X1 AOI21X1_2240 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe59), .B(_9701__bF_buf0), .C(micro_hash_ucr_3_pipe60_bF_buf2), .Y(_12812_) );
OAI21X1 OAI21X1_3651 ( .gnd(gnd), .vdd(vdd), .A(_12810_), .B(_12811_), .C(_12812_), .Y(_12813_) );
NAND2X1 NAND2X1_1696 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_7_bF_buf0_), .B(micro_hash_ucr_3_pipe60_bF_buf1), .Y(_12814_) );
NAND3X1 NAND3X1_656 ( .gnd(gnd), .vdd(vdd), .A(_9291_), .B(_12814_), .C(_12813_), .Y(_12815_) );
NAND3X1 NAND3X1_657 ( .gnd(gnd), .vdd(vdd), .A(_9287__bF_buf3), .B(_12721_), .C(_12815_), .Y(_12816_) );
NAND3X1 NAND3X1_658 ( .gnd(gnd), .vdd(vdd), .A(_9289__bF_buf3), .B(_12720_), .C(_12816_), .Y(_12817_) );
NAND3X1 NAND3X1_659 ( .gnd(gnd), .vdd(vdd), .A(_9288__bF_buf1), .B(_12719_), .C(_12817_), .Y(_12818_) );
AOI21X1 AOI21X1_2241 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_7_bF_buf3_), .B(micro_hash_ucr_3_pipe64_bF_buf3), .C(micro_hash_ucr_3_pipe65_bF_buf3), .Y(_12819_) );
AOI22X1 AOI22X1_93 ( .gnd(gnd), .vdd(vdd), .A(_9701__bF_buf3), .B(micro_hash_ucr_3_pipe65_bF_buf2), .C(_12818_), .D(_12819_), .Y(_12820_) );
AOI21X1 AOI21X1_2242 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe66_bF_buf2), .B(_12725_), .C(micro_hash_ucr_3_pipe67), .Y(_12821_) );
OAI21X1 OAI21X1_3652 ( .gnd(gnd), .vdd(vdd), .A(_12820_), .B(micro_hash_ucr_3_pipe66_bF_buf1), .C(_12821_), .Y(_12822_) );
AOI21X1 AOI21X1_2243 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_c_3_bF_buf2_), .B(micro_hash_ucr_3_pipe67), .C(micro_hash_ucr_3_pipe68_bF_buf2), .Y(_12823_) );
AND2X2 AND2X2_760 ( .gnd(gnd), .vdd(vdd), .A(_12822_), .B(_12823_), .Y(_12824_) );
OAI21X1 OAI21X1_3653 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_b_7_bF_buf2_), .B(_9282__bF_buf3), .C(_10380_), .Y(_12825_) );
OAI22X1 OAI22X1_155 ( .gnd(gnd), .vdd(vdd), .A(_9701__bF_buf2), .B(_11524_), .C(_12824_), .D(_12825_), .Y(_8701__7_) );
AOI21X1 AOI21X1_2244 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_176_), .B(_9183_), .C(micro_hash_ucr_3_Wx_224_), .Y(_12826_) );
OAI21X1 OAI21X1_3654 ( .gnd(gnd), .vdd(vdd), .A(_9183_), .B(micro_hash_ucr_3_Wx_176_), .C(_12826_), .Y(_12827_) );
AND2X2 AND2X2_761 ( .gnd(gnd), .vdd(vdd), .A(_12827_), .B(_8705__bF_buf1), .Y(_8699__248_) );
OAI21X1 OAI21X1_3655 ( .gnd(gnd), .vdd(vdd), .A(_9187_), .B(micro_hash_ucr_3_Wx_177_), .C(_10699_), .Y(_12828_) );
AOI21X1 AOI21X1_2245 ( .gnd(gnd), .vdd(vdd), .A(_9187_), .B(micro_hash_ucr_3_Wx_177_), .C(_12828_), .Y(_12829_) );
NOR2X1 NOR2X1_1987 ( .gnd(gnd), .vdd(vdd), .A(_12829_), .B(_8800__bF_buf1), .Y(_8699__249_) );
OAI21X1 OAI21X1_3656 ( .gnd(gnd), .vdd(vdd), .A(_9191_), .B(micro_hash_ucr_3_Wx_178_), .C(_10959_), .Y(_12830_) );
AOI21X1 AOI21X1_2246 ( .gnd(gnd), .vdd(vdd), .A(_9191_), .B(micro_hash_ucr_3_Wx_178_), .C(_12830_), .Y(_12831_) );
NOR2X1 NOR2X1_1988 ( .gnd(gnd), .vdd(vdd), .A(_12831_), .B(_8800__bF_buf0), .Y(_8699__250_) );
OAI21X1 OAI21X1_3657 ( .gnd(gnd), .vdd(vdd), .A(_9195_), .B(micro_hash_ucr_3_Wx_179_), .C(_11246_), .Y(_12832_) );
AOI21X1 AOI21X1_2247 ( .gnd(gnd), .vdd(vdd), .A(_9195_), .B(micro_hash_ucr_3_Wx_179_), .C(_12832_), .Y(_12833_) );
NOR2X1 NOR2X1_1989 ( .gnd(gnd), .vdd(vdd), .A(_12833_), .B(_8800__bF_buf12), .Y(_8699__251_) );
AOI21X1 AOI21X1_2248 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_180_), .B(_9199_), .C(micro_hash_ucr_3_Wx_228_), .Y(_12834_) );
OAI21X1 OAI21X1_3658 ( .gnd(gnd), .vdd(vdd), .A(_9199_), .B(micro_hash_ucr_3_Wx_180_), .C(_12834_), .Y(_12835_) );
AND2X2 AND2X2_762 ( .gnd(gnd), .vdd(vdd), .A(_12835_), .B(_8705__bF_buf0), .Y(_8699__252_) );
OAI21X1 OAI21X1_3659 ( .gnd(gnd), .vdd(vdd), .A(_9203_), .B(micro_hash_ucr_3_Wx_181_), .C(_11760_), .Y(_12836_) );
AOI21X1 AOI21X1_2249 ( .gnd(gnd), .vdd(vdd), .A(_9203_), .B(micro_hash_ucr_3_Wx_181_), .C(_12836_), .Y(_12837_) );
NOR2X1 NOR2X1_1990 ( .gnd(gnd), .vdd(vdd), .A(_12837_), .B(_8800__bF_buf11), .Y(_8699__253_) );
OAI21X1 OAI21X1_3660 ( .gnd(gnd), .vdd(vdd), .A(_9207_), .B(micro_hash_ucr_3_Wx_182_), .C(_11971_), .Y(_12838_) );
AOI21X1 AOI21X1_2250 ( .gnd(gnd), .vdd(vdd), .A(_9207_), .B(micro_hash_ucr_3_Wx_182_), .C(_12838_), .Y(_12839_) );
NOR2X1 NOR2X1_1991 ( .gnd(gnd), .vdd(vdd), .A(_12839_), .B(_8800__bF_buf10), .Y(_8699__254_) );
AOI21X1 AOI21X1_2251 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_Wx_183_), .B(_9211_), .C(micro_hash_ucr_3_Wx_231_), .Y(_12840_) );
OAI21X1 OAI21X1_3661 ( .gnd(gnd), .vdd(vdd), .A(_9211_), .B(micro_hash_ucr_3_Wx_183_), .C(_12840_), .Y(_12841_) );
AND2X2 AND2X2_763 ( .gnd(gnd), .vdd(vdd), .A(_12841_), .B(_8705__bF_buf13), .Y(_8699__255_) );
OAI21X1 OAI21X1_3662 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe70_bF_buf1), .B(comparador_3_valid_hash), .C(_8705__bF_buf12), .Y(_12842_) );
NOR2X1 NOR2X1_1992 ( .gnd(gnd), .vdd(vdd), .A(micro_hash_ucr_3_pipe71), .B(_12842_), .Y(_8777_) );
DFFPOSX1 DFFPOSX1_1177 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_8703__0_), .Q(H_3_0_) );
DFFPOSX1 DFFPOSX1_1178 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_8703__1_), .Q(H_3_1_) );
DFFPOSX1 DFFPOSX1_1179 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_8703__2_), .Q(H_3_2_) );
DFFPOSX1 DFFPOSX1_1180 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_8703__3_), .Q(H_3_3_) );
DFFPOSX1 DFFPOSX1_1181 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_8703__4_), .Q(H_3_4_) );
DFFPOSX1 DFFPOSX1_1182 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_8703__5_), .Q(H_3_5_) );
DFFPOSX1 DFFPOSX1_1183 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_8703__6_), .Q(H_3_6_) );
DFFPOSX1 DFFPOSX1_1184 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_8703__7_), .Q(H_3_7_) );
DFFPOSX1 DFFPOSX1_1185 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_8703__8_), .Q(H_3_8_) );
DFFPOSX1 DFFPOSX1_1186 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_8703__9_), .Q(H_3_9_) );
DFFPOSX1 DFFPOSX1_1187 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_8703__10_), .Q(H_3_10_) );
DFFPOSX1 DFFPOSX1_1188 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_8703__11_), .Q(H_3_11_) );
DFFPOSX1 DFFPOSX1_1189 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_8703__12_), .Q(H_3_12_) );
DFFPOSX1 DFFPOSX1_1190 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_8703__13_), .Q(H_3_13_) );
DFFPOSX1 DFFPOSX1_1191 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_8703__14_), .Q(H_3_14_) );
DFFPOSX1 DFFPOSX1_1192 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_8703__15_), .Q(H_3_15_) );
DFFPOSX1 DFFPOSX1_1193 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_8703__16_), .Q(H_3_16_) );
DFFPOSX1 DFFPOSX1_1194 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_8703__17_), .Q(H_3_17_) );
DFFPOSX1 DFFPOSX1_1195 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_8703__18_), .Q(H_3_18_) );
DFFPOSX1 DFFPOSX1_1196 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_8703__19_), .Q(H_3_19_) );
DFFPOSX1 DFFPOSX1_1197 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_8703__20_), .Q(H_3_20_) );
DFFPOSX1 DFFPOSX1_1198 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_8703__21_), .Q(H_3_21_) );
DFFPOSX1 DFFPOSX1_1199 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_8703__22_), .Q(H_3_22_) );
DFFPOSX1 DFFPOSX1_1200 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_8703__23_), .Q(H_3_23_) );
DFFPOSX1 DFFPOSX1_1201 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_8777_), .Q(comparador_3_valid_hash) );
DFFPOSX1 DFFPOSX1_1202 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_8701__0_), .Q(micro_hash_ucr_3_b_0_) );
DFFPOSX1 DFFPOSX1_1203 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_8701__1_), .Q(micro_hash_ucr_3_b_1_) );
DFFPOSX1 DFFPOSX1_1204 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_8701__2_), .Q(micro_hash_ucr_3_b_2_) );
DFFPOSX1 DFFPOSX1_1205 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_8701__3_), .Q(micro_hash_ucr_3_b_3_) );
DFFPOSX1 DFFPOSX1_1206 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_8701__4_), .Q(micro_hash_ucr_3_b_4_) );
DFFPOSX1 DFFPOSX1_1207 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_8701__5_), .Q(micro_hash_ucr_3_b_5_) );
DFFPOSX1 DFFPOSX1_1208 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_8701__6_), .Q(micro_hash_ucr_3_b_6_) );
DFFPOSX1 DFFPOSX1_1209 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_8701__7_), .Q(micro_hash_ucr_3_b_7_) );
DFFPOSX1 DFFPOSX1_1210 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_8702__0_), .Q(micro_hash_ucr_3_c_0_) );
DFFPOSX1 DFFPOSX1_1211 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_8702__1_), .Q(micro_hash_ucr_3_c_1_) );
DFFPOSX1 DFFPOSX1_1212 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_8702__2_), .Q(micro_hash_ucr_3_c_2_) );
DFFPOSX1 DFFPOSX1_1213 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_8702__3_), .Q(micro_hash_ucr_3_c_3_) );
DFFPOSX1 DFFPOSX1_1214 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_8702__4_), .Q(micro_hash_ucr_3_c_4_) );
DFFPOSX1 DFFPOSX1_1215 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_8702__5_), .Q(micro_hash_ucr_3_c_5_) );
DFFPOSX1 DFFPOSX1_1216 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_8702__6_), .Q(micro_hash_ucr_3_c_6_) );
DFFPOSX1 DFFPOSX1_1217 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_8702__7_), .Q(micro_hash_ucr_3_c_7_) );
DFFPOSX1 DFFPOSX1_1218 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_8778__0_), .Q(micro_hash_ucr_3_x_0_) );
DFFPOSX1 DFFPOSX1_1219 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_8778__1_), .Q(micro_hash_ucr_3_x_1_) );
DFFPOSX1 DFFPOSX1_1220 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_8778__2_), .Q(micro_hash_ucr_3_x_2_) );
DFFPOSX1 DFFPOSX1_1221 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_8778__3_), .Q(micro_hash_ucr_3_x_3_) );
DFFPOSX1 DFFPOSX1_1222 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_8778__4_), .Q(micro_hash_ucr_3_x_4_) );
DFFPOSX1 DFFPOSX1_1223 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_8778__5_), .Q(micro_hash_ucr_3_x_5_) );
DFFPOSX1 DFFPOSX1_1224 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_8778__6_), .Q(micro_hash_ucr_3_x_6_) );
DFFPOSX1 DFFPOSX1_1225 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_8778__7_), .Q(micro_hash_ucr_3_x_7_) );
DFFPOSX1 DFFPOSX1_1226 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_8704__0_), .Q(micro_hash_ucr_3_k_0_) );
DFFPOSX1 DFFPOSX1_1227 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_8704__1_), .Q(micro_hash_ucr_3_k_1_) );
DFFPOSX1 DFFPOSX1_1228 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_8704__2_), .Q(micro_hash_ucr_3_k_2_) );
DFFPOSX1 DFFPOSX1_1229 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_8704__3_), .Q(micro_hash_ucr_3_k_3_) );
DFFPOSX1 DFFPOSX1_1230 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_8704__4_), .Q(micro_hash_ucr_3_k_4_) );
DFFPOSX1 DFFPOSX1_1231 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_8704__5_), .Q(micro_hash_ucr_3_k_5_) );
DFFPOSX1 DFFPOSX1_1232 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_8704__6_), .Q(micro_hash_ucr_3_k_6_) );
DFFPOSX1 DFFPOSX1_1233 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_8704__7_), .Q(micro_hash_ucr_3_k_7_) );
DFFPOSX1 DFFPOSX1_1234 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_8700__0_), .Q(micro_hash_ucr_3_a_0_) );
DFFPOSX1 DFFPOSX1_1235 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_8700__1_), .Q(micro_hash_ucr_3_a_1_) );
DFFPOSX1 DFFPOSX1_1236 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_8700__2_), .Q(micro_hash_ucr_3_a_2_) );
DFFPOSX1 DFFPOSX1_1237 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_8700__3_), .Q(micro_hash_ucr_3_a_3_) );
DFFPOSX1 DFFPOSX1_1238 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_8700__4_), .Q(micro_hash_ucr_3_a_4_) );
DFFPOSX1 DFFPOSX1_1239 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_8700__5_), .Q(micro_hash_ucr_3_a_5_) );
DFFPOSX1 DFFPOSX1_1240 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_8700__6_), .Q(micro_hash_ucr_3_a_6_) );
DFFPOSX1 DFFPOSX1_1241 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_8700__7_), .Q(micro_hash_ucr_3_a_7_) );
DFFPOSX1 DFFPOSX1_1242 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_8705__bF_buf11), .Q(micro_hash_ucr_3_pipe0) );
DFFPOSX1 DFFPOSX1_1243 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_8699__0_), .Q(micro_hash_ucr_3_Wx_0_) );
DFFPOSX1 DFFPOSX1_1244 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_8699__1_), .Q(micro_hash_ucr_3_Wx_1_) );
DFFPOSX1 DFFPOSX1_1245 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_8699__2_), .Q(micro_hash_ucr_3_Wx_2_) );
DFFPOSX1 DFFPOSX1_1246 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_8699__3_), .Q(micro_hash_ucr_3_Wx_3_) );
DFFPOSX1 DFFPOSX1_1247 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_8699__4_), .Q(micro_hash_ucr_3_Wx_4_) );
DFFPOSX1 DFFPOSX1_1248 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_8699__5_), .Q(micro_hash_ucr_3_Wx_5_) );
DFFPOSX1 DFFPOSX1_1249 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_8699__6_), .Q(micro_hash_ucr_3_Wx_6_) );
DFFPOSX1 DFFPOSX1_1250 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_8699__7_), .Q(micro_hash_ucr_3_Wx_7_) );
DFFPOSX1 DFFPOSX1_1251 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_8699__8_), .Q(micro_hash_ucr_3_Wx_8_) );
DFFPOSX1 DFFPOSX1_1252 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_8699__9_), .Q(micro_hash_ucr_3_Wx_9_) );
DFFPOSX1 DFFPOSX1_1253 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_8699__10_), .Q(micro_hash_ucr_3_Wx_10_) );
DFFPOSX1 DFFPOSX1_1254 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_8699__11_), .Q(micro_hash_ucr_3_Wx_11_) );
DFFPOSX1 DFFPOSX1_1255 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_8699__12_), .Q(micro_hash_ucr_3_Wx_12_) );
DFFPOSX1 DFFPOSX1_1256 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_8699__13_), .Q(micro_hash_ucr_3_Wx_13_) );
DFFPOSX1 DFFPOSX1_1257 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_8699__14_), .Q(micro_hash_ucr_3_Wx_14_) );
DFFPOSX1 DFFPOSX1_1258 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_8699__15_), .Q(micro_hash_ucr_3_Wx_15_) );
DFFPOSX1 DFFPOSX1_1259 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_8699__16_), .Q(micro_hash_ucr_3_Wx_16_) );
DFFPOSX1 DFFPOSX1_1260 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_8699__17_), .Q(micro_hash_ucr_3_Wx_17_) );
DFFPOSX1 DFFPOSX1_1261 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_8699__18_), .Q(micro_hash_ucr_3_Wx_18_) );
DFFPOSX1 DFFPOSX1_1262 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_8699__19_), .Q(micro_hash_ucr_3_Wx_19_) );
DFFPOSX1 DFFPOSX1_1263 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_8699__20_), .Q(micro_hash_ucr_3_Wx_20_) );
DFFPOSX1 DFFPOSX1_1264 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_8699__21_), .Q(micro_hash_ucr_3_Wx_21_) );
DFFPOSX1 DFFPOSX1_1265 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf157), .D(_8699__22_), .Q(micro_hash_ucr_3_Wx_22_) );
DFFPOSX1 DFFPOSX1_1266 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf156), .D(_8699__23_), .Q(micro_hash_ucr_3_Wx_23_) );
DFFPOSX1 DFFPOSX1_1267 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf155), .D(_8699__24_), .Q(micro_hash_ucr_3_Wx_24_) );
DFFPOSX1 DFFPOSX1_1268 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf154), .D(_8699__25_), .Q(micro_hash_ucr_3_Wx_25_) );
DFFPOSX1 DFFPOSX1_1269 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf153), .D(_8699__26_), .Q(micro_hash_ucr_3_Wx_26_) );
DFFPOSX1 DFFPOSX1_1270 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf152), .D(_8699__27_), .Q(micro_hash_ucr_3_Wx_27_) );
DFFPOSX1 DFFPOSX1_1271 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf151), .D(_8699__28_), .Q(micro_hash_ucr_3_Wx_28_) );
DFFPOSX1 DFFPOSX1_1272 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf150), .D(_8699__29_), .Q(micro_hash_ucr_3_Wx_29_) );
DFFPOSX1 DFFPOSX1_1273 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf149), .D(_8699__30_), .Q(micro_hash_ucr_3_Wx_30_) );
DFFPOSX1 DFFPOSX1_1274 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf148), .D(_8699__31_), .Q(micro_hash_ucr_3_Wx_31_) );
DFFPOSX1 DFFPOSX1_1275 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf147), .D(_8699__32_), .Q(micro_hash_ucr_3_Wx_32_) );
DFFPOSX1 DFFPOSX1_1276 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf146), .D(_8699__33_), .Q(micro_hash_ucr_3_Wx_33_) );
DFFPOSX1 DFFPOSX1_1277 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf145), .D(_8699__34_), .Q(micro_hash_ucr_3_Wx_34_) );
DFFPOSX1 DFFPOSX1_1278 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf144), .D(_8699__35_), .Q(micro_hash_ucr_3_Wx_35_) );
DFFPOSX1 DFFPOSX1_1279 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf143), .D(_8699__36_), .Q(micro_hash_ucr_3_Wx_36_) );
DFFPOSX1 DFFPOSX1_1280 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf142), .D(_8699__37_), .Q(micro_hash_ucr_3_Wx_37_) );
DFFPOSX1 DFFPOSX1_1281 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf141), .D(_8699__38_), .Q(micro_hash_ucr_3_Wx_38_) );
DFFPOSX1 DFFPOSX1_1282 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf140), .D(_8699__39_), .Q(micro_hash_ucr_3_Wx_39_) );
DFFPOSX1 DFFPOSX1_1283 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf139), .D(_8699__40_), .Q(micro_hash_ucr_3_Wx_40_) );
DFFPOSX1 DFFPOSX1_1284 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf138), .D(_8699__41_), .Q(micro_hash_ucr_3_Wx_41_) );
DFFPOSX1 DFFPOSX1_1285 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf137), .D(_8699__42_), .Q(micro_hash_ucr_3_Wx_42_) );
DFFPOSX1 DFFPOSX1_1286 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf136), .D(_8699__43_), .Q(micro_hash_ucr_3_Wx_43_) );
DFFPOSX1 DFFPOSX1_1287 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf135), .D(_8699__44_), .Q(micro_hash_ucr_3_Wx_44_) );
DFFPOSX1 DFFPOSX1_1288 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf134), .D(_8699__45_), .Q(micro_hash_ucr_3_Wx_45_) );
DFFPOSX1 DFFPOSX1_1289 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf133), .D(_8699__46_), .Q(micro_hash_ucr_3_Wx_46_) );
DFFPOSX1 DFFPOSX1_1290 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf132), .D(_8699__47_), .Q(micro_hash_ucr_3_Wx_47_) );
DFFPOSX1 DFFPOSX1_1291 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf131), .D(_8699__48_), .Q(micro_hash_ucr_3_Wx_48_) );
DFFPOSX1 DFFPOSX1_1292 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf130), .D(_8699__49_), .Q(micro_hash_ucr_3_Wx_49_) );
DFFPOSX1 DFFPOSX1_1293 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf129), .D(_8699__50_), .Q(micro_hash_ucr_3_Wx_50_) );
DFFPOSX1 DFFPOSX1_1294 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf128), .D(_8699__51_), .Q(micro_hash_ucr_3_Wx_51_) );
DFFPOSX1 DFFPOSX1_1295 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf127), .D(_8699__52_), .Q(micro_hash_ucr_3_Wx_52_) );
DFFPOSX1 DFFPOSX1_1296 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf126), .D(_8699__53_), .Q(micro_hash_ucr_3_Wx_53_) );
DFFPOSX1 DFFPOSX1_1297 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf125), .D(_8699__54_), .Q(micro_hash_ucr_3_Wx_54_) );
DFFPOSX1 DFFPOSX1_1298 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf124), .D(_8699__55_), .Q(micro_hash_ucr_3_Wx_55_) );
DFFPOSX1 DFFPOSX1_1299 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf123), .D(_8699__56_), .Q(micro_hash_ucr_3_Wx_56_) );
DFFPOSX1 DFFPOSX1_1300 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf122), .D(_8699__57_), .Q(micro_hash_ucr_3_Wx_57_) );
DFFPOSX1 DFFPOSX1_1301 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf121), .D(_8699__58_), .Q(micro_hash_ucr_3_Wx_58_) );
DFFPOSX1 DFFPOSX1_1302 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf120), .D(_8699__59_), .Q(micro_hash_ucr_3_Wx_59_) );
DFFPOSX1 DFFPOSX1_1303 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf119), .D(_8699__60_), .Q(micro_hash_ucr_3_Wx_60_) );
DFFPOSX1 DFFPOSX1_1304 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf118), .D(_8699__61_), .Q(micro_hash_ucr_3_Wx_61_) );
DFFPOSX1 DFFPOSX1_1305 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf117), .D(_8699__62_), .Q(micro_hash_ucr_3_Wx_62_) );
DFFPOSX1 DFFPOSX1_1306 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf116), .D(_8699__63_), .Q(micro_hash_ucr_3_Wx_63_) );
DFFPOSX1 DFFPOSX1_1307 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf115), .D(_8699__64_), .Q(micro_hash_ucr_3_Wx_64_) );
DFFPOSX1 DFFPOSX1_1308 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf114), .D(_8699__65_), .Q(micro_hash_ucr_3_Wx_65_) );
DFFPOSX1 DFFPOSX1_1309 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf113), .D(_8699__66_), .Q(micro_hash_ucr_3_Wx_66_) );
DFFPOSX1 DFFPOSX1_1310 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf112), .D(_8699__67_), .Q(micro_hash_ucr_3_Wx_67_) );
DFFPOSX1 DFFPOSX1_1311 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf111), .D(_8699__68_), .Q(micro_hash_ucr_3_Wx_68_) );
DFFPOSX1 DFFPOSX1_1312 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf110), .D(_8699__69_), .Q(micro_hash_ucr_3_Wx_69_) );
DFFPOSX1 DFFPOSX1_1313 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf109), .D(_8699__70_), .Q(micro_hash_ucr_3_Wx_70_) );
DFFPOSX1 DFFPOSX1_1314 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf108), .D(_8699__71_), .Q(micro_hash_ucr_3_Wx_71_) );
DFFPOSX1 DFFPOSX1_1315 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf107), .D(_8699__72_), .Q(micro_hash_ucr_3_Wx_72_) );
DFFPOSX1 DFFPOSX1_1316 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(_8699__73_), .Q(micro_hash_ucr_3_Wx_73_) );
DFFPOSX1 DFFPOSX1_1317 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(_8699__74_), .Q(micro_hash_ucr_3_Wx_74_) );
DFFPOSX1 DFFPOSX1_1318 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(_8699__75_), .Q(micro_hash_ucr_3_Wx_75_) );
DFFPOSX1 DFFPOSX1_1319 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(_8699__76_), .Q(micro_hash_ucr_3_Wx_76_) );
DFFPOSX1 DFFPOSX1_1320 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(_8699__77_), .Q(micro_hash_ucr_3_Wx_77_) );
DFFPOSX1 DFFPOSX1_1321 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(_8699__78_), .Q(micro_hash_ucr_3_Wx_78_) );
DFFPOSX1 DFFPOSX1_1322 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(_8699__79_), .Q(micro_hash_ucr_3_Wx_79_) );
DFFPOSX1 DFFPOSX1_1323 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(_8699__80_), .Q(micro_hash_ucr_3_Wx_80_) );
DFFPOSX1 DFFPOSX1_1324 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_8699__81_), .Q(micro_hash_ucr_3_Wx_81_) );
DFFPOSX1 DFFPOSX1_1325 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_8699__82_), .Q(micro_hash_ucr_3_Wx_82_) );
DFFPOSX1 DFFPOSX1_1326 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_8699__83_), .Q(micro_hash_ucr_3_Wx_83_) );
DFFPOSX1 DFFPOSX1_1327 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_8699__84_), .Q(micro_hash_ucr_3_Wx_84_) );
DFFPOSX1 DFFPOSX1_1328 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_8699__85_), .Q(micro_hash_ucr_3_Wx_85_) );
DFFPOSX1 DFFPOSX1_1329 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_8699__86_), .Q(micro_hash_ucr_3_Wx_86_) );
DFFPOSX1 DFFPOSX1_1330 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_8699__87_), .Q(micro_hash_ucr_3_Wx_87_) );
DFFPOSX1 DFFPOSX1_1331 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_8699__88_), .Q(micro_hash_ucr_3_Wx_88_) );
DFFPOSX1 DFFPOSX1_1332 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_8699__89_), .Q(micro_hash_ucr_3_Wx_89_) );
DFFPOSX1 DFFPOSX1_1333 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_8699__90_), .Q(micro_hash_ucr_3_Wx_90_) );
DFFPOSX1 DFFPOSX1_1334 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_8699__91_), .Q(micro_hash_ucr_3_Wx_91_) );
DFFPOSX1 DFFPOSX1_1335 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_8699__92_), .Q(micro_hash_ucr_3_Wx_92_) );
DFFPOSX1 DFFPOSX1_1336 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_8699__93_), .Q(micro_hash_ucr_3_Wx_93_) );
DFFPOSX1 DFFPOSX1_1337 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_8699__94_), .Q(micro_hash_ucr_3_Wx_94_) );
DFFPOSX1 DFFPOSX1_1338 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_8699__95_), .Q(micro_hash_ucr_3_Wx_95_) );
DFFPOSX1 DFFPOSX1_1339 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_8699__96_), .Q(micro_hash_ucr_3_Wx_96_) );
DFFPOSX1 DFFPOSX1_1340 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_8699__97_), .Q(micro_hash_ucr_3_Wx_97_) );
DFFPOSX1 DFFPOSX1_1341 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_8699__98_), .Q(micro_hash_ucr_3_Wx_98_) );
DFFPOSX1 DFFPOSX1_1342 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_8699__99_), .Q(micro_hash_ucr_3_Wx_99_) );
DFFPOSX1 DFFPOSX1_1343 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_8699__100_), .Q(micro_hash_ucr_3_Wx_100_) );
DFFPOSX1 DFFPOSX1_1344 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_8699__101_), .Q(micro_hash_ucr_3_Wx_101_) );
DFFPOSX1 DFFPOSX1_1345 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_8699__102_), .Q(micro_hash_ucr_3_Wx_102_) );
DFFPOSX1 DFFPOSX1_1346 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_8699__103_), .Q(micro_hash_ucr_3_Wx_103_) );
DFFPOSX1 DFFPOSX1_1347 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_8699__104_), .Q(micro_hash_ucr_3_Wx_104_) );
DFFPOSX1 DFFPOSX1_1348 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_8699__105_), .Q(micro_hash_ucr_3_Wx_105_) );
DFFPOSX1 DFFPOSX1_1349 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_8699__106_), .Q(micro_hash_ucr_3_Wx_106_) );
DFFPOSX1 DFFPOSX1_1350 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_8699__107_), .Q(micro_hash_ucr_3_Wx_107_) );
DFFPOSX1 DFFPOSX1_1351 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_8699__108_), .Q(micro_hash_ucr_3_Wx_108_) );
DFFPOSX1 DFFPOSX1_1352 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_8699__109_), .Q(micro_hash_ucr_3_Wx_109_) );
DFFPOSX1 DFFPOSX1_1353 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_8699__110_), .Q(micro_hash_ucr_3_Wx_110_) );
DFFPOSX1 DFFPOSX1_1354 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_8699__111_), .Q(micro_hash_ucr_3_Wx_111_) );
DFFPOSX1 DFFPOSX1_1355 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_8699__112_), .Q(micro_hash_ucr_3_Wx_112_) );
DFFPOSX1 DFFPOSX1_1356 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_8699__113_), .Q(micro_hash_ucr_3_Wx_113_) );
DFFPOSX1 DFFPOSX1_1357 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_8699__114_), .Q(micro_hash_ucr_3_Wx_114_) );
DFFPOSX1 DFFPOSX1_1358 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_8699__115_), .Q(micro_hash_ucr_3_Wx_115_) );
DFFPOSX1 DFFPOSX1_1359 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_8699__116_), .Q(micro_hash_ucr_3_Wx_116_) );
DFFPOSX1 DFFPOSX1_1360 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_8699__117_), .Q(micro_hash_ucr_3_Wx_117_) );
DFFPOSX1 DFFPOSX1_1361 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_8699__118_), .Q(micro_hash_ucr_3_Wx_118_) );
DFFPOSX1 DFFPOSX1_1362 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_8699__119_), .Q(micro_hash_ucr_3_Wx_119_) );
DFFPOSX1 DFFPOSX1_1363 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_8699__120_), .Q(micro_hash_ucr_3_Wx_120_) );
DFFPOSX1 DFFPOSX1_1364 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_8699__121_), .Q(micro_hash_ucr_3_Wx_121_) );
DFFPOSX1 DFFPOSX1_1365 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_8699__122_), .Q(micro_hash_ucr_3_Wx_122_) );
DFFPOSX1 DFFPOSX1_1366 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_8699__123_), .Q(micro_hash_ucr_3_Wx_123_) );
DFFPOSX1 DFFPOSX1_1367 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_8699__124_), .Q(micro_hash_ucr_3_Wx_124_) );
DFFPOSX1 DFFPOSX1_1368 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_8699__125_), .Q(micro_hash_ucr_3_Wx_125_) );
DFFPOSX1 DFFPOSX1_1369 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_8699__126_), .Q(micro_hash_ucr_3_Wx_126_) );
DFFPOSX1 DFFPOSX1_1370 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_8699__127_), .Q(micro_hash_ucr_3_Wx_127_) );
DFFPOSX1 DFFPOSX1_1371 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_8699__128_), .Q(micro_hash_ucr_3_Wx_128_) );
DFFPOSX1 DFFPOSX1_1372 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_8699__129_), .Q(micro_hash_ucr_3_Wx_129_) );
DFFPOSX1 DFFPOSX1_1373 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_8699__130_), .Q(micro_hash_ucr_3_Wx_130_) );
DFFPOSX1 DFFPOSX1_1374 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_8699__131_), .Q(micro_hash_ucr_3_Wx_131_) );
DFFPOSX1 DFFPOSX1_1375 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_8699__132_), .Q(micro_hash_ucr_3_Wx_132_) );
DFFPOSX1 DFFPOSX1_1376 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_8699__133_), .Q(micro_hash_ucr_3_Wx_133_) );
DFFPOSX1 DFFPOSX1_1377 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_8699__134_), .Q(micro_hash_ucr_3_Wx_134_) );
DFFPOSX1 DFFPOSX1_1378 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_8699__135_), .Q(micro_hash_ucr_3_Wx_135_) );
DFFPOSX1 DFFPOSX1_1379 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_8699__136_), .Q(micro_hash_ucr_3_Wx_136_) );
DFFPOSX1 DFFPOSX1_1380 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_8699__137_), .Q(micro_hash_ucr_3_Wx_137_) );
DFFPOSX1 DFFPOSX1_1381 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_8699__138_), .Q(micro_hash_ucr_3_Wx_138_) );
DFFPOSX1 DFFPOSX1_1382 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_8699__139_), .Q(micro_hash_ucr_3_Wx_139_) );
DFFPOSX1 DFFPOSX1_1383 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_8699__140_), .Q(micro_hash_ucr_3_Wx_140_) );
DFFPOSX1 DFFPOSX1_1384 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_8699__141_), .Q(micro_hash_ucr_3_Wx_141_) );
DFFPOSX1 DFFPOSX1_1385 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_8699__142_), .Q(micro_hash_ucr_3_Wx_142_) );
DFFPOSX1 DFFPOSX1_1386 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_8699__143_), .Q(micro_hash_ucr_3_Wx_143_) );
DFFPOSX1 DFFPOSX1_1387 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_8699__144_), .Q(micro_hash_ucr_3_Wx_144_) );
DFFPOSX1 DFFPOSX1_1388 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_8699__145_), .Q(micro_hash_ucr_3_Wx_145_) );
DFFPOSX1 DFFPOSX1_1389 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_8699__146_), .Q(micro_hash_ucr_3_Wx_146_) );
DFFPOSX1 DFFPOSX1_1390 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_8699__147_), .Q(micro_hash_ucr_3_Wx_147_) );
DFFPOSX1 DFFPOSX1_1391 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_8699__148_), .Q(micro_hash_ucr_3_Wx_148_) );
DFFPOSX1 DFFPOSX1_1392 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_8699__149_), .Q(micro_hash_ucr_3_Wx_149_) );
DFFPOSX1 DFFPOSX1_1393 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_8699__150_), .Q(micro_hash_ucr_3_Wx_150_) );
DFFPOSX1 DFFPOSX1_1394 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_8699__151_), .Q(micro_hash_ucr_3_Wx_151_) );
DFFPOSX1 DFFPOSX1_1395 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_8699__152_), .Q(micro_hash_ucr_3_Wx_152_) );
DFFPOSX1 DFFPOSX1_1396 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_8699__153_), .Q(micro_hash_ucr_3_Wx_153_) );
DFFPOSX1 DFFPOSX1_1397 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_8699__154_), .Q(micro_hash_ucr_3_Wx_154_) );
DFFPOSX1 DFFPOSX1_1398 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_8699__155_), .Q(micro_hash_ucr_3_Wx_155_) );
DFFPOSX1 DFFPOSX1_1399 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_8699__156_), .Q(micro_hash_ucr_3_Wx_156_) );
DFFPOSX1 DFFPOSX1_1400 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_8699__157_), .Q(micro_hash_ucr_3_Wx_157_) );
DFFPOSX1 DFFPOSX1_1401 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_8699__158_), .Q(micro_hash_ucr_3_Wx_158_) );
DFFPOSX1 DFFPOSX1_1402 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_8699__159_), .Q(micro_hash_ucr_3_Wx_159_) );
DFFPOSX1 DFFPOSX1_1403 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_8699__160_), .Q(micro_hash_ucr_3_Wx_160_) );
DFFPOSX1 DFFPOSX1_1404 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_8699__161_), .Q(micro_hash_ucr_3_Wx_161_) );
DFFPOSX1 DFFPOSX1_1405 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_8699__162_), .Q(micro_hash_ucr_3_Wx_162_) );
DFFPOSX1 DFFPOSX1_1406 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_8699__163_), .Q(micro_hash_ucr_3_Wx_163_) );
DFFPOSX1 DFFPOSX1_1407 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_8699__164_), .Q(micro_hash_ucr_3_Wx_164_) );
DFFPOSX1 DFFPOSX1_1408 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_8699__165_), .Q(micro_hash_ucr_3_Wx_165_) );
DFFPOSX1 DFFPOSX1_1409 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_8699__166_), .Q(micro_hash_ucr_3_Wx_166_) );
DFFPOSX1 DFFPOSX1_1410 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_8699__167_), .Q(micro_hash_ucr_3_Wx_167_) );
DFFPOSX1 DFFPOSX1_1411 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_8699__168_), .Q(micro_hash_ucr_3_Wx_168_) );
DFFPOSX1 DFFPOSX1_1412 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_8699__169_), .Q(micro_hash_ucr_3_Wx_169_) );
DFFPOSX1 DFFPOSX1_1413 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_8699__170_), .Q(micro_hash_ucr_3_Wx_170_) );
DFFPOSX1 DFFPOSX1_1414 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_8699__171_), .Q(micro_hash_ucr_3_Wx_171_) );
DFFPOSX1 DFFPOSX1_1415 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_8699__172_), .Q(micro_hash_ucr_3_Wx_172_) );
DFFPOSX1 DFFPOSX1_1416 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_8699__173_), .Q(micro_hash_ucr_3_Wx_173_) );
DFFPOSX1 DFFPOSX1_1417 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_8699__174_), .Q(micro_hash_ucr_3_Wx_174_) );
DFFPOSX1 DFFPOSX1_1418 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_8699__175_), .Q(micro_hash_ucr_3_Wx_175_) );
DFFPOSX1 DFFPOSX1_1419 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_8699__176_), .Q(micro_hash_ucr_3_Wx_176_) );
DFFPOSX1 DFFPOSX1_1420 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_8699__177_), .Q(micro_hash_ucr_3_Wx_177_) );
DFFPOSX1 DFFPOSX1_1421 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_8699__178_), .Q(micro_hash_ucr_3_Wx_178_) );
DFFPOSX1 DFFPOSX1_1422 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_8699__179_), .Q(micro_hash_ucr_3_Wx_179_) );
DFFPOSX1 DFFPOSX1_1423 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf157), .D(_8699__180_), .Q(micro_hash_ucr_3_Wx_180_) );
DFFPOSX1 DFFPOSX1_1424 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf156), .D(_8699__181_), .Q(micro_hash_ucr_3_Wx_181_) );
DFFPOSX1 DFFPOSX1_1425 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf155), .D(_8699__182_), .Q(micro_hash_ucr_3_Wx_182_) );
DFFPOSX1 DFFPOSX1_1426 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf154), .D(_8699__183_), .Q(micro_hash_ucr_3_Wx_183_) );
DFFPOSX1 DFFPOSX1_1427 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf153), .D(_8699__184_), .Q(micro_hash_ucr_3_Wx_184_) );
DFFPOSX1 DFFPOSX1_1428 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf152), .D(_8699__185_), .Q(micro_hash_ucr_3_Wx_185_) );
DFFPOSX1 DFFPOSX1_1429 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf151), .D(_8699__186_), .Q(micro_hash_ucr_3_Wx_186_) );
DFFPOSX1 DFFPOSX1_1430 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf150), .D(_8699__187_), .Q(micro_hash_ucr_3_Wx_187_) );
DFFPOSX1 DFFPOSX1_1431 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf149), .D(_8699__188_), .Q(micro_hash_ucr_3_Wx_188_) );
DFFPOSX1 DFFPOSX1_1432 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf148), .D(_8699__189_), .Q(micro_hash_ucr_3_Wx_189_) );
DFFPOSX1 DFFPOSX1_1433 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf147), .D(_8699__190_), .Q(micro_hash_ucr_3_Wx_190_) );
DFFPOSX1 DFFPOSX1_1434 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf146), .D(_8699__191_), .Q(micro_hash_ucr_3_Wx_191_) );
DFFPOSX1 DFFPOSX1_1435 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf145), .D(_8699__192_), .Q(micro_hash_ucr_3_Wx_192_) );
DFFPOSX1 DFFPOSX1_1436 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf144), .D(_8699__193_), .Q(micro_hash_ucr_3_Wx_193_) );
DFFPOSX1 DFFPOSX1_1437 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf143), .D(_8699__194_), .Q(micro_hash_ucr_3_Wx_194_) );
DFFPOSX1 DFFPOSX1_1438 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf142), .D(_8699__195_), .Q(micro_hash_ucr_3_Wx_195_) );
DFFPOSX1 DFFPOSX1_1439 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf141), .D(_8699__196_), .Q(micro_hash_ucr_3_Wx_196_) );
DFFPOSX1 DFFPOSX1_1440 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf140), .D(_8699__197_), .Q(micro_hash_ucr_3_Wx_197_) );
DFFPOSX1 DFFPOSX1_1441 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf139), .D(_8699__198_), .Q(micro_hash_ucr_3_Wx_198_) );
DFFPOSX1 DFFPOSX1_1442 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf138), .D(_8699__199_), .Q(micro_hash_ucr_3_Wx_199_) );
DFFPOSX1 DFFPOSX1_1443 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf137), .D(_8699__200_), .Q(micro_hash_ucr_3_Wx_200_) );
DFFPOSX1 DFFPOSX1_1444 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf136), .D(_8699__201_), .Q(micro_hash_ucr_3_Wx_201_) );
DFFPOSX1 DFFPOSX1_1445 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf135), .D(_8699__202_), .Q(micro_hash_ucr_3_Wx_202_) );
DFFPOSX1 DFFPOSX1_1446 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf134), .D(_8699__203_), .Q(micro_hash_ucr_3_Wx_203_) );
DFFPOSX1 DFFPOSX1_1447 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf133), .D(_8699__204_), .Q(micro_hash_ucr_3_Wx_204_) );
DFFPOSX1 DFFPOSX1_1448 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf132), .D(_8699__205_), .Q(micro_hash_ucr_3_Wx_205_) );
DFFPOSX1 DFFPOSX1_1449 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf131), .D(_8699__206_), .Q(micro_hash_ucr_3_Wx_206_) );
DFFPOSX1 DFFPOSX1_1450 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf130), .D(_8699__207_), .Q(micro_hash_ucr_3_Wx_207_) );
DFFPOSX1 DFFPOSX1_1451 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf129), .D(_8699__208_), .Q(micro_hash_ucr_3_Wx_208_) );
DFFPOSX1 DFFPOSX1_1452 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf128), .D(_8699__209_), .Q(micro_hash_ucr_3_Wx_209_) );
DFFPOSX1 DFFPOSX1_1453 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf127), .D(_8699__210_), .Q(micro_hash_ucr_3_Wx_210_) );
DFFPOSX1 DFFPOSX1_1454 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf126), .D(_8699__211_), .Q(micro_hash_ucr_3_Wx_211_) );
DFFPOSX1 DFFPOSX1_1455 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf125), .D(_8699__212_), .Q(micro_hash_ucr_3_Wx_212_) );
DFFPOSX1 DFFPOSX1_1456 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf124), .D(_8699__213_), .Q(micro_hash_ucr_3_Wx_213_) );
DFFPOSX1 DFFPOSX1_1457 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf123), .D(_8699__214_), .Q(micro_hash_ucr_3_Wx_214_) );
DFFPOSX1 DFFPOSX1_1458 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf122), .D(_8699__215_), .Q(micro_hash_ucr_3_Wx_215_) );
DFFPOSX1 DFFPOSX1_1459 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf121), .D(_8699__216_), .Q(micro_hash_ucr_3_Wx_216_) );
DFFPOSX1 DFFPOSX1_1460 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf120), .D(_8699__217_), .Q(micro_hash_ucr_3_Wx_217_) );
DFFPOSX1 DFFPOSX1_1461 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf119), .D(_8699__218_), .Q(micro_hash_ucr_3_Wx_218_) );
DFFPOSX1 DFFPOSX1_1462 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf118), .D(_8699__219_), .Q(micro_hash_ucr_3_Wx_219_) );
DFFPOSX1 DFFPOSX1_1463 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf117), .D(_8699__220_), .Q(micro_hash_ucr_3_Wx_220_) );
DFFPOSX1 DFFPOSX1_1464 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf116), .D(_8699__221_), .Q(micro_hash_ucr_3_Wx_221_) );
DFFPOSX1 DFFPOSX1_1465 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf115), .D(_8699__222_), .Q(micro_hash_ucr_3_Wx_222_) );
DFFPOSX1 DFFPOSX1_1466 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf114), .D(_8699__223_), .Q(micro_hash_ucr_3_Wx_223_) );
DFFPOSX1 DFFPOSX1_1467 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf113), .D(_8699__224_), .Q(micro_hash_ucr_3_Wx_224_) );
DFFPOSX1 DFFPOSX1_1468 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf112), .D(_8699__225_), .Q(micro_hash_ucr_3_Wx_225_) );
DFFPOSX1 DFFPOSX1_1469 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf111), .D(_8699__226_), .Q(micro_hash_ucr_3_Wx_226_) );
DFFPOSX1 DFFPOSX1_1470 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf110), .D(_8699__227_), .Q(micro_hash_ucr_3_Wx_227_) );
DFFPOSX1 DFFPOSX1_1471 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf109), .D(_8699__228_), .Q(micro_hash_ucr_3_Wx_228_) );
DFFPOSX1 DFFPOSX1_1472 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf108), .D(_8699__229_), .Q(micro_hash_ucr_3_Wx_229_) );
DFFPOSX1 DFFPOSX1_1473 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf107), .D(_8699__230_), .Q(micro_hash_ucr_3_Wx_230_) );
DFFPOSX1 DFFPOSX1_1474 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(_8699__231_), .Q(micro_hash_ucr_3_Wx_231_) );
DFFPOSX1 DFFPOSX1_1475 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(_8699__232_), .Q(micro_hash_ucr_3_Wx_232_) );
DFFPOSX1 DFFPOSX1_1476 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(_8699__233_), .Q(micro_hash_ucr_3_Wx_233_) );
DFFPOSX1 DFFPOSX1_1477 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(_8699__234_), .Q(micro_hash_ucr_3_Wx_234_) );
DFFPOSX1 DFFPOSX1_1478 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(_8699__235_), .Q(micro_hash_ucr_3_Wx_235_) );
DFFPOSX1 DFFPOSX1_1479 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(_8699__236_), .Q(micro_hash_ucr_3_Wx_236_) );
DFFPOSX1 DFFPOSX1_1480 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(_8699__237_), .Q(micro_hash_ucr_3_Wx_237_) );
DFFPOSX1 DFFPOSX1_1481 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(_8699__238_), .Q(micro_hash_ucr_3_Wx_238_) );
DFFPOSX1 DFFPOSX1_1482 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_8699__239_), .Q(micro_hash_ucr_3_Wx_239_) );
DFFPOSX1 DFFPOSX1_1483 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_8699__240_), .Q(micro_hash_ucr_3_Wx_240_) );
DFFPOSX1 DFFPOSX1_1484 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_8699__241_), .Q(micro_hash_ucr_3_Wx_241_) );
DFFPOSX1 DFFPOSX1_1485 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_8699__242_), .Q(micro_hash_ucr_3_Wx_242_) );
DFFPOSX1 DFFPOSX1_1486 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_8699__243_), .Q(micro_hash_ucr_3_Wx_243_) );
DFFPOSX1 DFFPOSX1_1487 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_8699__244_), .Q(micro_hash_ucr_3_Wx_244_) );
DFFPOSX1 DFFPOSX1_1488 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_8699__245_), .Q(micro_hash_ucr_3_Wx_245_) );
DFFPOSX1 DFFPOSX1_1489 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_8699__246_), .Q(micro_hash_ucr_3_Wx_246_) );
DFFPOSX1 DFFPOSX1_1490 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_8699__247_), .Q(micro_hash_ucr_3_Wx_247_) );
DFFPOSX1 DFFPOSX1_1491 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_8699__248_), .Q(micro_hash_ucr_3_Wx_248_) );
DFFPOSX1 DFFPOSX1_1492 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_8699__249_), .Q(micro_hash_ucr_3_Wx_249_) );
DFFPOSX1 DFFPOSX1_1493 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_8699__250_), .Q(micro_hash_ucr_3_Wx_250_) );
DFFPOSX1 DFFPOSX1_1494 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_8699__251_), .Q(micro_hash_ucr_3_Wx_251_) );
DFFPOSX1 DFFPOSX1_1495 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_8699__252_), .Q(micro_hash_ucr_3_Wx_252_) );
DFFPOSX1 DFFPOSX1_1496 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_8699__253_), .Q(micro_hash_ucr_3_Wx_253_) );
DFFPOSX1 DFFPOSX1_1497 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_8699__254_), .Q(micro_hash_ucr_3_Wx_254_) );
DFFPOSX1 DFFPOSX1_1498 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_8699__255_), .Q(micro_hash_ucr_3_Wx_255_) );
DFFPOSX1 DFFPOSX1_1499 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_8716_), .Q(micro_hash_ucr_3_pipe1) );
DFFPOSX1 DFFPOSX1_1500 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_8727_), .Q(micro_hash_ucr_3_pipe2) );
DFFPOSX1 DFFPOSX1_1501 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_8738_), .Q(micro_hash_ucr_3_pipe3) );
DFFPOSX1 DFFPOSX1_1502 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_8749_), .Q(micro_hash_ucr_3_pipe4) );
DFFPOSX1 DFFPOSX1_1503 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_8760_), .Q(micro_hash_ucr_3_pipe5) );
DFFPOSX1 DFFPOSX1_1504 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_8771_), .Q(micro_hash_ucr_3_pipe6) );
DFFPOSX1 DFFPOSX1_1505 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_8774_), .Q(micro_hash_ucr_3_pipe7) );
DFFPOSX1 DFFPOSX1_1506 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_8775_), .Q(micro_hash_ucr_3_pipe8) );
DFFPOSX1 DFFPOSX1_1507 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_8776_), .Q(micro_hash_ucr_3_pipe9) );
DFFPOSX1 DFFPOSX1_1508 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_8706_), .Q(micro_hash_ucr_3_pipe10) );
DFFPOSX1 DFFPOSX1_1509 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_8707_), .Q(micro_hash_ucr_3_pipe11) );
DFFPOSX1 DFFPOSX1_1510 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_8708_), .Q(micro_hash_ucr_3_pipe12) );
DFFPOSX1 DFFPOSX1_1511 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_8709_), .Q(micro_hash_ucr_3_pipe13) );
DFFPOSX1 DFFPOSX1_1512 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_8710_), .Q(micro_hash_ucr_3_pipe14) );
DFFPOSX1 DFFPOSX1_1513 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_8711_), .Q(micro_hash_ucr_3_pipe15) );
DFFPOSX1 DFFPOSX1_1514 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_8712_), .Q(micro_hash_ucr_3_pipe16) );
DFFPOSX1 DFFPOSX1_1515 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_8713_), .Q(micro_hash_ucr_3_pipe17) );
DFFPOSX1 DFFPOSX1_1516 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_8714_), .Q(micro_hash_ucr_3_pipe18) );
DFFPOSX1 DFFPOSX1_1517 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_8715_), .Q(micro_hash_ucr_3_pipe19) );
DFFPOSX1 DFFPOSX1_1518 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_8717_), .Q(micro_hash_ucr_3_pipe20) );
DFFPOSX1 DFFPOSX1_1519 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_8718_), .Q(micro_hash_ucr_3_pipe21) );
DFFPOSX1 DFFPOSX1_1520 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_8719_), .Q(micro_hash_ucr_3_pipe22) );
DFFPOSX1 DFFPOSX1_1521 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_8720_), .Q(micro_hash_ucr_3_pipe23) );
DFFPOSX1 DFFPOSX1_1522 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_8721_), .Q(micro_hash_ucr_3_pipe24) );
DFFPOSX1 DFFPOSX1_1523 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_8722_), .Q(micro_hash_ucr_3_pipe25) );
DFFPOSX1 DFFPOSX1_1524 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_8723_), .Q(micro_hash_ucr_3_pipe26) );
DFFPOSX1 DFFPOSX1_1525 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_8724_), .Q(micro_hash_ucr_3_pipe27) );
DFFPOSX1 DFFPOSX1_1526 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_8725_), .Q(micro_hash_ucr_3_pipe28) );
DFFPOSX1 DFFPOSX1_1527 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_8726_), .Q(micro_hash_ucr_3_pipe29) );
DFFPOSX1 DFFPOSX1_1528 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_8728_), .Q(micro_hash_ucr_3_pipe30) );
DFFPOSX1 DFFPOSX1_1529 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_8729_), .Q(micro_hash_ucr_3_pipe31) );
DFFPOSX1 DFFPOSX1_1530 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_8730_), .Q(micro_hash_ucr_3_pipe32) );
DFFPOSX1 DFFPOSX1_1531 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_8731_), .Q(micro_hash_ucr_3_pipe33) );
DFFPOSX1 DFFPOSX1_1532 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_8732_), .Q(micro_hash_ucr_3_pipe34) );
DFFPOSX1 DFFPOSX1_1533 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_8733_), .Q(micro_hash_ucr_3_pipe35) );
DFFPOSX1 DFFPOSX1_1534 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_8734_), .Q(micro_hash_ucr_3_pipe36) );
DFFPOSX1 DFFPOSX1_1535 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_8735_), .Q(micro_hash_ucr_3_pipe37) );
DFFPOSX1 DFFPOSX1_1536 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_8736_), .Q(micro_hash_ucr_3_pipe38) );
DFFPOSX1 DFFPOSX1_1537 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_8737_), .Q(micro_hash_ucr_3_pipe39) );
DFFPOSX1 DFFPOSX1_1538 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_8739_), .Q(micro_hash_ucr_3_pipe40) );
DFFPOSX1 DFFPOSX1_1539 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_8740_), .Q(micro_hash_ucr_3_pipe41) );
DFFPOSX1 DFFPOSX1_1540 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_8741_), .Q(micro_hash_ucr_3_pipe42) );
DFFPOSX1 DFFPOSX1_1541 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_8742_), .Q(micro_hash_ucr_3_pipe43) );
DFFPOSX1 DFFPOSX1_1542 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_8743_), .Q(micro_hash_ucr_3_pipe44) );
DFFPOSX1 DFFPOSX1_1543 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_8744_), .Q(micro_hash_ucr_3_pipe45) );
DFFPOSX1 DFFPOSX1_1544 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_8745_), .Q(micro_hash_ucr_3_pipe46) );
DFFPOSX1 DFFPOSX1_1545 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_8746_), .Q(micro_hash_ucr_3_pipe47) );
DFFPOSX1 DFFPOSX1_1546 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_8747_), .Q(micro_hash_ucr_3_pipe48) );
DFFPOSX1 DFFPOSX1_1547 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_8748_), .Q(micro_hash_ucr_3_pipe49) );
DFFPOSX1 DFFPOSX1_1548 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_8750_), .Q(micro_hash_ucr_3_pipe50) );
DFFPOSX1 DFFPOSX1_1549 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_8751_), .Q(micro_hash_ucr_3_pipe51) );
DFFPOSX1 DFFPOSX1_1550 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_8752_), .Q(micro_hash_ucr_3_pipe52) );
DFFPOSX1 DFFPOSX1_1551 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_8753_), .Q(micro_hash_ucr_3_pipe53) );
DFFPOSX1 DFFPOSX1_1552 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_8754_), .Q(micro_hash_ucr_3_pipe54) );
DFFPOSX1 DFFPOSX1_1553 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_8755_), .Q(micro_hash_ucr_3_pipe55) );
DFFPOSX1 DFFPOSX1_1554 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_8756_), .Q(micro_hash_ucr_3_pipe56) );
DFFPOSX1 DFFPOSX1_1555 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_8757_), .Q(micro_hash_ucr_3_pipe57) );
DFFPOSX1 DFFPOSX1_1556 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_8758_), .Q(micro_hash_ucr_3_pipe58) );
DFFPOSX1 DFFPOSX1_1557 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_8759_), .Q(micro_hash_ucr_3_pipe59) );
DFFPOSX1 DFFPOSX1_1558 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_8761_), .Q(micro_hash_ucr_3_pipe60) );
DFFPOSX1 DFFPOSX1_1559 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_8762_), .Q(micro_hash_ucr_3_pipe61) );
DFFPOSX1 DFFPOSX1_1560 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_8763_), .Q(micro_hash_ucr_3_pipe62) );
DFFPOSX1 DFFPOSX1_1561 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_8764_), .Q(micro_hash_ucr_3_pipe63) );
DFFPOSX1 DFFPOSX1_1562 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_8765_), .Q(micro_hash_ucr_3_pipe64) );
DFFPOSX1 DFFPOSX1_1563 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_8766_), .Q(micro_hash_ucr_3_pipe65) );
DFFPOSX1 DFFPOSX1_1564 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_8767_), .Q(micro_hash_ucr_3_pipe66) );
DFFPOSX1 DFFPOSX1_1565 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_8768_), .Q(micro_hash_ucr_3_pipe67) );
DFFPOSX1 DFFPOSX1_1566 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_8769_), .Q(micro_hash_ucr_3_pipe68) );
DFFPOSX1 DFFPOSX1_1567 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_8770_), .Q(micro_hash_ucr_3_pipe69) );
DFFPOSX1 DFFPOSX1_1568 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_8772_), .Q(micro_hash_ucr_3_pipe70) );
DFFPOSX1 DFFPOSX1_1569 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_8773_), .Q(micro_hash_ucr_3_pipe71) );
INVX8 INVX8_287 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf4), .Y(_12916_) );
NAND2X1 NAND2X1_1697 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_0_), .B(_12916__bF_buf42), .Y(_12917_) );
MUX2X1 MUX2X1_37 ( .gnd(gnd), .vdd(vdd), .A(data_in[0]), .B(next_b_data_in_prev_0_), .S(_0__bF_buf5), .Y(_12918_) );
OAI21X1 OAI21X1_3663 ( .gnd(gnd), .vdd(vdd), .A(_12918_), .B(_12916__bF_buf41), .C(_12917_), .Y(_12914__0_) );
NAND2X1 NAND2X1_1698 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_1_), .B(_12916__bF_buf40), .Y(_12919_) );
MUX2X1 MUX2X1_38 ( .gnd(gnd), .vdd(vdd), .A(data_in[1]), .B(next_b_data_in_prev_1_), .S(_0__bF_buf4), .Y(_12920_) );
OAI21X1 OAI21X1_3664 ( .gnd(gnd), .vdd(vdd), .A(_12920_), .B(_12916__bF_buf39), .C(_12919_), .Y(_12914__1_) );
NAND2X1 NAND2X1_1699 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_2_), .B(_12916__bF_buf38), .Y(_12921_) );
MUX2X1 MUX2X1_39 ( .gnd(gnd), .vdd(vdd), .A(data_in[2]), .B(next_b_data_in_prev_2_), .S(_0__bF_buf3), .Y(_12922_) );
OAI21X1 OAI21X1_3665 ( .gnd(gnd), .vdd(vdd), .A(_12922_), .B(_12916__bF_buf37), .C(_12921_), .Y(_12914__2_) );
NAND2X1 NAND2X1_1700 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_3_), .B(_12916__bF_buf36), .Y(_12923_) );
MUX2X1 MUX2X1_40 ( .gnd(gnd), .vdd(vdd), .A(data_in[3]), .B(next_b_data_in_prev_3_), .S(_0__bF_buf2), .Y(_12924_) );
OAI21X1 OAI21X1_3666 ( .gnd(gnd), .vdd(vdd), .A(_12924_), .B(_12916__bF_buf35), .C(_12923_), .Y(_12914__3_) );
NAND2X1 NAND2X1_1701 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_4_), .B(_12916__bF_buf34), .Y(_12925_) );
MUX2X1 MUX2X1_41 ( .gnd(gnd), .vdd(vdd), .A(data_in[4]), .B(next_b_data_in_prev_4_), .S(_0__bF_buf1), .Y(_12926_) );
OAI21X1 OAI21X1_3667 ( .gnd(gnd), .vdd(vdd), .A(_12926_), .B(_12916__bF_buf33), .C(_12925_), .Y(_12914__4_) );
NAND2X1 NAND2X1_1702 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_5_), .B(_12916__bF_buf32), .Y(_12927_) );
MUX2X1 MUX2X1_42 ( .gnd(gnd), .vdd(vdd), .A(data_in[5]), .B(next_b_data_in_prev_5_), .S(_0__bF_buf0), .Y(_12928_) );
OAI21X1 OAI21X1_3668 ( .gnd(gnd), .vdd(vdd), .A(_12928_), .B(_12916__bF_buf31), .C(_12927_), .Y(_12914__5_) );
NAND2X1 NAND2X1_1703 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_6_), .B(_12916__bF_buf30), .Y(_12929_) );
MUX2X1 MUX2X1_43 ( .gnd(gnd), .vdd(vdd), .A(data_in[6]), .B(next_b_data_in_prev_6_), .S(_0__bF_buf9), .Y(_12930_) );
OAI21X1 OAI21X1_3669 ( .gnd(gnd), .vdd(vdd), .A(_12930_), .B(_12916__bF_buf29), .C(_12929_), .Y(_12914__6_) );
NAND2X1 NAND2X1_1704 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_7_), .B(_12916__bF_buf28), .Y(_12931_) );
MUX2X1 MUX2X1_44 ( .gnd(gnd), .vdd(vdd), .A(data_in[7]), .B(next_b_data_in_prev_7_), .S(_0__bF_buf8), .Y(_12932_) );
OAI21X1 OAI21X1_3670 ( .gnd(gnd), .vdd(vdd), .A(_12932_), .B(_12916__bF_buf27), .C(_12931_), .Y(_12914__7_) );
NAND2X1 NAND2X1_1705 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_8_), .B(_12916__bF_buf26), .Y(_12933_) );
MUX2X1 MUX2X1_45 ( .gnd(gnd), .vdd(vdd), .A(data_in[8]), .B(next_b_data_in_prev_8_), .S(_0__bF_buf7), .Y(_12934_) );
OAI21X1 OAI21X1_3671 ( .gnd(gnd), .vdd(vdd), .A(_12934_), .B(_12916__bF_buf25), .C(_12933_), .Y(_12914__8_) );
NAND2X1 NAND2X1_1706 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_9_), .B(_12916__bF_buf24), .Y(_12935_) );
MUX2X1 MUX2X1_46 ( .gnd(gnd), .vdd(vdd), .A(data_in[9]), .B(next_b_data_in_prev_9_), .S(_0__bF_buf6), .Y(_12936_) );
OAI21X1 OAI21X1_3672 ( .gnd(gnd), .vdd(vdd), .A(_12936_), .B(_12916__bF_buf23), .C(_12935_), .Y(_12914__9_) );
NAND2X1 NAND2X1_1707 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_10_), .B(_12916__bF_buf22), .Y(_12937_) );
MUX2X1 MUX2X1_47 ( .gnd(gnd), .vdd(vdd), .A(data_in[10]), .B(next_b_data_in_prev_10_), .S(_0__bF_buf5), .Y(_12938_) );
OAI21X1 OAI21X1_3673 ( .gnd(gnd), .vdd(vdd), .A(_12938_), .B(_12916__bF_buf21), .C(_12937_), .Y(_12914__10_) );
NAND2X1 NAND2X1_1708 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_11_), .B(_12916__bF_buf20), .Y(_12939_) );
MUX2X1 MUX2X1_48 ( .gnd(gnd), .vdd(vdd), .A(data_in[11]), .B(next_b_data_in_prev_11_), .S(_0__bF_buf4), .Y(_12940_) );
OAI21X1 OAI21X1_3674 ( .gnd(gnd), .vdd(vdd), .A(_12940_), .B(_12916__bF_buf19), .C(_12939_), .Y(_12914__11_) );
NAND2X1 NAND2X1_1709 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_12_), .B(_12916__bF_buf18), .Y(_12941_) );
MUX2X1 MUX2X1_49 ( .gnd(gnd), .vdd(vdd), .A(data_in[12]), .B(next_b_data_in_prev_12_), .S(_0__bF_buf3), .Y(_12942_) );
OAI21X1 OAI21X1_3675 ( .gnd(gnd), .vdd(vdd), .A(_12942_), .B(_12916__bF_buf17), .C(_12941_), .Y(_12914__12_) );
NAND2X1 NAND2X1_1710 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_13_), .B(_12916__bF_buf16), .Y(_12943_) );
MUX2X1 MUX2X1_50 ( .gnd(gnd), .vdd(vdd), .A(data_in[13]), .B(next_b_data_in_prev_13_), .S(_0__bF_buf2), .Y(_12944_) );
OAI21X1 OAI21X1_3676 ( .gnd(gnd), .vdd(vdd), .A(_12944_), .B(_12916__bF_buf15), .C(_12943_), .Y(_12914__13_) );
NAND2X1 NAND2X1_1711 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_14_), .B(_12916__bF_buf14), .Y(_12945_) );
MUX2X1 MUX2X1_51 ( .gnd(gnd), .vdd(vdd), .A(data_in[14]), .B(next_b_data_in_prev_14_), .S(_0__bF_buf1), .Y(_12946_) );
OAI21X1 OAI21X1_3677 ( .gnd(gnd), .vdd(vdd), .A(_12946_), .B(_12916__bF_buf13), .C(_12945_), .Y(_12914__14_) );
NAND2X1 NAND2X1_1712 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_15_), .B(_12916__bF_buf12), .Y(_12947_) );
MUX2X1 MUX2X1_52 ( .gnd(gnd), .vdd(vdd), .A(data_in[15]), .B(next_b_data_in_prev_15_), .S(_0__bF_buf0), .Y(_12948_) );
OAI21X1 OAI21X1_3678 ( .gnd(gnd), .vdd(vdd), .A(_12948_), .B(_12916__bF_buf11), .C(_12947_), .Y(_12914__15_) );
NAND2X1 NAND2X1_1713 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_16_), .B(_12916__bF_buf10), .Y(_12949_) );
MUX2X1 MUX2X1_53 ( .gnd(gnd), .vdd(vdd), .A(data_in[16]), .B(next_b_data_in_prev_16_), .S(_0__bF_buf9), .Y(_12950_) );
OAI21X1 OAI21X1_3679 ( .gnd(gnd), .vdd(vdd), .A(_12950_), .B(_12916__bF_buf9), .C(_12949_), .Y(_12914__16_) );
NAND2X1 NAND2X1_1714 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_17_), .B(_12916__bF_buf8), .Y(_12951_) );
MUX2X1 MUX2X1_54 ( .gnd(gnd), .vdd(vdd), .A(data_in[17]), .B(next_b_data_in_prev_17_), .S(_0__bF_buf8), .Y(_12952_) );
OAI21X1 OAI21X1_3680 ( .gnd(gnd), .vdd(vdd), .A(_12952_), .B(_12916__bF_buf7), .C(_12951_), .Y(_12914__17_) );
NAND2X1 NAND2X1_1715 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_18_), .B(_12916__bF_buf6), .Y(_12953_) );
MUX2X1 MUX2X1_55 ( .gnd(gnd), .vdd(vdd), .A(data_in[18]), .B(next_b_data_in_prev_18_), .S(_0__bF_buf7), .Y(_12954_) );
OAI21X1 OAI21X1_3681 ( .gnd(gnd), .vdd(vdd), .A(_12954_), .B(_12916__bF_buf5), .C(_12953_), .Y(_12914__18_) );
NAND2X1 NAND2X1_1716 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_19_), .B(_12916__bF_buf4), .Y(_12955_) );
MUX2X1 MUX2X1_56 ( .gnd(gnd), .vdd(vdd), .A(data_in[19]), .B(next_b_data_in_prev_19_), .S(_0__bF_buf6), .Y(_12956_) );
OAI21X1 OAI21X1_3682 ( .gnd(gnd), .vdd(vdd), .A(_12956_), .B(_12916__bF_buf3), .C(_12955_), .Y(_12914__19_) );
NAND2X1 NAND2X1_1717 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_20_), .B(_12916__bF_buf2), .Y(_12957_) );
MUX2X1 MUX2X1_57 ( .gnd(gnd), .vdd(vdd), .A(data_in[20]), .B(next_b_data_in_prev_20_), .S(_0__bF_buf5), .Y(_12958_) );
OAI21X1 OAI21X1_3683 ( .gnd(gnd), .vdd(vdd), .A(_12958_), .B(_12916__bF_buf1), .C(_12957_), .Y(_12914__20_) );
NAND2X1 NAND2X1_1718 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_21_), .B(_12916__bF_buf0), .Y(_12959_) );
MUX2X1 MUX2X1_58 ( .gnd(gnd), .vdd(vdd), .A(data_in[21]), .B(next_b_data_in_prev_21_), .S(_0__bF_buf4), .Y(_12960_) );
OAI21X1 OAI21X1_3684 ( .gnd(gnd), .vdd(vdd), .A(_12960_), .B(_12916__bF_buf42), .C(_12959_), .Y(_12914__21_) );
NAND2X1 NAND2X1_1719 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_22_), .B(_12916__bF_buf41), .Y(_12961_) );
MUX2X1 MUX2X1_59 ( .gnd(gnd), .vdd(vdd), .A(data_in[22]), .B(next_b_data_in_prev_22_), .S(_0__bF_buf3), .Y(_12962_) );
OAI21X1 OAI21X1_3685 ( .gnd(gnd), .vdd(vdd), .A(_12962_), .B(_12916__bF_buf40), .C(_12961_), .Y(_12914__22_) );
NAND2X1 NAND2X1_1720 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_23_), .B(_12916__bF_buf39), .Y(_12963_) );
MUX2X1 MUX2X1_60 ( .gnd(gnd), .vdd(vdd), .A(data_in[23]), .B(next_b_data_in_prev_23_), .S(_0__bF_buf2), .Y(_12964_) );
OAI21X1 OAI21X1_3686 ( .gnd(gnd), .vdd(vdd), .A(_12964_), .B(_12916__bF_buf38), .C(_12963_), .Y(_12914__23_) );
NAND2X1 NAND2X1_1721 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_24_), .B(_12916__bF_buf37), .Y(_12965_) );
MUX2X1 MUX2X1_61 ( .gnd(gnd), .vdd(vdd), .A(data_in[24]), .B(next_b_data_in_prev_24_), .S(_0__bF_buf1), .Y(_12966_) );
OAI21X1 OAI21X1_3687 ( .gnd(gnd), .vdd(vdd), .A(_12966_), .B(_12916__bF_buf36), .C(_12965_), .Y(_12914__24_) );
NAND2X1 NAND2X1_1722 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_25_), .B(_12916__bF_buf35), .Y(_12967_) );
MUX2X1 MUX2X1_62 ( .gnd(gnd), .vdd(vdd), .A(data_in[25]), .B(next_b_data_in_prev_25_), .S(_0__bF_buf0), .Y(_12968_) );
OAI21X1 OAI21X1_3688 ( .gnd(gnd), .vdd(vdd), .A(_12968_), .B(_12916__bF_buf34), .C(_12967_), .Y(_12914__25_) );
NAND2X1 NAND2X1_1723 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_26_), .B(_12916__bF_buf33), .Y(_12969_) );
MUX2X1 MUX2X1_63 ( .gnd(gnd), .vdd(vdd), .A(data_in[26]), .B(next_b_data_in_prev_26_), .S(_0__bF_buf9), .Y(_12970_) );
OAI21X1 OAI21X1_3689 ( .gnd(gnd), .vdd(vdd), .A(_12970_), .B(_12916__bF_buf32), .C(_12969_), .Y(_12914__26_) );
NAND2X1 NAND2X1_1724 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_27_), .B(_12916__bF_buf31), .Y(_12971_) );
MUX2X1 MUX2X1_64 ( .gnd(gnd), .vdd(vdd), .A(data_in[27]), .B(next_b_data_in_prev_27_), .S(_0__bF_buf8), .Y(_12972_) );
OAI21X1 OAI21X1_3690 ( .gnd(gnd), .vdd(vdd), .A(_12972_), .B(_12916__bF_buf30), .C(_12971_), .Y(_12914__27_) );
NAND2X1 NAND2X1_1725 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_28_), .B(_12916__bF_buf29), .Y(_12973_) );
MUX2X1 MUX2X1_65 ( .gnd(gnd), .vdd(vdd), .A(data_in[28]), .B(next_b_data_in_prev_28_), .S(_0__bF_buf7), .Y(_12974_) );
OAI21X1 OAI21X1_3691 ( .gnd(gnd), .vdd(vdd), .A(_12974_), .B(_12916__bF_buf28), .C(_12973_), .Y(_12914__28_) );
NAND2X1 NAND2X1_1726 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_29_), .B(_12916__bF_buf27), .Y(_12975_) );
MUX2X1 MUX2X1_66 ( .gnd(gnd), .vdd(vdd), .A(data_in[29]), .B(next_b_data_in_prev_29_), .S(_0__bF_buf6), .Y(_12976_) );
OAI21X1 OAI21X1_3692 ( .gnd(gnd), .vdd(vdd), .A(_12976_), .B(_12916__bF_buf26), .C(_12975_), .Y(_12914__29_) );
NAND2X1 NAND2X1_1727 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_30_), .B(_12916__bF_buf25), .Y(_12977_) );
MUX2X1 MUX2X1_67 ( .gnd(gnd), .vdd(vdd), .A(data_in[30]), .B(next_b_data_in_prev_30_), .S(_0__bF_buf5), .Y(_12978_) );
OAI21X1 OAI21X1_3693 ( .gnd(gnd), .vdd(vdd), .A(_12978_), .B(_12916__bF_buf24), .C(_12977_), .Y(_12914__30_) );
NAND2X1 NAND2X1_1728 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_31_), .B(_12916__bF_buf23), .Y(_12979_) );
MUX2X1 MUX2X1_68 ( .gnd(gnd), .vdd(vdd), .A(data_in[31]), .B(next_b_data_in_prev_31_), .S(_0__bF_buf4), .Y(_12980_) );
OAI21X1 OAI21X1_3694 ( .gnd(gnd), .vdd(vdd), .A(_12980_), .B(_12916__bF_buf22), .C(_12979_), .Y(_12914__31_) );
NAND2X1 NAND2X1_1729 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_32_), .B(_12916__bF_buf21), .Y(_12981_) );
MUX2X1 MUX2X1_69 ( .gnd(gnd), .vdd(vdd), .A(data_in[32]), .B(next_b_data_in_prev_32_), .S(_0__bF_buf3), .Y(_12982_) );
OAI21X1 OAI21X1_3695 ( .gnd(gnd), .vdd(vdd), .A(_12982_), .B(_12916__bF_buf20), .C(_12981_), .Y(_12914__32_) );
NAND2X1 NAND2X1_1730 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_33_), .B(_12916__bF_buf19), .Y(_12983_) );
MUX2X1 MUX2X1_70 ( .gnd(gnd), .vdd(vdd), .A(data_in[33]), .B(next_b_data_in_prev_33_), .S(_0__bF_buf2), .Y(_12984_) );
OAI21X1 OAI21X1_3696 ( .gnd(gnd), .vdd(vdd), .A(_12984_), .B(_12916__bF_buf18), .C(_12983_), .Y(_12914__33_) );
NAND2X1 NAND2X1_1731 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_34_), .B(_12916__bF_buf17), .Y(_12985_) );
MUX2X1 MUX2X1_71 ( .gnd(gnd), .vdd(vdd), .A(data_in[34]), .B(next_b_data_in_prev_34_), .S(_0__bF_buf1), .Y(_12986_) );
OAI21X1 OAI21X1_3697 ( .gnd(gnd), .vdd(vdd), .A(_12986_), .B(_12916__bF_buf16), .C(_12985_), .Y(_12914__34_) );
NAND2X1 NAND2X1_1732 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_35_), .B(_12916__bF_buf15), .Y(_12987_) );
MUX2X1 MUX2X1_72 ( .gnd(gnd), .vdd(vdd), .A(data_in[35]), .B(next_b_data_in_prev_35_), .S(_0__bF_buf0), .Y(_12988_) );
OAI21X1 OAI21X1_3698 ( .gnd(gnd), .vdd(vdd), .A(_12988_), .B(_12916__bF_buf14), .C(_12987_), .Y(_12914__35_) );
NAND2X1 NAND2X1_1733 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_36_), .B(_12916__bF_buf13), .Y(_12989_) );
MUX2X1 MUX2X1_73 ( .gnd(gnd), .vdd(vdd), .A(data_in[36]), .B(next_b_data_in_prev_36_), .S(_0__bF_buf9), .Y(_12990_) );
OAI21X1 OAI21X1_3699 ( .gnd(gnd), .vdd(vdd), .A(_12990_), .B(_12916__bF_buf12), .C(_12989_), .Y(_12914__36_) );
NAND2X1 NAND2X1_1734 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_37_), .B(_12916__bF_buf11), .Y(_12991_) );
MUX2X1 MUX2X1_74 ( .gnd(gnd), .vdd(vdd), .A(data_in[37]), .B(next_b_data_in_prev_37_), .S(_0__bF_buf8), .Y(_12992_) );
OAI21X1 OAI21X1_3700 ( .gnd(gnd), .vdd(vdd), .A(_12992_), .B(_12916__bF_buf10), .C(_12991_), .Y(_12914__37_) );
NAND2X1 NAND2X1_1735 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_38_), .B(_12916__bF_buf9), .Y(_12993_) );
MUX2X1 MUX2X1_75 ( .gnd(gnd), .vdd(vdd), .A(data_in[38]), .B(next_b_data_in_prev_38_), .S(_0__bF_buf7), .Y(_12994_) );
OAI21X1 OAI21X1_3701 ( .gnd(gnd), .vdd(vdd), .A(_12994_), .B(_12916__bF_buf8), .C(_12993_), .Y(_12914__38_) );
NAND2X1 NAND2X1_1736 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_39_), .B(_12916__bF_buf7), .Y(_12995_) );
MUX2X1 MUX2X1_76 ( .gnd(gnd), .vdd(vdd), .A(data_in[39]), .B(next_b_data_in_prev_39_), .S(_0__bF_buf6), .Y(_12996_) );
OAI21X1 OAI21X1_3702 ( .gnd(gnd), .vdd(vdd), .A(_12996_), .B(_12916__bF_buf6), .C(_12995_), .Y(_12914__39_) );
NAND2X1 NAND2X1_1737 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_40_), .B(_12916__bF_buf5), .Y(_12997_) );
MUX2X1 MUX2X1_77 ( .gnd(gnd), .vdd(vdd), .A(data_in[40]), .B(next_b_data_in_prev_40_), .S(_0__bF_buf5), .Y(_12998_) );
OAI21X1 OAI21X1_3703 ( .gnd(gnd), .vdd(vdd), .A(_12998_), .B(_12916__bF_buf4), .C(_12997_), .Y(_12914__40_) );
NAND2X1 NAND2X1_1738 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_41_), .B(_12916__bF_buf3), .Y(_12999_) );
MUX2X1 MUX2X1_78 ( .gnd(gnd), .vdd(vdd), .A(data_in[41]), .B(next_b_data_in_prev_41_), .S(_0__bF_buf4), .Y(_13000_) );
OAI21X1 OAI21X1_3704 ( .gnd(gnd), .vdd(vdd), .A(_13000_), .B(_12916__bF_buf2), .C(_12999_), .Y(_12914__41_) );
NAND2X1 NAND2X1_1739 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_42_), .B(_12916__bF_buf1), .Y(_13001_) );
MUX2X1 MUX2X1_79 ( .gnd(gnd), .vdd(vdd), .A(data_in[42]), .B(next_b_data_in_prev_42_), .S(_0__bF_buf3), .Y(_13002_) );
OAI21X1 OAI21X1_3705 ( .gnd(gnd), .vdd(vdd), .A(_13002_), .B(_12916__bF_buf0), .C(_13001_), .Y(_12914__42_) );
NAND2X1 NAND2X1_1740 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_43_), .B(_12916__bF_buf42), .Y(_13003_) );
MUX2X1 MUX2X1_80 ( .gnd(gnd), .vdd(vdd), .A(data_in[43]), .B(next_b_data_in_prev_43_), .S(_0__bF_buf2), .Y(_13004_) );
OAI21X1 OAI21X1_3706 ( .gnd(gnd), .vdd(vdd), .A(_13004_), .B(_12916__bF_buf41), .C(_13003_), .Y(_12914__43_) );
NAND2X1 NAND2X1_1741 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_44_), .B(_12916__bF_buf40), .Y(_13005_) );
MUX2X1 MUX2X1_81 ( .gnd(gnd), .vdd(vdd), .A(data_in[44]), .B(next_b_data_in_prev_44_), .S(_0__bF_buf1), .Y(_13006_) );
OAI21X1 OAI21X1_3707 ( .gnd(gnd), .vdd(vdd), .A(_13006_), .B(_12916__bF_buf39), .C(_13005_), .Y(_12914__44_) );
NAND2X1 NAND2X1_1742 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_45_), .B(_12916__bF_buf38), .Y(_13007_) );
MUX2X1 MUX2X1_82 ( .gnd(gnd), .vdd(vdd), .A(data_in[45]), .B(next_b_data_in_prev_45_), .S(_0__bF_buf0), .Y(_13008_) );
OAI21X1 OAI21X1_3708 ( .gnd(gnd), .vdd(vdd), .A(_13008_), .B(_12916__bF_buf37), .C(_13007_), .Y(_12914__45_) );
NAND2X1 NAND2X1_1743 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_46_), .B(_12916__bF_buf36), .Y(_13009_) );
MUX2X1 MUX2X1_83 ( .gnd(gnd), .vdd(vdd), .A(data_in[46]), .B(next_b_data_in_prev_46_), .S(_0__bF_buf9), .Y(_13010_) );
OAI21X1 OAI21X1_3709 ( .gnd(gnd), .vdd(vdd), .A(_13010_), .B(_12916__bF_buf35), .C(_13009_), .Y(_12914__46_) );
NAND2X1 NAND2X1_1744 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_47_), .B(_12916__bF_buf34), .Y(_13011_) );
MUX2X1 MUX2X1_84 ( .gnd(gnd), .vdd(vdd), .A(data_in[47]), .B(next_b_data_in_prev_47_), .S(_0__bF_buf8), .Y(_13012_) );
OAI21X1 OAI21X1_3710 ( .gnd(gnd), .vdd(vdd), .A(_13012_), .B(_12916__bF_buf33), .C(_13011_), .Y(_12914__47_) );
NAND2X1 NAND2X1_1745 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_48_), .B(_12916__bF_buf32), .Y(_13013_) );
MUX2X1 MUX2X1_85 ( .gnd(gnd), .vdd(vdd), .A(data_in[48]), .B(next_b_data_in_prev_48_), .S(_0__bF_buf7), .Y(_13014_) );
OAI21X1 OAI21X1_3711 ( .gnd(gnd), .vdd(vdd), .A(_13014_), .B(_12916__bF_buf31), .C(_13013_), .Y(_12914__48_) );
NAND2X1 NAND2X1_1746 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_49_), .B(_12916__bF_buf30), .Y(_13015_) );
MUX2X1 MUX2X1_86 ( .gnd(gnd), .vdd(vdd), .A(data_in[49]), .B(next_b_data_in_prev_49_), .S(_0__bF_buf6), .Y(_13016_) );
OAI21X1 OAI21X1_3712 ( .gnd(gnd), .vdd(vdd), .A(_13016_), .B(_12916__bF_buf29), .C(_13015_), .Y(_12914__49_) );
NAND2X1 NAND2X1_1747 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_50_), .B(_12916__bF_buf28), .Y(_13017_) );
MUX2X1 MUX2X1_87 ( .gnd(gnd), .vdd(vdd), .A(data_in[50]), .B(next_b_data_in_prev_50_), .S(_0__bF_buf5), .Y(_13018_) );
OAI21X1 OAI21X1_3713 ( .gnd(gnd), .vdd(vdd), .A(_13018_), .B(_12916__bF_buf27), .C(_13017_), .Y(_12914__50_) );
NAND2X1 NAND2X1_1748 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_51_), .B(_12916__bF_buf26), .Y(_13019_) );
MUX2X1 MUX2X1_88 ( .gnd(gnd), .vdd(vdd), .A(data_in[51]), .B(next_b_data_in_prev_51_), .S(_0__bF_buf4), .Y(_13020_) );
OAI21X1 OAI21X1_3714 ( .gnd(gnd), .vdd(vdd), .A(_13020_), .B(_12916__bF_buf25), .C(_13019_), .Y(_12914__51_) );
NAND2X1 NAND2X1_1749 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_52_), .B(_12916__bF_buf24), .Y(_13021_) );
MUX2X1 MUX2X1_89 ( .gnd(gnd), .vdd(vdd), .A(data_in[52]), .B(next_b_data_in_prev_52_), .S(_0__bF_buf3), .Y(_13022_) );
OAI21X1 OAI21X1_3715 ( .gnd(gnd), .vdd(vdd), .A(_13022_), .B(_12916__bF_buf23), .C(_13021_), .Y(_12914__52_) );
NAND2X1 NAND2X1_1750 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_53_), .B(_12916__bF_buf22), .Y(_13023_) );
MUX2X1 MUX2X1_90 ( .gnd(gnd), .vdd(vdd), .A(data_in[53]), .B(next_b_data_in_prev_53_), .S(_0__bF_buf2), .Y(_13024_) );
OAI21X1 OAI21X1_3716 ( .gnd(gnd), .vdd(vdd), .A(_13024_), .B(_12916__bF_buf21), .C(_13023_), .Y(_12914__53_) );
NAND2X1 NAND2X1_1751 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_54_), .B(_12916__bF_buf20), .Y(_13025_) );
MUX2X1 MUX2X1_91 ( .gnd(gnd), .vdd(vdd), .A(data_in[54]), .B(next_b_data_in_prev_54_), .S(_0__bF_buf1), .Y(_13026_) );
OAI21X1 OAI21X1_3717 ( .gnd(gnd), .vdd(vdd), .A(_13026_), .B(_12916__bF_buf19), .C(_13025_), .Y(_12914__54_) );
NAND2X1 NAND2X1_1752 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_55_), .B(_12916__bF_buf18), .Y(_13027_) );
MUX2X1 MUX2X1_92 ( .gnd(gnd), .vdd(vdd), .A(data_in[55]), .B(next_b_data_in_prev_55_), .S(_0__bF_buf0), .Y(_13028_) );
OAI21X1 OAI21X1_3718 ( .gnd(gnd), .vdd(vdd), .A(_13028_), .B(_12916__bF_buf17), .C(_13027_), .Y(_12914__55_) );
NAND2X1 NAND2X1_1753 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_56_), .B(_12916__bF_buf16), .Y(_13029_) );
MUX2X1 MUX2X1_93 ( .gnd(gnd), .vdd(vdd), .A(data_in[56]), .B(next_b_data_in_prev_56_), .S(_0__bF_buf9), .Y(_13030_) );
OAI21X1 OAI21X1_3719 ( .gnd(gnd), .vdd(vdd), .A(_13030_), .B(_12916__bF_buf15), .C(_13029_), .Y(_12914__56_) );
NAND2X1 NAND2X1_1754 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_57_), .B(_12916__bF_buf14), .Y(_13031_) );
MUX2X1 MUX2X1_94 ( .gnd(gnd), .vdd(vdd), .A(data_in[57]), .B(next_b_data_in_prev_57_), .S(_0__bF_buf8), .Y(_13032_) );
OAI21X1 OAI21X1_3720 ( .gnd(gnd), .vdd(vdd), .A(_13032_), .B(_12916__bF_buf13), .C(_13031_), .Y(_12914__57_) );
NAND2X1 NAND2X1_1755 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_58_), .B(_12916__bF_buf12), .Y(_13033_) );
MUX2X1 MUX2X1_95 ( .gnd(gnd), .vdd(vdd), .A(data_in[58]), .B(next_b_data_in_prev_58_), .S(_0__bF_buf7), .Y(_13034_) );
OAI21X1 OAI21X1_3721 ( .gnd(gnd), .vdd(vdd), .A(_13034_), .B(_12916__bF_buf11), .C(_13033_), .Y(_12914__58_) );
NAND2X1 NAND2X1_1756 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_59_), .B(_12916__bF_buf10), .Y(_13035_) );
MUX2X1 MUX2X1_96 ( .gnd(gnd), .vdd(vdd), .A(data_in[59]), .B(next_b_data_in_prev_59_), .S(_0__bF_buf6), .Y(_13036_) );
OAI21X1 OAI21X1_3722 ( .gnd(gnd), .vdd(vdd), .A(_13036_), .B(_12916__bF_buf9), .C(_13035_), .Y(_12914__59_) );
NAND2X1 NAND2X1_1757 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_60_), .B(_12916__bF_buf8), .Y(_13037_) );
MUX2X1 MUX2X1_97 ( .gnd(gnd), .vdd(vdd), .A(data_in[60]), .B(next_b_data_in_prev_60_), .S(_0__bF_buf5), .Y(_13038_) );
OAI21X1 OAI21X1_3723 ( .gnd(gnd), .vdd(vdd), .A(_13038_), .B(_12916__bF_buf7), .C(_13037_), .Y(_12914__60_) );
NAND2X1 NAND2X1_1758 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_61_), .B(_12916__bF_buf6), .Y(_13039_) );
MUX2X1 MUX2X1_98 ( .gnd(gnd), .vdd(vdd), .A(data_in[61]), .B(next_b_data_in_prev_61_), .S(_0__bF_buf4), .Y(_13040_) );
OAI21X1 OAI21X1_3724 ( .gnd(gnd), .vdd(vdd), .A(_13040_), .B(_12916__bF_buf5), .C(_13039_), .Y(_12914__61_) );
NAND2X1 NAND2X1_1759 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_62_), .B(_12916__bF_buf4), .Y(_13041_) );
MUX2X1 MUX2X1_99 ( .gnd(gnd), .vdd(vdd), .A(data_in[62]), .B(next_b_data_in_prev_62_), .S(_0__bF_buf3), .Y(_13042_) );
OAI21X1 OAI21X1_3725 ( .gnd(gnd), .vdd(vdd), .A(_13042_), .B(_12916__bF_buf3), .C(_13041_), .Y(_12914__62_) );
NAND2X1 NAND2X1_1760 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_63_), .B(_12916__bF_buf2), .Y(_13043_) );
MUX2X1 MUX2X1_100 ( .gnd(gnd), .vdd(vdd), .A(data_in[63]), .B(next_b_data_in_prev_63_), .S(_0__bF_buf2), .Y(_13044_) );
OAI21X1 OAI21X1_3726 ( .gnd(gnd), .vdd(vdd), .A(_13044_), .B(_12916__bF_buf1), .C(_13043_), .Y(_12914__63_) );
NAND2X1 NAND2X1_1761 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_64_), .B(_12916__bF_buf0), .Y(_13045_) );
MUX2X1 MUX2X1_101 ( .gnd(gnd), .vdd(vdd), .A(data_in[64]), .B(next_b_data_in_prev_64_), .S(_0__bF_buf1), .Y(_13046_) );
OAI21X1 OAI21X1_3727 ( .gnd(gnd), .vdd(vdd), .A(_13046_), .B(_12916__bF_buf42), .C(_13045_), .Y(_12914__64_) );
NAND2X1 NAND2X1_1762 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_65_), .B(_12916__bF_buf41), .Y(_13047_) );
MUX2X1 MUX2X1_102 ( .gnd(gnd), .vdd(vdd), .A(data_in[65]), .B(next_b_data_in_prev_65_), .S(_0__bF_buf0), .Y(_13048_) );
OAI21X1 OAI21X1_3728 ( .gnd(gnd), .vdd(vdd), .A(_13048_), .B(_12916__bF_buf40), .C(_13047_), .Y(_12914__65_) );
NAND2X1 NAND2X1_1763 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_66_), .B(_12916__bF_buf39), .Y(_13049_) );
MUX2X1 MUX2X1_103 ( .gnd(gnd), .vdd(vdd), .A(data_in[66]), .B(next_b_data_in_prev_66_), .S(_0__bF_buf9), .Y(_13050_) );
OAI21X1 OAI21X1_3729 ( .gnd(gnd), .vdd(vdd), .A(_13050_), .B(_12916__bF_buf38), .C(_13049_), .Y(_12914__66_) );
NAND2X1 NAND2X1_1764 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_67_), .B(_12916__bF_buf37), .Y(_13051_) );
MUX2X1 MUX2X1_104 ( .gnd(gnd), .vdd(vdd), .A(data_in[67]), .B(next_b_data_in_prev_67_), .S(_0__bF_buf8), .Y(_13052_) );
OAI21X1 OAI21X1_3730 ( .gnd(gnd), .vdd(vdd), .A(_13052_), .B(_12916__bF_buf36), .C(_13051_), .Y(_12914__67_) );
NAND2X1 NAND2X1_1765 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_68_), .B(_12916__bF_buf35), .Y(_13053_) );
MUX2X1 MUX2X1_105 ( .gnd(gnd), .vdd(vdd), .A(data_in[68]), .B(next_b_data_in_prev_68_), .S(_0__bF_buf7), .Y(_13054_) );
OAI21X1 OAI21X1_3731 ( .gnd(gnd), .vdd(vdd), .A(_13054_), .B(_12916__bF_buf34), .C(_13053_), .Y(_12914__68_) );
NAND2X1 NAND2X1_1766 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_69_), .B(_12916__bF_buf33), .Y(_13055_) );
MUX2X1 MUX2X1_106 ( .gnd(gnd), .vdd(vdd), .A(data_in[69]), .B(next_b_data_in_prev_69_), .S(_0__bF_buf6), .Y(_13056_) );
OAI21X1 OAI21X1_3732 ( .gnd(gnd), .vdd(vdd), .A(_13056_), .B(_12916__bF_buf32), .C(_13055_), .Y(_12914__69_) );
NAND2X1 NAND2X1_1767 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_70_), .B(_12916__bF_buf31), .Y(_13057_) );
MUX2X1 MUX2X1_107 ( .gnd(gnd), .vdd(vdd), .A(data_in[70]), .B(next_b_data_in_prev_70_), .S(_0__bF_buf5), .Y(_13058_) );
OAI21X1 OAI21X1_3733 ( .gnd(gnd), .vdd(vdd), .A(_13058_), .B(_12916__bF_buf30), .C(_13057_), .Y(_12914__70_) );
NAND2X1 NAND2X1_1768 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_71_), .B(_12916__bF_buf29), .Y(_13059_) );
MUX2X1 MUX2X1_108 ( .gnd(gnd), .vdd(vdd), .A(data_in[71]), .B(next_b_data_in_prev_71_), .S(_0__bF_buf4), .Y(_13060_) );
OAI21X1 OAI21X1_3734 ( .gnd(gnd), .vdd(vdd), .A(_13060_), .B(_12916__bF_buf28), .C(_13059_), .Y(_12914__71_) );
NAND2X1 NAND2X1_1769 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_72_), .B(_12916__bF_buf27), .Y(_13061_) );
MUX2X1 MUX2X1_109 ( .gnd(gnd), .vdd(vdd), .A(data_in[72]), .B(next_b_data_in_prev_72_), .S(_0__bF_buf3), .Y(_13062_) );
OAI21X1 OAI21X1_3735 ( .gnd(gnd), .vdd(vdd), .A(_13062_), .B(_12916__bF_buf26), .C(_13061_), .Y(_12914__72_) );
NAND2X1 NAND2X1_1770 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_73_), .B(_12916__bF_buf25), .Y(_13063_) );
MUX2X1 MUX2X1_110 ( .gnd(gnd), .vdd(vdd), .A(data_in[73]), .B(next_b_data_in_prev_73_), .S(_0__bF_buf2), .Y(_13064_) );
OAI21X1 OAI21X1_3736 ( .gnd(gnd), .vdd(vdd), .A(_13064_), .B(_12916__bF_buf24), .C(_13063_), .Y(_12914__73_) );
NAND2X1 NAND2X1_1771 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_74_), .B(_12916__bF_buf23), .Y(_13065_) );
MUX2X1 MUX2X1_111 ( .gnd(gnd), .vdd(vdd), .A(data_in[74]), .B(next_b_data_in_prev_74_), .S(_0__bF_buf1), .Y(_13066_) );
OAI21X1 OAI21X1_3737 ( .gnd(gnd), .vdd(vdd), .A(_13066_), .B(_12916__bF_buf22), .C(_13065_), .Y(_12914__74_) );
NAND2X1 NAND2X1_1772 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_75_), .B(_12916__bF_buf21), .Y(_13067_) );
MUX2X1 MUX2X1_112 ( .gnd(gnd), .vdd(vdd), .A(data_in[75]), .B(next_b_data_in_prev_75_), .S(_0__bF_buf0), .Y(_13068_) );
OAI21X1 OAI21X1_3738 ( .gnd(gnd), .vdd(vdd), .A(_13068_), .B(_12916__bF_buf20), .C(_13067_), .Y(_12914__75_) );
NAND2X1 NAND2X1_1773 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_76_), .B(_12916__bF_buf19), .Y(_13069_) );
MUX2X1 MUX2X1_113 ( .gnd(gnd), .vdd(vdd), .A(data_in[76]), .B(next_b_data_in_prev_76_), .S(_0__bF_buf9), .Y(_13070_) );
OAI21X1 OAI21X1_3739 ( .gnd(gnd), .vdd(vdd), .A(_13070_), .B(_12916__bF_buf18), .C(_13069_), .Y(_12914__76_) );
NAND2X1 NAND2X1_1774 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_77_), .B(_12916__bF_buf17), .Y(_13071_) );
MUX2X1 MUX2X1_114 ( .gnd(gnd), .vdd(vdd), .A(data_in[77]), .B(next_b_data_in_prev_77_), .S(_0__bF_buf8), .Y(_13072_) );
OAI21X1 OAI21X1_3740 ( .gnd(gnd), .vdd(vdd), .A(_13072_), .B(_12916__bF_buf16), .C(_13071_), .Y(_12914__77_) );
NAND2X1 NAND2X1_1775 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_78_), .B(_12916__bF_buf15), .Y(_13073_) );
MUX2X1 MUX2X1_115 ( .gnd(gnd), .vdd(vdd), .A(data_in[78]), .B(next_b_data_in_prev_78_), .S(_0__bF_buf7), .Y(_13074_) );
OAI21X1 OAI21X1_3741 ( .gnd(gnd), .vdd(vdd), .A(_13074_), .B(_12916__bF_buf14), .C(_13073_), .Y(_12914__78_) );
NAND2X1 NAND2X1_1776 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_79_), .B(_12916__bF_buf13), .Y(_13075_) );
MUX2X1 MUX2X1_116 ( .gnd(gnd), .vdd(vdd), .A(data_in[79]), .B(next_b_data_in_prev_79_), .S(_0__bF_buf6), .Y(_13076_) );
OAI21X1 OAI21X1_3742 ( .gnd(gnd), .vdd(vdd), .A(_13076_), .B(_12916__bF_buf12), .C(_13075_), .Y(_12914__79_) );
NAND2X1 NAND2X1_1777 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_80_), .B(_12916__bF_buf11), .Y(_13077_) );
MUX2X1 MUX2X1_117 ( .gnd(gnd), .vdd(vdd), .A(data_in[80]), .B(next_b_data_in_prev_80_), .S(_0__bF_buf5), .Y(_13078_) );
OAI21X1 OAI21X1_3743 ( .gnd(gnd), .vdd(vdd), .A(_13078_), .B(_12916__bF_buf10), .C(_13077_), .Y(_12914__80_) );
NAND2X1 NAND2X1_1778 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_81_), .B(_12916__bF_buf9), .Y(_13079_) );
MUX2X1 MUX2X1_118 ( .gnd(gnd), .vdd(vdd), .A(data_in[81]), .B(next_b_data_in_prev_81_), .S(_0__bF_buf4), .Y(_13080_) );
OAI21X1 OAI21X1_3744 ( .gnd(gnd), .vdd(vdd), .A(_13080_), .B(_12916__bF_buf8), .C(_13079_), .Y(_12914__81_) );
NAND2X1 NAND2X1_1779 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_82_), .B(_12916__bF_buf7), .Y(_13081_) );
MUX2X1 MUX2X1_119 ( .gnd(gnd), .vdd(vdd), .A(data_in[82]), .B(next_b_data_in_prev_82_), .S(_0__bF_buf3), .Y(_13082_) );
OAI21X1 OAI21X1_3745 ( .gnd(gnd), .vdd(vdd), .A(_13082_), .B(_12916__bF_buf6), .C(_13081_), .Y(_12914__82_) );
NAND2X1 NAND2X1_1780 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_83_), .B(_12916__bF_buf5), .Y(_13083_) );
MUX2X1 MUX2X1_120 ( .gnd(gnd), .vdd(vdd), .A(data_in[83]), .B(next_b_data_in_prev_83_), .S(_0__bF_buf2), .Y(_13084_) );
OAI21X1 OAI21X1_3746 ( .gnd(gnd), .vdd(vdd), .A(_13084_), .B(_12916__bF_buf4), .C(_13083_), .Y(_12914__83_) );
NAND2X1 NAND2X1_1781 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_84_), .B(_12916__bF_buf3), .Y(_13085_) );
MUX2X1 MUX2X1_121 ( .gnd(gnd), .vdd(vdd), .A(data_in[84]), .B(next_b_data_in_prev_84_), .S(_0__bF_buf1), .Y(_13086_) );
OAI21X1 OAI21X1_3747 ( .gnd(gnd), .vdd(vdd), .A(_13086_), .B(_12916__bF_buf2), .C(_13085_), .Y(_12914__84_) );
NAND2X1 NAND2X1_1782 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_85_), .B(_12916__bF_buf1), .Y(_13087_) );
MUX2X1 MUX2X1_122 ( .gnd(gnd), .vdd(vdd), .A(data_in[85]), .B(next_b_data_in_prev_85_), .S(_0__bF_buf0), .Y(_13088_) );
OAI21X1 OAI21X1_3748 ( .gnd(gnd), .vdd(vdd), .A(_13088_), .B(_12916__bF_buf0), .C(_13087_), .Y(_12914__85_) );
NAND2X1 NAND2X1_1783 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_86_), .B(_12916__bF_buf42), .Y(_13089_) );
MUX2X1 MUX2X1_123 ( .gnd(gnd), .vdd(vdd), .A(data_in[86]), .B(next_b_data_in_prev_86_), .S(_0__bF_buf9), .Y(_13090_) );
OAI21X1 OAI21X1_3749 ( .gnd(gnd), .vdd(vdd), .A(_13090_), .B(_12916__bF_buf41), .C(_13089_), .Y(_12914__86_) );
NAND2X1 NAND2X1_1784 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_87_), .B(_12916__bF_buf40), .Y(_13091_) );
MUX2X1 MUX2X1_124 ( .gnd(gnd), .vdd(vdd), .A(data_in[87]), .B(next_b_data_in_prev_87_), .S(_0__bF_buf8), .Y(_13092_) );
OAI21X1 OAI21X1_3750 ( .gnd(gnd), .vdd(vdd), .A(_13092_), .B(_12916__bF_buf39), .C(_13091_), .Y(_12914__87_) );
NAND2X1 NAND2X1_1785 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_88_), .B(_12916__bF_buf38), .Y(_13093_) );
MUX2X1 MUX2X1_125 ( .gnd(gnd), .vdd(vdd), .A(data_in[88]), .B(next_b_data_in_prev_88_), .S(_0__bF_buf7), .Y(_13094_) );
OAI21X1 OAI21X1_3751 ( .gnd(gnd), .vdd(vdd), .A(_13094_), .B(_12916__bF_buf37), .C(_13093_), .Y(_12914__88_) );
NAND2X1 NAND2X1_1786 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_89_), .B(_12916__bF_buf36), .Y(_13095_) );
MUX2X1 MUX2X1_126 ( .gnd(gnd), .vdd(vdd), .A(data_in[89]), .B(next_b_data_in_prev_89_), .S(_0__bF_buf6), .Y(_13096_) );
OAI21X1 OAI21X1_3752 ( .gnd(gnd), .vdd(vdd), .A(_13096_), .B(_12916__bF_buf35), .C(_13095_), .Y(_12914__89_) );
NAND2X1 NAND2X1_1787 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_90_), .B(_12916__bF_buf34), .Y(_13097_) );
MUX2X1 MUX2X1_127 ( .gnd(gnd), .vdd(vdd), .A(data_in[90]), .B(next_b_data_in_prev_90_), .S(_0__bF_buf5), .Y(_13098_) );
OAI21X1 OAI21X1_3753 ( .gnd(gnd), .vdd(vdd), .A(_13098_), .B(_12916__bF_buf33), .C(_13097_), .Y(_12914__90_) );
NAND2X1 NAND2X1_1788 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_91_), .B(_12916__bF_buf32), .Y(_13099_) );
MUX2X1 MUX2X1_128 ( .gnd(gnd), .vdd(vdd), .A(data_in[91]), .B(next_b_data_in_prev_91_), .S(_0__bF_buf4), .Y(_13100_) );
OAI21X1 OAI21X1_3754 ( .gnd(gnd), .vdd(vdd), .A(_13100_), .B(_12916__bF_buf31), .C(_13099_), .Y(_12914__91_) );
NAND2X1 NAND2X1_1789 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_92_), .B(_12916__bF_buf30), .Y(_13101_) );
MUX2X1 MUX2X1_129 ( .gnd(gnd), .vdd(vdd), .A(data_in[92]), .B(next_b_data_in_prev_92_), .S(_0__bF_buf3), .Y(_13102_) );
OAI21X1 OAI21X1_3755 ( .gnd(gnd), .vdd(vdd), .A(_13102_), .B(_12916__bF_buf29), .C(_13101_), .Y(_12914__92_) );
NAND2X1 NAND2X1_1790 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_93_), .B(_12916__bF_buf28), .Y(_13103_) );
MUX2X1 MUX2X1_130 ( .gnd(gnd), .vdd(vdd), .A(data_in[93]), .B(next_b_data_in_prev_93_), .S(_0__bF_buf2), .Y(_13104_) );
OAI21X1 OAI21X1_3756 ( .gnd(gnd), .vdd(vdd), .A(_13104_), .B(_12916__bF_buf27), .C(_13103_), .Y(_12914__93_) );
NAND2X1 NAND2X1_1791 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_94_), .B(_12916__bF_buf26), .Y(_13105_) );
MUX2X1 MUX2X1_131 ( .gnd(gnd), .vdd(vdd), .A(data_in[94]), .B(next_b_data_in_prev_94_), .S(_0__bF_buf1), .Y(_13106_) );
OAI21X1 OAI21X1_3757 ( .gnd(gnd), .vdd(vdd), .A(_13106_), .B(_12916__bF_buf25), .C(_13105_), .Y(_12914__94_) );
NAND2X1 NAND2X1_1792 ( .gnd(gnd), .vdd(vdd), .A(next_b_data_in_prev_95_), .B(_12916__bF_buf24), .Y(_13107_) );
MUX2X1 MUX2X1_132 ( .gnd(gnd), .vdd(vdd), .A(data_in[95]), .B(next_b_data_in_prev_95_), .S(_0__bF_buf0), .Y(_13108_) );
OAI21X1 OAI21X1_3758 ( .gnd(gnd), .vdd(vdd), .A(_13108_), .B(_12916__bF_buf23), .C(_13107_), .Y(_12914__95_) );
NOR2X1 NOR2X1_1993 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf22), .B(_12918_), .Y(_12915__0_) );
NOR2X1 NOR2X1_1994 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf21), .B(_12920_), .Y(_12915__1_) );
NOR2X1 NOR2X1_1995 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf20), .B(_12922_), .Y(_12915__2_) );
NOR2X1 NOR2X1_1996 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf19), .B(_12924_), .Y(_12915__3_) );
NOR2X1 NOR2X1_1997 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf18), .B(_12926_), .Y(_12915__4_) );
NOR2X1 NOR2X1_1998 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf17), .B(_12928_), .Y(_12915__5_) );
NOR2X1 NOR2X1_1999 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf16), .B(_12930_), .Y(_12915__6_) );
NOR2X1 NOR2X1_2000 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf15), .B(_12932_), .Y(_12915__7_) );
NOR2X1 NOR2X1_2001 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf14), .B(_12934_), .Y(_12915__8_) );
NOR2X1 NOR2X1_2002 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf13), .B(_12936_), .Y(_12915__9_) );
NOR2X1 NOR2X1_2003 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf12), .B(_12938_), .Y(_12915__10_) );
NOR2X1 NOR2X1_2004 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf11), .B(_12940_), .Y(_12915__11_) );
NOR2X1 NOR2X1_2005 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf10), .B(_12942_), .Y(_12915__12_) );
NOR2X1 NOR2X1_2006 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf9), .B(_12944_), .Y(_12915__13_) );
NOR2X1 NOR2X1_2007 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf8), .B(_12946_), .Y(_12915__14_) );
NOR2X1 NOR2X1_2008 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf7), .B(_12948_), .Y(_12915__15_) );
NOR2X1 NOR2X1_2009 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf6), .B(_12950_), .Y(_12915__16_) );
NOR2X1 NOR2X1_2010 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf5), .B(_12952_), .Y(_12915__17_) );
NOR2X1 NOR2X1_2011 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf4), .B(_12954_), .Y(_12915__18_) );
NOR2X1 NOR2X1_2012 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf3), .B(_12956_), .Y(_12915__19_) );
NOR2X1 NOR2X1_2013 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf2), .B(_12958_), .Y(_12915__20_) );
NOR2X1 NOR2X1_2014 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf1), .B(_12960_), .Y(_12915__21_) );
NOR2X1 NOR2X1_2015 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf0), .B(_12962_), .Y(_12915__22_) );
NOR2X1 NOR2X1_2016 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf42), .B(_12964_), .Y(_12915__23_) );
NOR2X1 NOR2X1_2017 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf41), .B(_12966_), .Y(_12915__24_) );
NOR2X1 NOR2X1_2018 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf40), .B(_12968_), .Y(_12915__25_) );
NOR2X1 NOR2X1_2019 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf39), .B(_12970_), .Y(_12915__26_) );
NOR2X1 NOR2X1_2020 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf38), .B(_12972_), .Y(_12915__27_) );
NOR2X1 NOR2X1_2021 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf37), .B(_12974_), .Y(_12915__28_) );
NOR2X1 NOR2X1_2022 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf36), .B(_12976_), .Y(_12915__29_) );
NOR2X1 NOR2X1_2023 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf35), .B(_12978_), .Y(_12915__30_) );
NOR2X1 NOR2X1_2024 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf34), .B(_12980_), .Y(_12915__31_) );
NOR2X1 NOR2X1_2025 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf33), .B(_12982_), .Y(_12915__32_) );
NOR2X1 NOR2X1_2026 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf32), .B(_12984_), .Y(_12915__33_) );
NOR2X1 NOR2X1_2027 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf31), .B(_12986_), .Y(_12915__34_) );
NOR2X1 NOR2X1_2028 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf30), .B(_12988_), .Y(_12915__35_) );
NOR2X1 NOR2X1_2029 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf29), .B(_12990_), .Y(_12915__36_) );
NOR2X1 NOR2X1_2030 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf28), .B(_12992_), .Y(_12915__37_) );
NOR2X1 NOR2X1_2031 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf27), .B(_12994_), .Y(_12915__38_) );
NOR2X1 NOR2X1_2032 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf26), .B(_12996_), .Y(_12915__39_) );
NOR2X1 NOR2X1_2033 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf25), .B(_12998_), .Y(_12915__40_) );
NOR2X1 NOR2X1_2034 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf24), .B(_13000_), .Y(_12915__41_) );
NOR2X1 NOR2X1_2035 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf23), .B(_13002_), .Y(_12915__42_) );
NOR2X1 NOR2X1_2036 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf22), .B(_13004_), .Y(_12915__43_) );
NOR2X1 NOR2X1_2037 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf21), .B(_13006_), .Y(_12915__44_) );
NOR2X1 NOR2X1_2038 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf20), .B(_13008_), .Y(_12915__45_) );
NOR2X1 NOR2X1_2039 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf19), .B(_13010_), .Y(_12915__46_) );
NOR2X1 NOR2X1_2040 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf18), .B(_13012_), .Y(_12915__47_) );
NOR2X1 NOR2X1_2041 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf17), .B(_13014_), .Y(_12915__48_) );
NOR2X1 NOR2X1_2042 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf16), .B(_13016_), .Y(_12915__49_) );
NOR2X1 NOR2X1_2043 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf15), .B(_13018_), .Y(_12915__50_) );
NOR2X1 NOR2X1_2044 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf14), .B(_13020_), .Y(_12915__51_) );
NOR2X1 NOR2X1_2045 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf13), .B(_13022_), .Y(_12915__52_) );
NOR2X1 NOR2X1_2046 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf12), .B(_13024_), .Y(_12915__53_) );
NOR2X1 NOR2X1_2047 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf11), .B(_13026_), .Y(_12915__54_) );
NOR2X1 NOR2X1_2048 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf10), .B(_13028_), .Y(_12915__55_) );
NOR2X1 NOR2X1_2049 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf9), .B(_13030_), .Y(_12915__56_) );
NOR2X1 NOR2X1_2050 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf8), .B(_13032_), .Y(_12915__57_) );
NOR2X1 NOR2X1_2051 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf7), .B(_13034_), .Y(_12915__58_) );
NOR2X1 NOR2X1_2052 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf6), .B(_13036_), .Y(_12915__59_) );
NOR2X1 NOR2X1_2053 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf5), .B(_13038_), .Y(_12915__60_) );
NOR2X1 NOR2X1_2054 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf4), .B(_13040_), .Y(_12915__61_) );
NOR2X1 NOR2X1_2055 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf3), .B(_13042_), .Y(_12915__62_) );
NOR2X1 NOR2X1_2056 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf2), .B(_13044_), .Y(_12915__63_) );
NOR2X1 NOR2X1_2057 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf1), .B(_13046_), .Y(_12915__64_) );
NOR2X1 NOR2X1_2058 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf0), .B(_13048_), .Y(_12915__65_) );
NOR2X1 NOR2X1_2059 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf42), .B(_13050_), .Y(_12915__66_) );
NOR2X1 NOR2X1_2060 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf41), .B(_13052_), .Y(_12915__67_) );
NOR2X1 NOR2X1_2061 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf40), .B(_13054_), .Y(_12915__68_) );
NOR2X1 NOR2X1_2062 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf39), .B(_13056_), .Y(_12915__69_) );
NOR2X1 NOR2X1_2063 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf38), .B(_13058_), .Y(_12915__70_) );
NOR2X1 NOR2X1_2064 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf37), .B(_13060_), .Y(_12915__71_) );
NOR2X1 NOR2X1_2065 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf36), .B(_13062_), .Y(_12915__72_) );
NOR2X1 NOR2X1_2066 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf35), .B(_13064_), .Y(_12915__73_) );
NOR2X1 NOR2X1_2067 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf34), .B(_13066_), .Y(_12915__74_) );
NOR2X1 NOR2X1_2068 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf33), .B(_13068_), .Y(_12915__75_) );
NOR2X1 NOR2X1_2069 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf32), .B(_13070_), .Y(_12915__76_) );
NOR2X1 NOR2X1_2070 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf31), .B(_13072_), .Y(_12915__77_) );
NOR2X1 NOR2X1_2071 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf30), .B(_13074_), .Y(_12915__78_) );
NOR2X1 NOR2X1_2072 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf29), .B(_13076_), .Y(_12915__79_) );
NOR2X1 NOR2X1_2073 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf28), .B(_13078_), .Y(_12915__80_) );
NOR2X1 NOR2X1_2074 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf27), .B(_13080_), .Y(_12915__81_) );
NOR2X1 NOR2X1_2075 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf26), .B(_13082_), .Y(_12915__82_) );
NOR2X1 NOR2X1_2076 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf25), .B(_13084_), .Y(_12915__83_) );
NOR2X1 NOR2X1_2077 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf24), .B(_13086_), .Y(_12915__84_) );
NOR2X1 NOR2X1_2078 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf23), .B(_13088_), .Y(_12915__85_) );
NOR2X1 NOR2X1_2079 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf22), .B(_13090_), .Y(_12915__86_) );
NOR2X1 NOR2X1_2080 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf21), .B(_13092_), .Y(_12915__87_) );
NOR2X1 NOR2X1_2081 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf20), .B(_13094_), .Y(_12915__88_) );
NOR2X1 NOR2X1_2082 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf19), .B(_13096_), .Y(_12915__89_) );
NOR2X1 NOR2X1_2083 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf18), .B(_13098_), .Y(_12915__90_) );
NOR2X1 NOR2X1_2084 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf17), .B(_13100_), .Y(_12915__91_) );
NOR2X1 NOR2X1_2085 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf16), .B(_13102_), .Y(_12915__92_) );
NOR2X1 NOR2X1_2086 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf15), .B(_13104_), .Y(_12915__93_) );
NOR2X1 NOR2X1_2087 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf14), .B(_13106_), .Y(_12915__94_) );
NOR2X1 NOR2X1_2088 ( .gnd(gnd), .vdd(vdd), .A(_12916__bF_buf13), .B(_13108_), .Y(_12915__95_) );
DFFPOSX1 DFFPOSX1_1570 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_12915__0_), .Q(concatenador_bloque_0_) );
DFFPOSX1 DFFPOSX1_1571 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_12915__1_), .Q(concatenador_bloque_1_) );
DFFPOSX1 DFFPOSX1_1572 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_12915__2_), .Q(concatenador_bloque_2_) );
DFFPOSX1 DFFPOSX1_1573 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_12915__3_), .Q(concatenador_bloque_3_) );
DFFPOSX1 DFFPOSX1_1574 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_12915__4_), .Q(concatenador_bloque_4_) );
DFFPOSX1 DFFPOSX1_1575 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_12915__5_), .Q(concatenador_bloque_5_) );
DFFPOSX1 DFFPOSX1_1576 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_12915__6_), .Q(concatenador_bloque_6_) );
DFFPOSX1 DFFPOSX1_1577 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_12915__7_), .Q(concatenador_bloque_7_) );
DFFPOSX1 DFFPOSX1_1578 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_12915__8_), .Q(concatenador_bloque_8_) );
DFFPOSX1 DFFPOSX1_1579 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_12915__9_), .Q(concatenador_bloque_9_) );
DFFPOSX1 DFFPOSX1_1580 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_12915__10_), .Q(concatenador_bloque_10_) );
DFFPOSX1 DFFPOSX1_1581 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf157), .D(_12915__11_), .Q(concatenador_bloque_11_) );
DFFPOSX1 DFFPOSX1_1582 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf156), .D(_12915__12_), .Q(concatenador_bloque_12_) );
DFFPOSX1 DFFPOSX1_1583 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf155), .D(_12915__13_), .Q(concatenador_bloque_13_) );
DFFPOSX1 DFFPOSX1_1584 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf154), .D(_12915__14_), .Q(concatenador_bloque_14_) );
DFFPOSX1 DFFPOSX1_1585 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf153), .D(_12915__15_), .Q(concatenador_bloque_15_) );
DFFPOSX1 DFFPOSX1_1586 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf152), .D(_12915__16_), .Q(concatenador_bloque_16_) );
DFFPOSX1 DFFPOSX1_1587 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf151), .D(_12915__17_), .Q(concatenador_bloque_17_) );
DFFPOSX1 DFFPOSX1_1588 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf150), .D(_12915__18_), .Q(concatenador_bloque_18_) );
DFFPOSX1 DFFPOSX1_1589 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf149), .D(_12915__19_), .Q(concatenador_bloque_19_) );
DFFPOSX1 DFFPOSX1_1590 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf148), .D(_12915__20_), .Q(concatenador_bloque_20_) );
DFFPOSX1 DFFPOSX1_1591 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf147), .D(_12915__21_), .Q(concatenador_bloque_21_) );
DFFPOSX1 DFFPOSX1_1592 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf146), .D(_12915__22_), .Q(concatenador_bloque_22_) );
DFFPOSX1 DFFPOSX1_1593 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf145), .D(_12915__23_), .Q(concatenador_bloque_23_) );
DFFPOSX1 DFFPOSX1_1594 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf144), .D(_12915__24_), .Q(concatenador_bloque_24_) );
DFFPOSX1 DFFPOSX1_1595 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf143), .D(_12915__25_), .Q(concatenador_bloque_25_) );
DFFPOSX1 DFFPOSX1_1596 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf142), .D(_12915__26_), .Q(concatenador_bloque_26_) );
DFFPOSX1 DFFPOSX1_1597 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf141), .D(_12915__27_), .Q(concatenador_bloque_27_) );
DFFPOSX1 DFFPOSX1_1598 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf140), .D(_12915__28_), .Q(concatenador_bloque_28_) );
DFFPOSX1 DFFPOSX1_1599 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf139), .D(_12915__29_), .Q(concatenador_bloque_29_) );
DFFPOSX1 DFFPOSX1_1600 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf138), .D(_12915__30_), .Q(concatenador_bloque_30_) );
DFFPOSX1 DFFPOSX1_1601 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf137), .D(_12915__31_), .Q(concatenador_bloque_31_) );
DFFPOSX1 DFFPOSX1_1602 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf136), .D(_12915__32_), .Q(concatenador_bloque_32_) );
DFFPOSX1 DFFPOSX1_1603 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf135), .D(_12915__33_), .Q(concatenador_bloque_33_) );
DFFPOSX1 DFFPOSX1_1604 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf134), .D(_12915__34_), .Q(concatenador_bloque_34_) );
DFFPOSX1 DFFPOSX1_1605 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf133), .D(_12915__35_), .Q(concatenador_bloque_35_) );
DFFPOSX1 DFFPOSX1_1606 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf132), .D(_12915__36_), .Q(concatenador_bloque_36_) );
DFFPOSX1 DFFPOSX1_1607 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf131), .D(_12915__37_), .Q(concatenador_bloque_37_) );
DFFPOSX1 DFFPOSX1_1608 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf130), .D(_12915__38_), .Q(concatenador_bloque_38_) );
DFFPOSX1 DFFPOSX1_1609 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf129), .D(_12915__39_), .Q(concatenador_bloque_39_) );
DFFPOSX1 DFFPOSX1_1610 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf128), .D(_12915__40_), .Q(concatenador_bloque_40_) );
DFFPOSX1 DFFPOSX1_1611 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf127), .D(_12915__41_), .Q(concatenador_bloque_41_) );
DFFPOSX1 DFFPOSX1_1612 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf126), .D(_12915__42_), .Q(concatenador_bloque_42_) );
DFFPOSX1 DFFPOSX1_1613 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf125), .D(_12915__43_), .Q(concatenador_bloque_43_) );
DFFPOSX1 DFFPOSX1_1614 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf124), .D(_12915__44_), .Q(concatenador_bloque_44_) );
DFFPOSX1 DFFPOSX1_1615 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf123), .D(_12915__45_), .Q(concatenador_bloque_45_) );
DFFPOSX1 DFFPOSX1_1616 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf122), .D(_12915__46_), .Q(concatenador_bloque_46_) );
DFFPOSX1 DFFPOSX1_1617 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf121), .D(_12915__47_), .Q(concatenador_bloque_47_) );
DFFPOSX1 DFFPOSX1_1618 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf120), .D(_12915__48_), .Q(concatenador_bloque_48_) );
DFFPOSX1 DFFPOSX1_1619 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf119), .D(_12915__49_), .Q(concatenador_bloque_49_) );
DFFPOSX1 DFFPOSX1_1620 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf118), .D(_12915__50_), .Q(concatenador_bloque_50_) );
DFFPOSX1 DFFPOSX1_1621 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf117), .D(_12915__51_), .Q(concatenador_bloque_51_) );
DFFPOSX1 DFFPOSX1_1622 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf116), .D(_12915__52_), .Q(concatenador_bloque_52_) );
DFFPOSX1 DFFPOSX1_1623 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf115), .D(_12915__53_), .Q(concatenador_bloque_53_) );
DFFPOSX1 DFFPOSX1_1624 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf114), .D(_12915__54_), .Q(concatenador_bloque_54_) );
DFFPOSX1 DFFPOSX1_1625 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf113), .D(_12915__55_), .Q(concatenador_bloque_55_) );
DFFPOSX1 DFFPOSX1_1626 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf112), .D(_12915__56_), .Q(concatenador_bloque_56_) );
DFFPOSX1 DFFPOSX1_1627 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf111), .D(_12915__57_), .Q(concatenador_bloque_57_) );
DFFPOSX1 DFFPOSX1_1628 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf110), .D(_12915__58_), .Q(concatenador_bloque_58_) );
DFFPOSX1 DFFPOSX1_1629 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf109), .D(_12915__59_), .Q(concatenador_bloque_59_) );
DFFPOSX1 DFFPOSX1_1630 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf108), .D(_12915__60_), .Q(concatenador_bloque_60_) );
DFFPOSX1 DFFPOSX1_1631 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf107), .D(_12915__61_), .Q(concatenador_bloque_61_) );
DFFPOSX1 DFFPOSX1_1632 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(_12915__62_), .Q(concatenador_bloque_62_) );
DFFPOSX1 DFFPOSX1_1633 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(_12915__63_), .Q(concatenador_bloque_63_) );
DFFPOSX1 DFFPOSX1_1634 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(_12915__64_), .Q(concatenador_bloque_64_) );
DFFPOSX1 DFFPOSX1_1635 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(_12915__65_), .Q(concatenador_bloque_65_) );
DFFPOSX1 DFFPOSX1_1636 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(_12915__66_), .Q(concatenador_bloque_66_) );
DFFPOSX1 DFFPOSX1_1637 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(_12915__67_), .Q(concatenador_bloque_67_) );
DFFPOSX1 DFFPOSX1_1638 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(_12915__68_), .Q(concatenador_bloque_68_) );
DFFPOSX1 DFFPOSX1_1639 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(_12915__69_), .Q(concatenador_bloque_69_) );
DFFPOSX1 DFFPOSX1_1640 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_12915__70_), .Q(concatenador_bloque_70_) );
DFFPOSX1 DFFPOSX1_1641 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_12915__71_), .Q(concatenador_bloque_71_) );
DFFPOSX1 DFFPOSX1_1642 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_12915__72_), .Q(concatenador_bloque_72_) );
DFFPOSX1 DFFPOSX1_1643 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_12915__73_), .Q(concatenador_bloque_73_) );
DFFPOSX1 DFFPOSX1_1644 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_12915__74_), .Q(concatenador_bloque_74_) );
DFFPOSX1 DFFPOSX1_1645 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_12915__75_), .Q(concatenador_bloque_75_) );
DFFPOSX1 DFFPOSX1_1646 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_12915__76_), .Q(concatenador_bloque_76_) );
DFFPOSX1 DFFPOSX1_1647 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_12915__77_), .Q(concatenador_bloque_77_) );
DFFPOSX1 DFFPOSX1_1648 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_12915__78_), .Q(concatenador_bloque_78_) );
DFFPOSX1 DFFPOSX1_1649 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_12915__79_), .Q(concatenador_bloque_79_) );
DFFPOSX1 DFFPOSX1_1650 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_12915__80_), .Q(concatenador_bloque_80_) );
DFFPOSX1 DFFPOSX1_1651 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_12915__81_), .Q(concatenador_bloque_81_) );
DFFPOSX1 DFFPOSX1_1652 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_12915__82_), .Q(concatenador_bloque_82_) );
DFFPOSX1 DFFPOSX1_1653 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_12915__83_), .Q(concatenador_bloque_83_) );
DFFPOSX1 DFFPOSX1_1654 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_12915__84_), .Q(concatenador_bloque_84_) );
DFFPOSX1 DFFPOSX1_1655 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_12915__85_), .Q(concatenador_bloque_85_) );
DFFPOSX1 DFFPOSX1_1656 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_12915__86_), .Q(concatenador_bloque_86_) );
DFFPOSX1 DFFPOSX1_1657 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_12915__87_), .Q(concatenador_bloque_87_) );
DFFPOSX1 DFFPOSX1_1658 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_12915__88_), .Q(concatenador_bloque_88_) );
DFFPOSX1 DFFPOSX1_1659 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_12915__89_), .Q(concatenador_bloque_89_) );
DFFPOSX1 DFFPOSX1_1660 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_12915__90_), .Q(concatenador_bloque_90_) );
DFFPOSX1 DFFPOSX1_1661 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_12915__91_), .Q(concatenador_bloque_91_) );
DFFPOSX1 DFFPOSX1_1662 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_12915__92_), .Q(concatenador_bloque_92_) );
DFFPOSX1 DFFPOSX1_1663 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_12915__93_), .Q(concatenador_bloque_93_) );
DFFPOSX1 DFFPOSX1_1664 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_12915__94_), .Q(concatenador_bloque_94_) );
DFFPOSX1 DFFPOSX1_1665 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_12915__95_), .Q(concatenador_bloque_95_) );
DFFPOSX1 DFFPOSX1_1666 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_12914__0_), .Q(next_b_data_in_prev_0_) );
DFFPOSX1 DFFPOSX1_1667 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_12914__1_), .Q(next_b_data_in_prev_1_) );
DFFPOSX1 DFFPOSX1_1668 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_12914__2_), .Q(next_b_data_in_prev_2_) );
DFFPOSX1 DFFPOSX1_1669 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_12914__3_), .Q(next_b_data_in_prev_3_) );
DFFPOSX1 DFFPOSX1_1670 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_12914__4_), .Q(next_b_data_in_prev_4_) );
DFFPOSX1 DFFPOSX1_1671 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_12914__5_), .Q(next_b_data_in_prev_5_) );
DFFPOSX1 DFFPOSX1_1672 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_12914__6_), .Q(next_b_data_in_prev_6_) );
DFFPOSX1 DFFPOSX1_1673 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_12914__7_), .Q(next_b_data_in_prev_7_) );
DFFPOSX1 DFFPOSX1_1674 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_12914__8_), .Q(next_b_data_in_prev_8_) );
DFFPOSX1 DFFPOSX1_1675 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_12914__9_), .Q(next_b_data_in_prev_9_) );
DFFPOSX1 DFFPOSX1_1676 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_12914__10_), .Q(next_b_data_in_prev_10_) );
DFFPOSX1 DFFPOSX1_1677 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_12914__11_), .Q(next_b_data_in_prev_11_) );
DFFPOSX1 DFFPOSX1_1678 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_12914__12_), .Q(next_b_data_in_prev_12_) );
DFFPOSX1 DFFPOSX1_1679 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_12914__13_), .Q(next_b_data_in_prev_13_) );
DFFPOSX1 DFFPOSX1_1680 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_12914__14_), .Q(next_b_data_in_prev_14_) );
DFFPOSX1 DFFPOSX1_1681 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_12914__15_), .Q(next_b_data_in_prev_15_) );
DFFPOSX1 DFFPOSX1_1682 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_12914__16_), .Q(next_b_data_in_prev_16_) );
DFFPOSX1 DFFPOSX1_1683 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_12914__17_), .Q(next_b_data_in_prev_17_) );
DFFPOSX1 DFFPOSX1_1684 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_12914__18_), .Q(next_b_data_in_prev_18_) );
DFFPOSX1 DFFPOSX1_1685 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_12914__19_), .Q(next_b_data_in_prev_19_) );
DFFPOSX1 DFFPOSX1_1686 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_12914__20_), .Q(next_b_data_in_prev_20_) );
DFFPOSX1 DFFPOSX1_1687 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_12914__21_), .Q(next_b_data_in_prev_21_) );
DFFPOSX1 DFFPOSX1_1688 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_12914__22_), .Q(next_b_data_in_prev_22_) );
DFFPOSX1 DFFPOSX1_1689 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_12914__23_), .Q(next_b_data_in_prev_23_) );
DFFPOSX1 DFFPOSX1_1690 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_12914__24_), .Q(next_b_data_in_prev_24_) );
DFFPOSX1 DFFPOSX1_1691 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_12914__25_), .Q(next_b_data_in_prev_25_) );
DFFPOSX1 DFFPOSX1_1692 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_12914__26_), .Q(next_b_data_in_prev_26_) );
DFFPOSX1 DFFPOSX1_1693 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_12914__27_), .Q(next_b_data_in_prev_27_) );
DFFPOSX1 DFFPOSX1_1694 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_12914__28_), .Q(next_b_data_in_prev_28_) );
DFFPOSX1 DFFPOSX1_1695 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_12914__29_), .Q(next_b_data_in_prev_29_) );
DFFPOSX1 DFFPOSX1_1696 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_12914__30_), .Q(next_b_data_in_prev_30_) );
DFFPOSX1 DFFPOSX1_1697 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_12914__31_), .Q(next_b_data_in_prev_31_) );
DFFPOSX1 DFFPOSX1_1698 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_12914__32_), .Q(next_b_data_in_prev_32_) );
DFFPOSX1 DFFPOSX1_1699 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_12914__33_), .Q(next_b_data_in_prev_33_) );
DFFPOSX1 DFFPOSX1_1700 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_12914__34_), .Q(next_b_data_in_prev_34_) );
DFFPOSX1 DFFPOSX1_1701 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_12914__35_), .Q(next_b_data_in_prev_35_) );
DFFPOSX1 DFFPOSX1_1702 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_12914__36_), .Q(next_b_data_in_prev_36_) );
DFFPOSX1 DFFPOSX1_1703 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_12914__37_), .Q(next_b_data_in_prev_37_) );
DFFPOSX1 DFFPOSX1_1704 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_12914__38_), .Q(next_b_data_in_prev_38_) );
DFFPOSX1 DFFPOSX1_1705 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_12914__39_), .Q(next_b_data_in_prev_39_) );
DFFPOSX1 DFFPOSX1_1706 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_12914__40_), .Q(next_b_data_in_prev_40_) );
DFFPOSX1 DFFPOSX1_1707 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_12914__41_), .Q(next_b_data_in_prev_41_) );
DFFPOSX1 DFFPOSX1_1708 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_12914__42_), .Q(next_b_data_in_prev_42_) );
DFFPOSX1 DFFPOSX1_1709 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_12914__43_), .Q(next_b_data_in_prev_43_) );
DFFPOSX1 DFFPOSX1_1710 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_12914__44_), .Q(next_b_data_in_prev_44_) );
DFFPOSX1 DFFPOSX1_1711 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_12914__45_), .Q(next_b_data_in_prev_45_) );
DFFPOSX1 DFFPOSX1_1712 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_12914__46_), .Q(next_b_data_in_prev_46_) );
DFFPOSX1 DFFPOSX1_1713 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_12914__47_), .Q(next_b_data_in_prev_47_) );
DFFPOSX1 DFFPOSX1_1714 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_12914__48_), .Q(next_b_data_in_prev_48_) );
DFFPOSX1 DFFPOSX1_1715 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_12914__49_), .Q(next_b_data_in_prev_49_) );
DFFPOSX1 DFFPOSX1_1716 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_12914__50_), .Q(next_b_data_in_prev_50_) );
DFFPOSX1 DFFPOSX1_1717 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_12914__51_), .Q(next_b_data_in_prev_51_) );
DFFPOSX1 DFFPOSX1_1718 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_12914__52_), .Q(next_b_data_in_prev_52_) );
DFFPOSX1 DFFPOSX1_1719 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_12914__53_), .Q(next_b_data_in_prev_53_) );
DFFPOSX1 DFFPOSX1_1720 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_12914__54_), .Q(next_b_data_in_prev_54_) );
DFFPOSX1 DFFPOSX1_1721 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_12914__55_), .Q(next_b_data_in_prev_55_) );
DFFPOSX1 DFFPOSX1_1722 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_12914__56_), .Q(next_b_data_in_prev_56_) );
DFFPOSX1 DFFPOSX1_1723 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_12914__57_), .Q(next_b_data_in_prev_57_) );
DFFPOSX1 DFFPOSX1_1724 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_12914__58_), .Q(next_b_data_in_prev_58_) );
DFFPOSX1 DFFPOSX1_1725 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_12914__59_), .Q(next_b_data_in_prev_59_) );
DFFPOSX1 DFFPOSX1_1726 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_12914__60_), .Q(next_b_data_in_prev_60_) );
DFFPOSX1 DFFPOSX1_1727 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_12914__61_), .Q(next_b_data_in_prev_61_) );
DFFPOSX1 DFFPOSX1_1728 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_12914__62_), .Q(next_b_data_in_prev_62_) );
DFFPOSX1 DFFPOSX1_1729 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_12914__63_), .Q(next_b_data_in_prev_63_) );
DFFPOSX1 DFFPOSX1_1730 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_12914__64_), .Q(next_b_data_in_prev_64_) );
DFFPOSX1 DFFPOSX1_1731 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_12914__65_), .Q(next_b_data_in_prev_65_) );
DFFPOSX1 DFFPOSX1_1732 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_12914__66_), .Q(next_b_data_in_prev_66_) );
DFFPOSX1 DFFPOSX1_1733 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_12914__67_), .Q(next_b_data_in_prev_67_) );
DFFPOSX1 DFFPOSX1_1734 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_12914__68_), .Q(next_b_data_in_prev_68_) );
DFFPOSX1 DFFPOSX1_1735 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_12914__69_), .Q(next_b_data_in_prev_69_) );
DFFPOSX1 DFFPOSX1_1736 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_12914__70_), .Q(next_b_data_in_prev_70_) );
DFFPOSX1 DFFPOSX1_1737 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_12914__71_), .Q(next_b_data_in_prev_71_) );
DFFPOSX1 DFFPOSX1_1738 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_12914__72_), .Q(next_b_data_in_prev_72_) );
DFFPOSX1 DFFPOSX1_1739 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf157), .D(_12914__73_), .Q(next_b_data_in_prev_73_) );
DFFPOSX1 DFFPOSX1_1740 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf156), .D(_12914__74_), .Q(next_b_data_in_prev_74_) );
DFFPOSX1 DFFPOSX1_1741 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf155), .D(_12914__75_), .Q(next_b_data_in_prev_75_) );
DFFPOSX1 DFFPOSX1_1742 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf154), .D(_12914__76_), .Q(next_b_data_in_prev_76_) );
DFFPOSX1 DFFPOSX1_1743 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf153), .D(_12914__77_), .Q(next_b_data_in_prev_77_) );
DFFPOSX1 DFFPOSX1_1744 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf152), .D(_12914__78_), .Q(next_b_data_in_prev_78_) );
DFFPOSX1 DFFPOSX1_1745 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf151), .D(_12914__79_), .Q(next_b_data_in_prev_79_) );
DFFPOSX1 DFFPOSX1_1746 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf150), .D(_12914__80_), .Q(next_b_data_in_prev_80_) );
DFFPOSX1 DFFPOSX1_1747 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf149), .D(_12914__81_), .Q(next_b_data_in_prev_81_) );
DFFPOSX1 DFFPOSX1_1748 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf148), .D(_12914__82_), .Q(next_b_data_in_prev_82_) );
DFFPOSX1 DFFPOSX1_1749 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf147), .D(_12914__83_), .Q(next_b_data_in_prev_83_) );
DFFPOSX1 DFFPOSX1_1750 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf146), .D(_12914__84_), .Q(next_b_data_in_prev_84_) );
DFFPOSX1 DFFPOSX1_1751 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf145), .D(_12914__85_), .Q(next_b_data_in_prev_85_) );
DFFPOSX1 DFFPOSX1_1752 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf144), .D(_12914__86_), .Q(next_b_data_in_prev_86_) );
DFFPOSX1 DFFPOSX1_1753 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf143), .D(_12914__87_), .Q(next_b_data_in_prev_87_) );
DFFPOSX1 DFFPOSX1_1754 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf142), .D(_12914__88_), .Q(next_b_data_in_prev_88_) );
DFFPOSX1 DFFPOSX1_1755 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf141), .D(_12914__89_), .Q(next_b_data_in_prev_89_) );
DFFPOSX1 DFFPOSX1_1756 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf140), .D(_12914__90_), .Q(next_b_data_in_prev_90_) );
DFFPOSX1 DFFPOSX1_1757 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf139), .D(_12914__91_), .Q(next_b_data_in_prev_91_) );
DFFPOSX1 DFFPOSX1_1758 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf138), .D(_12914__92_), .Q(next_b_data_in_prev_92_) );
DFFPOSX1 DFFPOSX1_1759 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf137), .D(_12914__93_), .Q(next_b_data_in_prev_93_) );
DFFPOSX1 DFFPOSX1_1760 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf136), .D(_12914__94_), .Q(next_b_data_in_prev_94_) );
DFFPOSX1 DFFPOSX1_1761 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf135), .D(_12914__95_), .Q(next_b_data_in_prev_95_) );
INVX1 INVX1_845 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf3), .Y(_13216_) );
NOR2X1 NOR2X1_2089 ( .gnd(gnd), .vdd(vdd), .A(_0__bF_buf9), .B(_13216_), .Y(_13217_) );
INVX4 INVX4_155 ( .gnd(gnd), .vdd(vdd), .A(_13217__bF_buf4), .Y(_13218_) );
INVX1 INVX1_846 ( .gnd(gnd), .vdd(vdd), .A(comparador_next_bF_buf0), .Y(_13219_) );
NOR2X1 NOR2X1_2090 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_0_), .B(_13219_), .Y(_13220_) );
INVX1 INVX1_847 ( .gnd(gnd), .vdd(vdd), .A(_13220_), .Y(_13221_) );
NAND2X1 NAND2X1_1793 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_0_), .B(_13219_), .Y(_13222_) );
AOI21X1 AOI21X1_2252 ( .gnd(gnd), .vdd(vdd), .A(_13222_), .B(_13221_), .C(_13218_), .Y(_13109__0_) );
OAI21X1 OAI21X1_3759 ( .gnd(gnd), .vdd(vdd), .A(_13220_), .B(concatenador_nonce_1_), .C(_13217__bF_buf3), .Y(_13223_) );
AOI21X1 AOI21X1_2253 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_1_), .B(_13220_), .C(_13223_), .Y(_13109__1_) );
OAI21X1 OAI21X1_3760 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_0_), .B(concatenador_nonce_1_), .C(comparador_next_bF_buf3), .Y(_13224_) );
INVX1 INVX1_848 ( .gnd(gnd), .vdd(vdd), .A(_13224_), .Y(_13225_) );
AND2X2 AND2X2_764 ( .gnd(gnd), .vdd(vdd), .A(_13225_), .B(concatenador_nonce_2_), .Y(_13226_) );
OAI21X1 OAI21X1_3761 ( .gnd(gnd), .vdd(vdd), .A(_13225_), .B(concatenador_nonce_2_), .C(_13217__bF_buf2), .Y(_13227_) );
NOR2X1 NOR2X1_2091 ( .gnd(gnd), .vdd(vdd), .A(_13227_), .B(_13226_), .Y(_13109__2_) );
NOR2X1 NOR2X1_2092 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_3_), .B(_13226_), .Y(_13228_) );
NAND2X1 NAND2X1_1794 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_2_), .B(concatenador_nonce_3_), .Y(_13229_) );
OAI21X1 OAI21X1_3762 ( .gnd(gnd), .vdd(vdd), .A(_13224_), .B(_13229_), .C(_13217__bF_buf1), .Y(_13230_) );
NOR2X1 NOR2X1_2093 ( .gnd(gnd), .vdd(vdd), .A(_13230_), .B(_13228_), .Y(_13109__3_) );
NOR2X1 NOR2X1_2094 ( .gnd(gnd), .vdd(vdd), .A(_13229_), .B(_13224_), .Y(_13231_) );
AND2X2 AND2X2_765 ( .gnd(gnd), .vdd(vdd), .A(_13231_), .B(concatenador_nonce_4_), .Y(_13232_) );
OAI21X1 OAI21X1_3763 ( .gnd(gnd), .vdd(vdd), .A(_13231_), .B(concatenador_nonce_4_), .C(_13217__bF_buf0), .Y(_13233_) );
NOR2X1 NOR2X1_2095 ( .gnd(gnd), .vdd(vdd), .A(_13233_), .B(_13232_), .Y(_13109__4_) );
AND2X2 AND2X2_766 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_2_), .B(concatenador_nonce_3_), .Y(_13234_) );
NAND3X1 NAND3X1_660 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_4_), .B(concatenador_nonce_5_), .C(_13234_), .Y(_13235_) );
NOR2X1 NOR2X1_2096 ( .gnd(gnd), .vdd(vdd), .A(_13224_), .B(_13235_), .Y(_13236_) );
OAI21X1 OAI21X1_3764 ( .gnd(gnd), .vdd(vdd), .A(_13232_), .B(concatenador_nonce_5_), .C(_13217__bF_buf4), .Y(_13237_) );
NOR2X1 NOR2X1_2097 ( .gnd(gnd), .vdd(vdd), .A(_13236_), .B(_13237_), .Y(_13109__5_) );
AND2X2 AND2X2_767 ( .gnd(gnd), .vdd(vdd), .A(_13236_), .B(concatenador_nonce_6_), .Y(_13238_) );
OAI21X1 OAI21X1_3765 ( .gnd(gnd), .vdd(vdd), .A(_13236_), .B(concatenador_nonce_6_), .C(_13217__bF_buf3), .Y(_13239_) );
NOR2X1 NOR2X1_2098 ( .gnd(gnd), .vdd(vdd), .A(_13239_), .B(_13238_), .Y(_13109__6_) );
NOR2X1 NOR2X1_2099 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_7_), .B(_13238_), .Y(_13240_) );
AND2X2 AND2X2_768 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_6_), .B(concatenador_nonce_7_), .Y(_13110_) );
NAND2X1 NAND2X1_1795 ( .gnd(gnd), .vdd(vdd), .A(_13110_), .B(_13236_), .Y(_13111_) );
NAND2X1 NAND2X1_1796 ( .gnd(gnd), .vdd(vdd), .A(_13217__bF_buf2), .B(_13111_), .Y(_13112_) );
NOR2X1 NOR2X1_2100 ( .gnd(gnd), .vdd(vdd), .A(_13112_), .B(_13240_), .Y(_13109__7_) );
INVX1 INVX1_849 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_8_), .Y(_13113_) );
OR2X2 OR2X2_79 ( .gnd(gnd), .vdd(vdd), .A(_13111_), .B(_13113_), .Y(_13114_) );
AOI21X1 AOI21X1_2254 ( .gnd(gnd), .vdd(vdd), .A(_13113_), .B(_13111_), .C(_13218_), .Y(_13115_) );
AND2X2 AND2X2_769 ( .gnd(gnd), .vdd(vdd), .A(_13114_), .B(_13115_), .Y(_13109__8_) );
INVX1 INVX1_850 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_9_), .Y(_13116_) );
NAND2X1 NAND2X1_1797 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_8_), .B(concatenador_nonce_9_), .Y(_13117_) );
OAI21X1 OAI21X1_3766 ( .gnd(gnd), .vdd(vdd), .A(_13111_), .B(_13117_), .C(_13217__bF_buf1), .Y(_13118_) );
AOI21X1 AOI21X1_2255 ( .gnd(gnd), .vdd(vdd), .A(_13116_), .B(_13114_), .C(_13118_), .Y(_13109__9_) );
OAI21X1 OAI21X1_3767 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_0_), .B(concatenador_nonce_1_), .C(_13234_), .Y(_13119_) );
NAND3X1 NAND3X1_661 ( .gnd(gnd), .vdd(vdd), .A(comparador_next_bF_buf2), .B(concatenador_nonce_4_), .C(concatenador_nonce_5_), .Y(_13120_) );
AND2X2 AND2X2_770 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_8_), .B(concatenador_nonce_9_), .Y(_13121_) );
NAND2X1 NAND2X1_1798 ( .gnd(gnd), .vdd(vdd), .A(_13110_), .B(_13121_), .Y(_13122_) );
NOR3X1 NOR3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_13122_), .B(_13120_), .C(_13119_), .Y(_13123_) );
OAI21X1 OAI21X1_3768 ( .gnd(gnd), .vdd(vdd), .A(_13123_), .B(concatenador_nonce_10_), .C(_13217__bF_buf0), .Y(_13124_) );
AOI21X1 AOI21X1_2256 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_10_), .B(_13123_), .C(_13124_), .Y(_13109__10_) );
AOI21X1 AOI21X1_2257 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_10_), .B(_13123_), .C(concatenador_nonce_11_), .Y(_13125_) );
NOR2X1 NOR2X1_2101 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_0_), .B(concatenador_nonce_1_), .Y(_13126_) );
NOR2X1 NOR2X1_2102 ( .gnd(gnd), .vdd(vdd), .A(_13229_), .B(_13126_), .Y(_13127_) );
INVX1 INVX1_851 ( .gnd(gnd), .vdd(vdd), .A(_13120_), .Y(_13128_) );
NAND2X1 NAND2X1_1799 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_6_), .B(concatenador_nonce_7_), .Y(_13129_) );
NOR2X1 NOR2X1_2103 ( .gnd(gnd), .vdd(vdd), .A(_13129_), .B(_13117_), .Y(_13130_) );
NAND3X1 NAND3X1_662 ( .gnd(gnd), .vdd(vdd), .A(_13128_), .B(_13130_), .C(_13127_), .Y(_13131_) );
NAND2X1 NAND2X1_1800 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_10_), .B(concatenador_nonce_11_), .Y(_13132_) );
OAI21X1 OAI21X1_3769 ( .gnd(gnd), .vdd(vdd), .A(_13131_), .B(_13132_), .C(_13217__bF_buf4), .Y(_13133_) );
NOR2X1 NOR2X1_2104 ( .gnd(gnd), .vdd(vdd), .A(_13133_), .B(_13125_), .Y(_13109__11_) );
NOR2X1 NOR2X1_2105 ( .gnd(gnd), .vdd(vdd), .A(_13132_), .B(_13131_), .Y(_13134_) );
OAI21X1 OAI21X1_3770 ( .gnd(gnd), .vdd(vdd), .A(_13134_), .B(concatenador_nonce_12_), .C(_13217__bF_buf3), .Y(_13135_) );
AND2X2 AND2X2_771 ( .gnd(gnd), .vdd(vdd), .A(_13134_), .B(concatenador_nonce_12_), .Y(_13136_) );
NOR2X1 NOR2X1_2106 ( .gnd(gnd), .vdd(vdd), .A(_13135_), .B(_13136_), .Y(_13109__12_) );
OAI21X1 OAI21X1_3771 ( .gnd(gnd), .vdd(vdd), .A(_13136_), .B(concatenador_nonce_13_), .C(_13217__bF_buf2), .Y(_13137_) );
AOI21X1 AOI21X1_2258 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_13_), .B(_13136_), .C(_13137_), .Y(_13109__13_) );
OR2X2 OR2X2_80 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_0_), .B(concatenador_nonce_1_), .Y(_13138_) );
NAND3X1 NAND3X1_663 ( .gnd(gnd), .vdd(vdd), .A(_13110_), .B(_13121_), .C(_13138_), .Y(_13139_) );
NOR2X1 NOR2X1_2107 ( .gnd(gnd), .vdd(vdd), .A(_13235_), .B(_13139_), .Y(_13140_) );
NAND2X1 NAND2X1_1801 ( .gnd(gnd), .vdd(vdd), .A(comparador_next_bF_buf1), .B(_13140_), .Y(_13141_) );
NAND2X1 NAND2X1_1802 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_12_), .B(concatenador_nonce_13_), .Y(_13142_) );
NOR2X1 NOR2X1_2108 ( .gnd(gnd), .vdd(vdd), .A(_13132_), .B(_13142_), .Y(_13143_) );
INVX1 INVX1_852 ( .gnd(gnd), .vdd(vdd), .A(_13143_), .Y(_13144_) );
NOR2X1 NOR2X1_2109 ( .gnd(gnd), .vdd(vdd), .A(_13144_), .B(_13141_), .Y(_13145_) );
OAI21X1 OAI21X1_3772 ( .gnd(gnd), .vdd(vdd), .A(_13145_), .B(concatenador_nonce_14_), .C(_13217__bF_buf1), .Y(_13146_) );
AOI21X1 AOI21X1_2259 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_14_), .B(_13145_), .C(_13146_), .Y(_13109__14_) );
NAND3X1 NAND3X1_664 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_14_), .B(concatenador_nonce_15_), .C(_13143_), .Y(_13147_) );
NOR2X1 NOR2X1_2110 ( .gnd(gnd), .vdd(vdd), .A(_13147_), .B(_13141_), .Y(_13148_) );
AOI21X1 AOI21X1_2260 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_14_), .B(_13145_), .C(concatenador_nonce_15_), .Y(_13149_) );
NOR3X1 NOR3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_13218_), .B(_13148_), .C(_13149_), .Y(_13109__15_) );
OAI21X1 OAI21X1_3773 ( .gnd(gnd), .vdd(vdd), .A(_13148_), .B(concatenador_nonce_16_), .C(_13217__bF_buf0), .Y(_13150_) );
AOI21X1 AOI21X1_2261 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_16_), .B(_13148_), .C(_13150_), .Y(_13109__16_) );
AND2X2 AND2X2_772 ( .gnd(gnd), .vdd(vdd), .A(_13140_), .B(comparador_next_bF_buf0), .Y(_13151_) );
NAND2X1 NAND2X1_1803 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_16_), .B(concatenador_nonce_17_), .Y(_13152_) );
NOR2X1 NOR2X1_2111 ( .gnd(gnd), .vdd(vdd), .A(_13152_), .B(_13147_), .Y(_13153_) );
AND2X2 AND2X2_773 ( .gnd(gnd), .vdd(vdd), .A(_13151_), .B(_13153_), .Y(_13154_) );
AOI21X1 AOI21X1_2262 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_16_), .B(_13148_), .C(concatenador_nonce_17_), .Y(_13155_) );
NOR3X1 NOR3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_13218_), .B(_13154_), .C(_13155_), .Y(_13109__17_) );
OAI21X1 OAI21X1_3774 ( .gnd(gnd), .vdd(vdd), .A(_13154_), .B(concatenador_nonce_18_), .C(_13217__bF_buf4), .Y(_13156_) );
AOI21X1 AOI21X1_2263 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_18_), .B(_13154_), .C(_13156_), .Y(_13109__18_) );
NAND3X1 NAND3X1_665 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_18_), .B(_13153_), .C(_13151_), .Y(_13157_) );
NAND2X1 NAND2X1_1804 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_19_), .B(_13157_), .Y(_13158_) );
OR2X2 OR2X2_81 ( .gnd(gnd), .vdd(vdd), .A(_13157_), .B(concatenador_nonce_19_), .Y(_13159_) );
AOI21X1 AOI21X1_2264 ( .gnd(gnd), .vdd(vdd), .A(_13158_), .B(_13159_), .C(_13218_), .Y(_13109__19_) );
INVX1 INVX1_853 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_20_), .Y(_13160_) );
NAND3X1 NAND3X1_666 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_13_), .B(concatenador_nonce_14_), .C(concatenador_nonce_15_), .Y(_13161_) );
NOR2X1 NOR2X1_2112 ( .gnd(gnd), .vdd(vdd), .A(_13152_), .B(_13161_), .Y(_13162_) );
NAND3X1 NAND3X1_667 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_12_), .B(concatenador_nonce_18_), .C(concatenador_nonce_19_), .Y(_13163_) );
NOR2X1 NOR2X1_2113 ( .gnd(gnd), .vdd(vdd), .A(_13132_), .B(_13163_), .Y(_13164_) );
NAND2X1 NAND2X1_1805 ( .gnd(gnd), .vdd(vdd), .A(_13162_), .B(_13164_), .Y(_13165_) );
OAI21X1 OAI21X1_3775 ( .gnd(gnd), .vdd(vdd), .A(_13131_), .B(_13165_), .C(_13160_), .Y(_13166_) );
NAND2X1 NAND2X1_1806 ( .gnd(gnd), .vdd(vdd), .A(_13217__bF_buf3), .B(_13166_), .Y(_13167_) );
AND2X2 AND2X2_774 ( .gnd(gnd), .vdd(vdd), .A(_13162_), .B(_13164_), .Y(_13168_) );
NAND2X1 NAND2X1_1807 ( .gnd(gnd), .vdd(vdd), .A(_13168_), .B(_13123_), .Y(_13169_) );
NOR2X1 NOR2X1_2114 ( .gnd(gnd), .vdd(vdd), .A(_13160_), .B(_13169_), .Y(_13170_) );
NOR2X1 NOR2X1_2115 ( .gnd(gnd), .vdd(vdd), .A(_13167_), .B(_13170_), .Y(_13109__20_) );
NOR2X1 NOR2X1_2116 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_21_), .B(_13170_), .Y(_13171_) );
NAND2X1 NAND2X1_1808 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_20_), .B(concatenador_nonce_21_), .Y(_13172_) );
OAI21X1 OAI21X1_3776 ( .gnd(gnd), .vdd(vdd), .A(_13169_), .B(_13172_), .C(_13217__bF_buf2), .Y(_13173_) );
NOR2X1 NOR2X1_2117 ( .gnd(gnd), .vdd(vdd), .A(_13173_), .B(_13171_), .Y(_13109__21_) );
NOR3X1 NOR3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_13165_), .B(_13172_), .C(_13131_), .Y(_13174_) );
OAI21X1 OAI21X1_3777 ( .gnd(gnd), .vdd(vdd), .A(_13174_), .B(concatenador_nonce_22_), .C(_13217__bF_buf1), .Y(_13175_) );
INVX2 INVX2_393 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_22_), .Y(_13176_) );
INVX1 INVX1_854 ( .gnd(gnd), .vdd(vdd), .A(_13172_), .Y(_13177_) );
NAND3X1 NAND3X1_668 ( .gnd(gnd), .vdd(vdd), .A(_13168_), .B(_13177_), .C(_13123_), .Y(_13178_) );
NOR2X1 NOR2X1_2118 ( .gnd(gnd), .vdd(vdd), .A(_13176_), .B(_13178_), .Y(_13179_) );
NOR2X1 NOR2X1_2119 ( .gnd(gnd), .vdd(vdd), .A(_13179_), .B(_13175_), .Y(_13109__22_) );
INVX1 INVX1_855 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_23_), .Y(_13180_) );
NOR3X1 NOR3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_13176_), .B(_13180_), .C(_13178_), .Y(_13181_) );
OAI21X1 OAI21X1_3778 ( .gnd(gnd), .vdd(vdd), .A(_13179_), .B(concatenador_nonce_23_), .C(_13217__bF_buf0), .Y(_13182_) );
NOR2X1 NOR2X1_2120 ( .gnd(gnd), .vdd(vdd), .A(_13181_), .B(_13182_), .Y(_13109__23_) );
OAI21X1 OAI21X1_3779 ( .gnd(gnd), .vdd(vdd), .A(_13181_), .B(concatenador_nonce_24_), .C(_13217__bF_buf4), .Y(_13183_) );
AOI21X1 AOI21X1_2265 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_24_), .B(_13181_), .C(_13183_), .Y(_13109__24_) );
INVX1 INVX1_856 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_24_), .Y(_13184_) );
NAND3X1 NAND3X1_669 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_22_), .B(concatenador_nonce_23_), .C(_13174_), .Y(_13185_) );
OAI21X1 OAI21X1_3780 ( .gnd(gnd), .vdd(vdd), .A(_13185_), .B(_13184_), .C(concatenador_nonce_25_), .Y(_13186_) );
INVX1 INVX1_857 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_25_), .Y(_13187_) );
NAND3X1 NAND3X1_670 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_24_), .B(_13187_), .C(_13181_), .Y(_13188_) );
AOI21X1 AOI21X1_2266 ( .gnd(gnd), .vdd(vdd), .A(_13186_), .B(_13188_), .C(_13218_), .Y(_13109__25_) );
NAND3X1 NAND3X1_671 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_23_), .B(concatenador_nonce_24_), .C(concatenador_nonce_25_), .Y(_13189_) );
NOR3X1 NOR3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_13176_), .B(_13189_), .C(_13178_), .Y(_13190_) );
OAI21X1 OAI21X1_3781 ( .gnd(gnd), .vdd(vdd), .A(_13190_), .B(concatenador_nonce_26_), .C(_13217__bF_buf3), .Y(_13191_) );
AOI21X1 AOI21X1_2267 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_26_), .B(_13190_), .C(_13191_), .Y(_13109__26_) );
INVX1 INVX1_858 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_26_), .Y(_13192_) );
INVX1 INVX1_859 ( .gnd(gnd), .vdd(vdd), .A(_13189_), .Y(_13193_) );
NAND3X1 NAND3X1_672 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_22_), .B(_13193_), .C(_13174_), .Y(_13194_) );
OAI21X1 OAI21X1_3782 ( .gnd(gnd), .vdd(vdd), .A(_13194_), .B(_13192_), .C(concatenador_nonce_27_), .Y(_13195_) );
INVX1 INVX1_860 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_27_), .Y(_13196_) );
NAND3X1 NAND3X1_673 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_26_), .B(_13196_), .C(_13190_), .Y(_13197_) );
AOI21X1 AOI21X1_2268 ( .gnd(gnd), .vdd(vdd), .A(_13195_), .B(_13197_), .C(_13218_), .Y(_13109__27_) );
NAND3X1 NAND3X1_674 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_22_), .B(concatenador_nonce_26_), .C(concatenador_nonce_27_), .Y(_13198_) );
NOR2X1 NOR2X1_2121 ( .gnd(gnd), .vdd(vdd), .A(_13172_), .B(_13198_), .Y(_13199_) );
NAND2X1 NAND2X1_1809 ( .gnd(gnd), .vdd(vdd), .A(_13193_), .B(_13199_), .Y(_13200_) );
NOR3X1 NOR3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_13165_), .B(_13200_), .C(_13131_), .Y(_13201_) );
OAI21X1 OAI21X1_3783 ( .gnd(gnd), .vdd(vdd), .A(_13201_), .B(concatenador_nonce_28_), .C(_13217__bF_buf2), .Y(_13202_) );
INVX1 INVX1_861 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_28_), .Y(_13203_) );
AND2X2 AND2X2_775 ( .gnd(gnd), .vdd(vdd), .A(_13199_), .B(_13193_), .Y(_13204_) );
NAND3X1 NAND3X1_675 ( .gnd(gnd), .vdd(vdd), .A(_13168_), .B(_13204_), .C(_13123_), .Y(_13205_) );
NOR2X1 NOR2X1_2122 ( .gnd(gnd), .vdd(vdd), .A(_13203_), .B(_13205_), .Y(_13206_) );
NOR2X1 NOR2X1_2123 ( .gnd(gnd), .vdd(vdd), .A(_13206_), .B(_13202_), .Y(_13109__28_) );
INVX1 INVX1_862 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_29_), .Y(_13207_) );
NOR3X1 NOR3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_13203_), .B(_13207_), .C(_13205_), .Y(_13208_) );
OAI21X1 OAI21X1_3784 ( .gnd(gnd), .vdd(vdd), .A(_13206_), .B(concatenador_nonce_29_), .C(_13217__bF_buf1), .Y(_13209_) );
NOR2X1 NOR2X1_2124 ( .gnd(gnd), .vdd(vdd), .A(_13208_), .B(_13209_), .Y(_13109__29_) );
OAI21X1 OAI21X1_3785 ( .gnd(gnd), .vdd(vdd), .A(_13208_), .B(concatenador_nonce_30_), .C(_13217__bF_buf0), .Y(_13210_) );
AOI21X1 AOI21X1_2269 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_30_), .B(_13208_), .C(_13210_), .Y(_13109__30_) );
INVX1 INVX1_863 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_30_), .Y(_13211_) );
NAND3X1 NAND3X1_676 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_28_), .B(concatenador_nonce_29_), .C(_13201_), .Y(_13212_) );
OAI21X1 OAI21X1_3786 ( .gnd(gnd), .vdd(vdd), .A(_13212_), .B(_13211_), .C(concatenador_nonce_31_), .Y(_13213_) );
INVX1 INVX1_864 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_31_), .Y(_13214_) );
NAND3X1 NAND3X1_677 ( .gnd(gnd), .vdd(vdd), .A(concatenador_nonce_30_), .B(_13214_), .C(_13208_), .Y(_13215_) );
AOI21X1 AOI21X1_2270 ( .gnd(gnd), .vdd(vdd), .A(_13213_), .B(_13215_), .C(_13218_), .Y(_13109__31_) );
DFFPOSX1 DFFPOSX1_1762 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf134), .D(_13109__0_), .Q(concatenador_nonce_0_) );
DFFPOSX1 DFFPOSX1_1763 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf133), .D(_13109__1_), .Q(concatenador_nonce_1_) );
DFFPOSX1 DFFPOSX1_1764 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf132), .D(_13109__2_), .Q(concatenador_nonce_2_) );
DFFPOSX1 DFFPOSX1_1765 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf131), .D(_13109__3_), .Q(concatenador_nonce_3_) );
DFFPOSX1 DFFPOSX1_1766 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf130), .D(_13109__4_), .Q(concatenador_nonce_4_) );
DFFPOSX1 DFFPOSX1_1767 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf129), .D(_13109__5_), .Q(concatenador_nonce_5_) );
DFFPOSX1 DFFPOSX1_1768 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf128), .D(_13109__6_), .Q(concatenador_nonce_6_) );
DFFPOSX1 DFFPOSX1_1769 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf127), .D(_13109__7_), .Q(concatenador_nonce_7_) );
DFFPOSX1 DFFPOSX1_1770 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf126), .D(_13109__8_), .Q(concatenador_nonce_8_) );
DFFPOSX1 DFFPOSX1_1771 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf125), .D(_13109__9_), .Q(concatenador_nonce_9_) );
DFFPOSX1 DFFPOSX1_1772 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf124), .D(_13109__10_), .Q(concatenador_nonce_10_) );
DFFPOSX1 DFFPOSX1_1773 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf123), .D(_13109__11_), .Q(concatenador_nonce_11_) );
DFFPOSX1 DFFPOSX1_1774 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf122), .D(_13109__12_), .Q(concatenador_nonce_12_) );
DFFPOSX1 DFFPOSX1_1775 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf121), .D(_13109__13_), .Q(concatenador_nonce_13_) );
DFFPOSX1 DFFPOSX1_1776 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf120), .D(_13109__14_), .Q(concatenador_nonce_14_) );
DFFPOSX1 DFFPOSX1_1777 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf119), .D(_13109__15_), .Q(concatenador_nonce_15_) );
DFFPOSX1 DFFPOSX1_1778 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf118), .D(_13109__16_), .Q(concatenador_nonce_16_) );
DFFPOSX1 DFFPOSX1_1779 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf117), .D(_13109__17_), .Q(concatenador_nonce_17_) );
DFFPOSX1 DFFPOSX1_1780 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf116), .D(_13109__18_), .Q(concatenador_nonce_18_) );
DFFPOSX1 DFFPOSX1_1781 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf115), .D(_13109__19_), .Q(concatenador_nonce_19_) );
DFFPOSX1 DFFPOSX1_1782 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf114), .D(_13109__20_), .Q(concatenador_nonce_20_) );
DFFPOSX1 DFFPOSX1_1783 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf113), .D(_13109__21_), .Q(concatenador_nonce_21_) );
DFFPOSX1 DFFPOSX1_1784 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf112), .D(_13109__22_), .Q(concatenador_nonce_22_) );
DFFPOSX1 DFFPOSX1_1785 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf111), .D(_13109__23_), .Q(concatenador_nonce_23_) );
DFFPOSX1 DFFPOSX1_1786 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf110), .D(_13109__24_), .Q(concatenador_nonce_24_) );
DFFPOSX1 DFFPOSX1_1787 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf109), .D(_13109__25_), .Q(concatenador_nonce_25_) );
DFFPOSX1 DFFPOSX1_1788 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf108), .D(_13109__26_), .Q(concatenador_nonce_26_) );
DFFPOSX1 DFFPOSX1_1789 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf107), .D(_13109__27_), .Q(concatenador_nonce_27_) );
DFFPOSX1 DFFPOSX1_1790 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(_13109__28_), .Q(concatenador_nonce_28_) );
DFFPOSX1 DFFPOSX1_1791 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(_13109__29_), .Q(concatenador_nonce_29_) );
DFFPOSX1 DFFPOSX1_1792 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(_13109__30_), .Q(concatenador_nonce_30_) );
DFFPOSX1 DFFPOSX1_1793 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(_13109__31_), .Q(concatenador_nonce_31_) );
INVX1 INVX1_865 ( .gnd(gnd), .vdd(vdd), .A(comparador_next_bF_buf3), .Y(_13352_) );
NOR2X1 NOR2X1_2125 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_0_), .B(_13352_), .Y(_13353_) );
INVX1 INVX1_866 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_0_), .Y(_13354_) );
INVX1 INVX1_867 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf2), .Y(_13355_) );
NOR2X1 NOR2X1_2126 ( .gnd(gnd), .vdd(vdd), .A(_0__bF_buf8), .B(_13355_), .Y(_13356_) );
OAI21X1 OAI21X1_3787 ( .gnd(gnd), .vdd(vdd), .A(comparador_next_bF_buf2), .B(_13354_), .C(_13356__bF_buf4), .Y(_13357_) );
OR2X2 OR2X2_82 ( .gnd(gnd), .vdd(vdd), .A(_13357_), .B(_13353_), .Y(_13241__0_) );
OAI21X1 OAI21X1_3788 ( .gnd(gnd), .vdd(vdd), .A(_13353_), .B(concatenador_2_nonce_1_), .C(_13356__bF_buf3), .Y(_13358_) );
AOI21X1 AOI21X1_2271 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_1_), .B(_13353_), .C(_13358_), .Y(_13241__1_) );
OAI21X1 OAI21X1_3789 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_0_), .B(concatenador_2_nonce_1_), .C(comparador_next_bF_buf1), .Y(_13359_) );
INVX1 INVX1_868 ( .gnd(gnd), .vdd(vdd), .A(_13359_), .Y(_13360_) );
AND2X2 AND2X2_776 ( .gnd(gnd), .vdd(vdd), .A(_13360_), .B(concatenador_2_nonce_2_), .Y(_13361_) );
OAI21X1 OAI21X1_3790 ( .gnd(gnd), .vdd(vdd), .A(_13360_), .B(concatenador_2_nonce_2_), .C(_13356__bF_buf2), .Y(_13362_) );
NOR2X1 NOR2X1_2127 ( .gnd(gnd), .vdd(vdd), .A(_13362_), .B(_13361_), .Y(_13241__2_) );
NOR2X1 NOR2X1_2128 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_3_), .B(_13361_), .Y(_13363_) );
NAND2X1 NAND2X1_1810 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_2_), .B(concatenador_2_nonce_3_), .Y(_13364_) );
OAI21X1 OAI21X1_3791 ( .gnd(gnd), .vdd(vdd), .A(_13359_), .B(_13364_), .C(_13356__bF_buf1), .Y(_13365_) );
NOR2X1 NOR2X1_2129 ( .gnd(gnd), .vdd(vdd), .A(_13365_), .B(_13363_), .Y(_13241__3_) );
NOR2X1 NOR2X1_2130 ( .gnd(gnd), .vdd(vdd), .A(_13364_), .B(_13359_), .Y(_13366_) );
AND2X2 AND2X2_777 ( .gnd(gnd), .vdd(vdd), .A(_13366_), .B(concatenador_2_nonce_4_), .Y(_13367_) );
OAI21X1 OAI21X1_3792 ( .gnd(gnd), .vdd(vdd), .A(_13366_), .B(concatenador_2_nonce_4_), .C(_13356__bF_buf0), .Y(_13368_) );
NOR2X1 NOR2X1_2131 ( .gnd(gnd), .vdd(vdd), .A(_13368_), .B(_13367_), .Y(_13241__4_) );
AND2X2 AND2X2_778 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_2_), .B(concatenador_2_nonce_3_), .Y(_13369_) );
NAND3X1 NAND3X1_678 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_4_), .B(concatenador_2_nonce_5_), .C(_13369_), .Y(_13370_) );
NOR2X1 NOR2X1_2132 ( .gnd(gnd), .vdd(vdd), .A(_13359_), .B(_13370_), .Y(_13371_) );
OAI21X1 OAI21X1_3793 ( .gnd(gnd), .vdd(vdd), .A(_13367_), .B(concatenador_2_nonce_5_), .C(_13356__bF_buf4), .Y(_13372_) );
NOR2X1 NOR2X1_2133 ( .gnd(gnd), .vdd(vdd), .A(_13371_), .B(_13372_), .Y(_13241__5_) );
AND2X2 AND2X2_779 ( .gnd(gnd), .vdd(vdd), .A(_13371_), .B(concatenador_2_nonce_6_), .Y(_13373_) );
OAI21X1 OAI21X1_3794 ( .gnd(gnd), .vdd(vdd), .A(_13371_), .B(concatenador_2_nonce_6_), .C(_13356__bF_buf3), .Y(_13374_) );
NOR2X1 NOR2X1_2134 ( .gnd(gnd), .vdd(vdd), .A(_13374_), .B(_13373_), .Y(_13241__6_) );
NOR2X1 NOR2X1_2135 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_7_), .B(_13373_), .Y(_13375_) );
AND2X2 AND2X2_780 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_6_), .B(concatenador_2_nonce_7_), .Y(_13376_) );
NAND2X1 NAND2X1_1811 ( .gnd(gnd), .vdd(vdd), .A(_13376_), .B(_13371_), .Y(_13242_) );
NAND2X1 NAND2X1_1812 ( .gnd(gnd), .vdd(vdd), .A(_13356__bF_buf2), .B(_13242_), .Y(_13243_) );
NOR2X1 NOR2X1_2136 ( .gnd(gnd), .vdd(vdd), .A(_13243_), .B(_13375_), .Y(_13241__7_) );
INVX1 INVX1_869 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_8_), .Y(_13244_) );
OR2X2 OR2X2_83 ( .gnd(gnd), .vdd(vdd), .A(_13242_), .B(_13244_), .Y(_13245_) );
INVX4 INVX4_156 ( .gnd(gnd), .vdd(vdd), .A(_13356__bF_buf1), .Y(_13246_) );
AOI21X1 AOI21X1_2272 ( .gnd(gnd), .vdd(vdd), .A(_13244_), .B(_13242_), .C(_13246_), .Y(_13247_) );
AND2X2 AND2X2_781 ( .gnd(gnd), .vdd(vdd), .A(_13245_), .B(_13247_), .Y(_13241__8_) );
INVX1 INVX1_870 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_9_), .Y(_13248_) );
NAND2X1 NAND2X1_1813 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_8_), .B(concatenador_2_nonce_9_), .Y(_13249_) );
OAI21X1 OAI21X1_3795 ( .gnd(gnd), .vdd(vdd), .A(_13242_), .B(_13249_), .C(_13356__bF_buf0), .Y(_13250_) );
AOI21X1 AOI21X1_2273 ( .gnd(gnd), .vdd(vdd), .A(_13248_), .B(_13245_), .C(_13250_), .Y(_13241__9_) );
OAI21X1 OAI21X1_3796 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_0_), .B(concatenador_2_nonce_1_), .C(_13369_), .Y(_13251_) );
NAND3X1 NAND3X1_679 ( .gnd(gnd), .vdd(vdd), .A(comparador_next_bF_buf0), .B(concatenador_2_nonce_4_), .C(concatenador_2_nonce_5_), .Y(_13252_) );
AND2X2 AND2X2_782 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_8_), .B(concatenador_2_nonce_9_), .Y(_13253_) );
NAND2X1 NAND2X1_1814 ( .gnd(gnd), .vdd(vdd), .A(_13376_), .B(_13253_), .Y(_13254_) );
NOR3X1 NOR3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_13254_), .B(_13252_), .C(_13251_), .Y(_13255_) );
OAI21X1 OAI21X1_3797 ( .gnd(gnd), .vdd(vdd), .A(_13255_), .B(concatenador_2_nonce_10_), .C(_13356__bF_buf4), .Y(_13256_) );
AOI21X1 AOI21X1_2274 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_10_), .B(_13255_), .C(_13256_), .Y(_13241__10_) );
AOI21X1 AOI21X1_2275 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_10_), .B(_13255_), .C(concatenador_2_nonce_11_), .Y(_13257_) );
INVX1 INVX1_871 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_1_), .Y(_13258_) );
AOI21X1 AOI21X1_2276 ( .gnd(gnd), .vdd(vdd), .A(_13354_), .B(_13258_), .C(_13364_), .Y(_13259_) );
INVX1 INVX1_872 ( .gnd(gnd), .vdd(vdd), .A(_13252_), .Y(_13260_) );
NAND2X1 NAND2X1_1815 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_6_), .B(concatenador_2_nonce_7_), .Y(_13261_) );
NOR2X1 NOR2X1_2137 ( .gnd(gnd), .vdd(vdd), .A(_13261_), .B(_13249_), .Y(_13262_) );
NAND3X1 NAND3X1_680 ( .gnd(gnd), .vdd(vdd), .A(_13260_), .B(_13259_), .C(_13262_), .Y(_13263_) );
NAND2X1 NAND2X1_1816 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_10_), .B(concatenador_2_nonce_11_), .Y(_13264_) );
OAI21X1 OAI21X1_3798 ( .gnd(gnd), .vdd(vdd), .A(_13263_), .B(_13264_), .C(_13356__bF_buf3), .Y(_13265_) );
NOR2X1 NOR2X1_2138 ( .gnd(gnd), .vdd(vdd), .A(_13265_), .B(_13257_), .Y(_13241__11_) );
NOR2X1 NOR2X1_2139 ( .gnd(gnd), .vdd(vdd), .A(_13264_), .B(_13263_), .Y(_13266_) );
OAI21X1 OAI21X1_3799 ( .gnd(gnd), .vdd(vdd), .A(_13266_), .B(concatenador_2_nonce_12_), .C(_13356__bF_buf2), .Y(_13267_) );
AND2X2 AND2X2_783 ( .gnd(gnd), .vdd(vdd), .A(_13266_), .B(concatenador_2_nonce_12_), .Y(_13268_) );
NOR2X1 NOR2X1_2140 ( .gnd(gnd), .vdd(vdd), .A(_13267_), .B(_13268_), .Y(_13241__12_) );
OAI21X1 OAI21X1_3800 ( .gnd(gnd), .vdd(vdd), .A(_13268_), .B(concatenador_2_nonce_13_), .C(_13356__bF_buf1), .Y(_13269_) );
AOI21X1 AOI21X1_2277 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_13_), .B(_13268_), .C(_13269_), .Y(_13241__13_) );
OR2X2 OR2X2_84 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_0_), .B(concatenador_2_nonce_1_), .Y(_13270_) );
NAND3X1 NAND3X1_681 ( .gnd(gnd), .vdd(vdd), .A(_13376_), .B(_13253_), .C(_13270_), .Y(_13271_) );
NOR3X1 NOR3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_13370_), .B(_13352_), .C(_13271_), .Y(_13272_) );
NAND2X1 NAND2X1_1817 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_12_), .B(concatenador_2_nonce_13_), .Y(_13273_) );
NOR2X1 NOR2X1_2141 ( .gnd(gnd), .vdd(vdd), .A(_13264_), .B(_13273_), .Y(_13274_) );
AND2X2 AND2X2_784 ( .gnd(gnd), .vdd(vdd), .A(_13272_), .B(_13274_), .Y(_13275_) );
OAI21X1 OAI21X1_3801 ( .gnd(gnd), .vdd(vdd), .A(_13275_), .B(concatenador_2_nonce_14_), .C(_13356__bF_buf0), .Y(_13276_) );
AOI21X1 AOI21X1_2278 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_14_), .B(_13275_), .C(_13276_), .Y(_13241__14_) );
INVX1 INVX1_873 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_15_), .Y(_13277_) );
NAND3X1 NAND3X1_682 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_14_), .B(_13274_), .C(_13272_), .Y(_13278_) );
NOR2X1 NOR2X1_2142 ( .gnd(gnd), .vdd(vdd), .A(_13277_), .B(_13278_), .Y(_13279_) );
AND2X2 AND2X2_785 ( .gnd(gnd), .vdd(vdd), .A(_13278_), .B(_13277_), .Y(_13280_) );
NOR3X1 NOR3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_13279_), .B(_13246_), .C(_13280_), .Y(_13241__15_) );
AND2X2 AND2X2_786 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_14_), .B(concatenador_2_nonce_15_), .Y(_13281_) );
NAND2X1 NAND2X1_1818 ( .gnd(gnd), .vdd(vdd), .A(_13281_), .B(_13274_), .Y(_13282_) );
INVX1 INVX1_874 ( .gnd(gnd), .vdd(vdd), .A(_13282_), .Y(_13283_) );
AND2X2 AND2X2_787 ( .gnd(gnd), .vdd(vdd), .A(_13272_), .B(_13283_), .Y(_13284_) );
OAI21X1 OAI21X1_3802 ( .gnd(gnd), .vdd(vdd), .A(_13284_), .B(concatenador_2_nonce_16_), .C(_13356__bF_buf4), .Y(_13285_) );
AOI21X1 AOI21X1_2279 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_16_), .B(_13284_), .C(_13285_), .Y(_13241__16_) );
INVX2 INVX2_394 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_17_), .Y(_13286_) );
NAND3X1 NAND3X1_683 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_16_), .B(_13283_), .C(_13272_), .Y(_13287_) );
XNOR2X1 XNOR2X1_562 ( .gnd(gnd), .vdd(vdd), .A(_13287_), .B(_13286_), .Y(_13288_) );
NOR2X1 NOR2X1_2143 ( .gnd(gnd), .vdd(vdd), .A(_13246_), .B(_13288_), .Y(_13241__17_) );
NOR2X1 NOR2X1_2144 ( .gnd(gnd), .vdd(vdd), .A(_13286_), .B(_13287_), .Y(_13289_) );
OAI21X1 OAI21X1_3803 ( .gnd(gnd), .vdd(vdd), .A(_13289_), .B(concatenador_2_nonce_18_), .C(_13356__bF_buf3), .Y(_13290_) );
AOI21X1 AOI21X1_2280 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_18_), .B(_13289_), .C(_13290_), .Y(_13241__18_) );
NAND2X1 NAND2X1_1819 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_16_), .B(concatenador_2_nonce_17_), .Y(_13291_) );
NOR2X1 NOR2X1_2145 ( .gnd(gnd), .vdd(vdd), .A(_13291_), .B(_13282_), .Y(_13292_) );
NAND3X1 NAND3X1_684 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_18_), .B(_13272_), .C(_13292_), .Y(_13293_) );
NAND2X1 NAND2X1_1820 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_19_), .B(_13293_), .Y(_13294_) );
OR2X2 OR2X2_85 ( .gnd(gnd), .vdd(vdd), .A(_13293_), .B(concatenador_2_nonce_19_), .Y(_13295_) );
AOI21X1 AOI21X1_2281 ( .gnd(gnd), .vdd(vdd), .A(_13294_), .B(_13295_), .C(_13246_), .Y(_13241__19_) );
INVX1 INVX1_875 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_20_), .Y(_13296_) );
NAND3X1 NAND3X1_685 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_13_), .B(concatenador_2_nonce_14_), .C(concatenador_2_nonce_15_), .Y(_13297_) );
NOR2X1 NOR2X1_2146 ( .gnd(gnd), .vdd(vdd), .A(_13291_), .B(_13297_), .Y(_13298_) );
NAND3X1 NAND3X1_686 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_12_), .B(concatenador_2_nonce_18_), .C(concatenador_2_nonce_19_), .Y(_13299_) );
NOR2X1 NOR2X1_2147 ( .gnd(gnd), .vdd(vdd), .A(_13264_), .B(_13299_), .Y(_13300_) );
NAND2X1 NAND2X1_1821 ( .gnd(gnd), .vdd(vdd), .A(_13298_), .B(_13300_), .Y(_13301_) );
OAI21X1 OAI21X1_3804 ( .gnd(gnd), .vdd(vdd), .A(_13301_), .B(_13263_), .C(_13296_), .Y(_13302_) );
NAND2X1 NAND2X1_1822 ( .gnd(gnd), .vdd(vdd), .A(_13356__bF_buf2), .B(_13302_), .Y(_13303_) );
AND2X2 AND2X2_788 ( .gnd(gnd), .vdd(vdd), .A(_13298_), .B(_13300_), .Y(_13304_) );
NAND2X1 NAND2X1_1823 ( .gnd(gnd), .vdd(vdd), .A(_13304_), .B(_13255_), .Y(_13305_) );
NOR2X1 NOR2X1_2148 ( .gnd(gnd), .vdd(vdd), .A(_13296_), .B(_13305_), .Y(_13306_) );
NOR2X1 NOR2X1_2149 ( .gnd(gnd), .vdd(vdd), .A(_13303_), .B(_13306_), .Y(_13241__20_) );
NOR2X1 NOR2X1_2150 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_21_), .B(_13306_), .Y(_13307_) );
NAND2X1 NAND2X1_1824 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_20_), .B(concatenador_2_nonce_21_), .Y(_13308_) );
OAI21X1 OAI21X1_3805 ( .gnd(gnd), .vdd(vdd), .A(_13305_), .B(_13308_), .C(_13356__bF_buf1), .Y(_13309_) );
NOR2X1 NOR2X1_2151 ( .gnd(gnd), .vdd(vdd), .A(_13309_), .B(_13307_), .Y(_13241__21_) );
NOR3X1 NOR3X1_21 ( .gnd(gnd), .vdd(vdd), .A(_13263_), .B(_13308_), .C(_13301_), .Y(_13310_) );
OAI21X1 OAI21X1_3806 ( .gnd(gnd), .vdd(vdd), .A(_13310_), .B(concatenador_2_nonce_22_), .C(_13356__bF_buf0), .Y(_13311_) );
INVX2 INVX2_395 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_22_), .Y(_13312_) );
INVX1 INVX1_876 ( .gnd(gnd), .vdd(vdd), .A(_13308_), .Y(_13313_) );
NAND3X1 NAND3X1_687 ( .gnd(gnd), .vdd(vdd), .A(_13304_), .B(_13313_), .C(_13255_), .Y(_13314_) );
NOR2X1 NOR2X1_2152 ( .gnd(gnd), .vdd(vdd), .A(_13312_), .B(_13314_), .Y(_13315_) );
NOR2X1 NOR2X1_2153 ( .gnd(gnd), .vdd(vdd), .A(_13315_), .B(_13311_), .Y(_13241__22_) );
INVX1 INVX1_877 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_23_), .Y(_13316_) );
NOR3X1 NOR3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_13312_), .B(_13316_), .C(_13314_), .Y(_13317_) );
OAI21X1 OAI21X1_3807 ( .gnd(gnd), .vdd(vdd), .A(_13315_), .B(concatenador_2_nonce_23_), .C(_13356__bF_buf4), .Y(_13318_) );
NOR2X1 NOR2X1_2154 ( .gnd(gnd), .vdd(vdd), .A(_13317_), .B(_13318_), .Y(_13241__23_) );
OAI21X1 OAI21X1_3808 ( .gnd(gnd), .vdd(vdd), .A(_13317_), .B(concatenador_2_nonce_24_), .C(_13356__bF_buf3), .Y(_13319_) );
AOI21X1 AOI21X1_2282 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_24_), .B(_13317_), .C(_13319_), .Y(_13241__24_) );
INVX1 INVX1_878 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_24_), .Y(_13320_) );
NAND3X1 NAND3X1_688 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_22_), .B(concatenador_2_nonce_23_), .C(_13310_), .Y(_13321_) );
OAI21X1 OAI21X1_3809 ( .gnd(gnd), .vdd(vdd), .A(_13321_), .B(_13320_), .C(concatenador_2_nonce_25_), .Y(_13322_) );
INVX1 INVX1_879 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_25_), .Y(_13323_) );
NAND3X1 NAND3X1_689 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_24_), .B(_13323_), .C(_13317_), .Y(_13324_) );
AOI21X1 AOI21X1_2283 ( .gnd(gnd), .vdd(vdd), .A(_13322_), .B(_13324_), .C(_13246_), .Y(_13241__25_) );
NAND3X1 NAND3X1_690 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_23_), .B(concatenador_2_nonce_24_), .C(concatenador_2_nonce_25_), .Y(_13325_) );
NOR3X1 NOR3X1_23 ( .gnd(gnd), .vdd(vdd), .A(_13312_), .B(_13325_), .C(_13314_), .Y(_13326_) );
OAI21X1 OAI21X1_3810 ( .gnd(gnd), .vdd(vdd), .A(_13326_), .B(concatenador_2_nonce_26_), .C(_13356__bF_buf2), .Y(_13327_) );
AOI21X1 AOI21X1_2284 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_26_), .B(_13326_), .C(_13327_), .Y(_13241__26_) );
INVX1 INVX1_880 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_26_), .Y(_13328_) );
INVX1 INVX1_881 ( .gnd(gnd), .vdd(vdd), .A(_13325_), .Y(_13329_) );
NAND3X1 NAND3X1_691 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_22_), .B(_13329_), .C(_13310_), .Y(_13330_) );
OAI21X1 OAI21X1_3811 ( .gnd(gnd), .vdd(vdd), .A(_13330_), .B(_13328_), .C(concatenador_2_nonce_27_), .Y(_13331_) );
INVX1 INVX1_882 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_27_), .Y(_13332_) );
NAND3X1 NAND3X1_692 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_26_), .B(_13332_), .C(_13326_), .Y(_13333_) );
AOI21X1 AOI21X1_2285 ( .gnd(gnd), .vdd(vdd), .A(_13331_), .B(_13333_), .C(_13246_), .Y(_13241__27_) );
NAND3X1 NAND3X1_693 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_22_), .B(concatenador_2_nonce_26_), .C(concatenador_2_nonce_27_), .Y(_13334_) );
NOR2X1 NOR2X1_2155 ( .gnd(gnd), .vdd(vdd), .A(_13308_), .B(_13334_), .Y(_13335_) );
NAND2X1 NAND2X1_1825 ( .gnd(gnd), .vdd(vdd), .A(_13329_), .B(_13335_), .Y(_13336_) );
NOR3X1 NOR3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_13263_), .B(_13336_), .C(_13301_), .Y(_13337_) );
OAI21X1 OAI21X1_3812 ( .gnd(gnd), .vdd(vdd), .A(_13337_), .B(concatenador_2_nonce_28_), .C(_13356__bF_buf1), .Y(_13338_) );
INVX1 INVX1_883 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_28_), .Y(_13339_) );
AND2X2 AND2X2_789 ( .gnd(gnd), .vdd(vdd), .A(_13335_), .B(_13329_), .Y(_13340_) );
NAND3X1 NAND3X1_694 ( .gnd(gnd), .vdd(vdd), .A(_13304_), .B(_13340_), .C(_13255_), .Y(_13341_) );
NOR2X1 NOR2X1_2156 ( .gnd(gnd), .vdd(vdd), .A(_13339_), .B(_13341_), .Y(_13342_) );
NOR2X1 NOR2X1_2157 ( .gnd(gnd), .vdd(vdd), .A(_13342_), .B(_13338_), .Y(_13241__28_) );
INVX1 INVX1_884 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_29_), .Y(_13343_) );
NOR3X1 NOR3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_13339_), .B(_13343_), .C(_13341_), .Y(_13344_) );
OAI21X1 OAI21X1_3813 ( .gnd(gnd), .vdd(vdd), .A(_13342_), .B(concatenador_2_nonce_29_), .C(_13356__bF_buf0), .Y(_13345_) );
NOR2X1 NOR2X1_2158 ( .gnd(gnd), .vdd(vdd), .A(_13344_), .B(_13345_), .Y(_13241__29_) );
OAI21X1 OAI21X1_3814 ( .gnd(gnd), .vdd(vdd), .A(_13344_), .B(concatenador_2_nonce_30_), .C(_13356__bF_buf4), .Y(_13346_) );
AOI21X1 AOI21X1_2286 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_30_), .B(_13344_), .C(_13346_), .Y(_13241__30_) );
INVX1 INVX1_885 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_30_), .Y(_13347_) );
NAND3X1 NAND3X1_695 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_28_), .B(concatenador_2_nonce_29_), .C(_13337_), .Y(_13348_) );
OAI21X1 OAI21X1_3815 ( .gnd(gnd), .vdd(vdd), .A(_13348_), .B(_13347_), .C(concatenador_2_nonce_31_), .Y(_13349_) );
INVX1 INVX1_886 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_31_), .Y(_13350_) );
NAND3X1 NAND3X1_696 ( .gnd(gnd), .vdd(vdd), .A(concatenador_2_nonce_30_), .B(_13350_), .C(_13344_), .Y(_13351_) );
AOI21X1 AOI21X1_2287 ( .gnd(gnd), .vdd(vdd), .A(_13349_), .B(_13351_), .C(_13246_), .Y(_13241__31_) );
DFFPOSX1 DFFPOSX1_1794 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(_13241__0_), .Q(concatenador_2_nonce_0_) );
DFFPOSX1 DFFPOSX1_1795 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(_13241__1_), .Q(concatenador_2_nonce_1_) );
DFFPOSX1 DFFPOSX1_1796 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(_13241__2_), .Q(concatenador_2_nonce_2_) );
DFFPOSX1 DFFPOSX1_1797 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(_13241__3_), .Q(concatenador_2_nonce_3_) );
DFFPOSX1 DFFPOSX1_1798 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_13241__4_), .Q(concatenador_2_nonce_4_) );
DFFPOSX1 DFFPOSX1_1799 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_13241__5_), .Q(concatenador_2_nonce_5_) );
DFFPOSX1 DFFPOSX1_1800 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_13241__6_), .Q(concatenador_2_nonce_6_) );
DFFPOSX1 DFFPOSX1_1801 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_13241__7_), .Q(concatenador_2_nonce_7_) );
DFFPOSX1 DFFPOSX1_1802 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_13241__8_), .Q(concatenador_2_nonce_8_) );
DFFPOSX1 DFFPOSX1_1803 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_13241__9_), .Q(concatenador_2_nonce_9_) );
DFFPOSX1 DFFPOSX1_1804 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_13241__10_), .Q(concatenador_2_nonce_10_) );
DFFPOSX1 DFFPOSX1_1805 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_13241__11_), .Q(concatenador_2_nonce_11_) );
DFFPOSX1 DFFPOSX1_1806 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_13241__12_), .Q(concatenador_2_nonce_12_) );
DFFPOSX1 DFFPOSX1_1807 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_13241__13_), .Q(concatenador_2_nonce_13_) );
DFFPOSX1 DFFPOSX1_1808 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_13241__14_), .Q(concatenador_2_nonce_14_) );
DFFPOSX1 DFFPOSX1_1809 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_13241__15_), .Q(concatenador_2_nonce_15_) );
DFFPOSX1 DFFPOSX1_1810 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_13241__16_), .Q(concatenador_2_nonce_16_) );
DFFPOSX1 DFFPOSX1_1811 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_13241__17_), .Q(concatenador_2_nonce_17_) );
DFFPOSX1 DFFPOSX1_1812 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_13241__18_), .Q(concatenador_2_nonce_18_) );
DFFPOSX1 DFFPOSX1_1813 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_13241__19_), .Q(concatenador_2_nonce_19_) );
DFFPOSX1 DFFPOSX1_1814 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_13241__20_), .Q(concatenador_2_nonce_20_) );
DFFPOSX1 DFFPOSX1_1815 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_13241__21_), .Q(concatenador_2_nonce_21_) );
DFFPOSX1 DFFPOSX1_1816 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_13241__22_), .Q(concatenador_2_nonce_22_) );
DFFPOSX1 DFFPOSX1_1817 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_13241__23_), .Q(concatenador_2_nonce_23_) );
DFFPOSX1 DFFPOSX1_1818 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_13241__24_), .Q(concatenador_2_nonce_24_) );
DFFPOSX1 DFFPOSX1_1819 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_13241__25_), .Q(concatenador_2_nonce_25_) );
DFFPOSX1 DFFPOSX1_1820 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_13241__26_), .Q(concatenador_2_nonce_26_) );
DFFPOSX1 DFFPOSX1_1821 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_13241__27_), .Q(concatenador_2_nonce_27_) );
DFFPOSX1 DFFPOSX1_1822 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_13241__28_), .Q(concatenador_2_nonce_28_) );
DFFPOSX1 DFFPOSX1_1823 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_13241__29_), .Q(concatenador_2_nonce_29_) );
DFFPOSX1 DFFPOSX1_1824 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_13241__30_), .Q(concatenador_2_nonce_30_) );
DFFPOSX1 DFFPOSX1_1825 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_13241__31_), .Q(concatenador_2_nonce_31_) );
INVX1 INVX1_887 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf1), .Y(_13483_) );
NOR2X1 NOR2X1_2159 ( .gnd(gnd), .vdd(vdd), .A(_0__bF_buf7), .B(_13483_), .Y(_13484_) );
INVX4 INVX4_157 ( .gnd(gnd), .vdd(vdd), .A(_13484__bF_buf3), .Y(_13485_) );
INVX2 INVX2_396 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_0_), .Y(_13486_) );
NAND2X1 NAND2X1_1826 ( .gnd(gnd), .vdd(vdd), .A(comparador_next_bF_buf3), .B(_13486_), .Y(_13487_) );
OR2X2 OR2X2_86 ( .gnd(gnd), .vdd(vdd), .A(_13486_), .B(comparador_next_bF_buf2), .Y(_13488_) );
AOI21X1 AOI21X1_2288 ( .gnd(gnd), .vdd(vdd), .A(_13487_), .B(_13488_), .C(_13485_), .Y(_13377__0_) );
AOI21X1 AOI21X1_2289 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_1_), .B(_13487_), .C(_13485_), .Y(_13489_) );
OAI21X1 OAI21X1_3816 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_1_), .B(_13487_), .C(_13489_), .Y(_13377__1_) );
OAI21X1 OAI21X1_3817 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_0_), .B(concatenador_3_nonce_1_), .C(comparador_next_bF_buf1), .Y(_13490_) );
INVX1 INVX1_888 ( .gnd(gnd), .vdd(vdd), .A(_13490_), .Y(_13491_) );
AND2X2 AND2X2_790 ( .gnd(gnd), .vdd(vdd), .A(_13491_), .B(concatenador_3_nonce_2_), .Y(_13492_) );
OAI21X1 OAI21X1_3818 ( .gnd(gnd), .vdd(vdd), .A(_13491_), .B(concatenador_3_nonce_2_), .C(_13484__bF_buf2), .Y(_13493_) );
NOR2X1 NOR2X1_2160 ( .gnd(gnd), .vdd(vdd), .A(_13493_), .B(_13492_), .Y(_13377__2_) );
NOR2X1 NOR2X1_2161 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_3_), .B(_13492_), .Y(_13494_) );
NAND2X1 NAND2X1_1827 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_2_), .B(concatenador_3_nonce_3_), .Y(_13495_) );
OAI21X1 OAI21X1_3819 ( .gnd(gnd), .vdd(vdd), .A(_13490_), .B(_13495_), .C(_13484__bF_buf1), .Y(_13496_) );
NOR2X1 NOR2X1_2162 ( .gnd(gnd), .vdd(vdd), .A(_13496_), .B(_13494_), .Y(_13377__3_) );
NOR2X1 NOR2X1_2163 ( .gnd(gnd), .vdd(vdd), .A(_13495_), .B(_13490_), .Y(_13497_) );
AND2X2 AND2X2_791 ( .gnd(gnd), .vdd(vdd), .A(_13497_), .B(concatenador_3_nonce_4_), .Y(_13498_) );
OAI21X1 OAI21X1_3820 ( .gnd(gnd), .vdd(vdd), .A(_13497_), .B(concatenador_3_nonce_4_), .C(_13484__bF_buf0), .Y(_13499_) );
NOR2X1 NOR2X1_2164 ( .gnd(gnd), .vdd(vdd), .A(_13499_), .B(_13498_), .Y(_13377__4_) );
AND2X2 AND2X2_792 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_2_), .B(concatenador_3_nonce_3_), .Y(_13500_) );
NAND3X1 NAND3X1_697 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_4_), .B(concatenador_3_nonce_5_), .C(_13500_), .Y(_13501_) );
NOR2X1 NOR2X1_2165 ( .gnd(gnd), .vdd(vdd), .A(_13490_), .B(_13501_), .Y(_13502_) );
OAI21X1 OAI21X1_3821 ( .gnd(gnd), .vdd(vdd), .A(_13498_), .B(concatenador_3_nonce_5_), .C(_13484__bF_buf3), .Y(_13503_) );
NOR2X1 NOR2X1_2166 ( .gnd(gnd), .vdd(vdd), .A(_13502_), .B(_13503_), .Y(_13377__5_) );
AND2X2 AND2X2_793 ( .gnd(gnd), .vdd(vdd), .A(_13502_), .B(concatenador_3_nonce_6_), .Y(_13504_) );
OAI21X1 OAI21X1_3822 ( .gnd(gnd), .vdd(vdd), .A(_13502_), .B(concatenador_3_nonce_6_), .C(_13484__bF_buf2), .Y(_13505_) );
NOR2X1 NOR2X1_2167 ( .gnd(gnd), .vdd(vdd), .A(_13505_), .B(_13504_), .Y(_13377__6_) );
NOR2X1 NOR2X1_2168 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_7_), .B(_13504_), .Y(_13506_) );
AND2X2 AND2X2_794 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_6_), .B(concatenador_3_nonce_7_), .Y(_13507_) );
NAND2X1 NAND2X1_1828 ( .gnd(gnd), .vdd(vdd), .A(_13507_), .B(_13502_), .Y(_13378_) );
NAND2X1 NAND2X1_1829 ( .gnd(gnd), .vdd(vdd), .A(_13484__bF_buf1), .B(_13378_), .Y(_13379_) );
NOR2X1 NOR2X1_2169 ( .gnd(gnd), .vdd(vdd), .A(_13379_), .B(_13506_), .Y(_13377__7_) );
INVX1 INVX1_889 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_8_), .Y(_13380_) );
OR2X2 OR2X2_87 ( .gnd(gnd), .vdd(vdd), .A(_13378_), .B(_13380_), .Y(_13381_) );
AOI21X1 AOI21X1_2290 ( .gnd(gnd), .vdd(vdd), .A(_13380_), .B(_13378_), .C(_13485_), .Y(_13382_) );
AND2X2 AND2X2_795 ( .gnd(gnd), .vdd(vdd), .A(_13381_), .B(_13382_), .Y(_13377__8_) );
INVX1 INVX1_890 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_9_), .Y(_13383_) );
NAND2X1 NAND2X1_1830 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_8_), .B(concatenador_3_nonce_9_), .Y(_13384_) );
OAI21X1 OAI21X1_3823 ( .gnd(gnd), .vdd(vdd), .A(_13378_), .B(_13384_), .C(_13484__bF_buf0), .Y(_13385_) );
AOI21X1 AOI21X1_2291 ( .gnd(gnd), .vdd(vdd), .A(_13383_), .B(_13381_), .C(_13385_), .Y(_13377__9_) );
OAI21X1 OAI21X1_3824 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_0_), .B(concatenador_3_nonce_1_), .C(_13500_), .Y(_13386_) );
NAND3X1 NAND3X1_698 ( .gnd(gnd), .vdd(vdd), .A(comparador_next_bF_buf0), .B(concatenador_3_nonce_4_), .C(concatenador_3_nonce_5_), .Y(_13387_) );
AND2X2 AND2X2_796 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_8_), .B(concatenador_3_nonce_9_), .Y(_13388_) );
NAND2X1 NAND2X1_1831 ( .gnd(gnd), .vdd(vdd), .A(_13507_), .B(_13388_), .Y(_13389_) );
NOR3X1 NOR3X1_26 ( .gnd(gnd), .vdd(vdd), .A(_13389_), .B(_13387_), .C(_13386_), .Y(_13390_) );
OAI21X1 OAI21X1_3825 ( .gnd(gnd), .vdd(vdd), .A(_13390_), .B(concatenador_3_nonce_10_), .C(_13484__bF_buf3), .Y(_13391_) );
AOI21X1 AOI21X1_2292 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_10_), .B(_13390_), .C(_13391_), .Y(_13377__10_) );
AOI21X1 AOI21X1_2293 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_10_), .B(_13390_), .C(concatenador_3_nonce_11_), .Y(_13392_) );
INVX1 INVX1_891 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_1_), .Y(_13393_) );
AOI21X1 AOI21X1_2294 ( .gnd(gnd), .vdd(vdd), .A(_13486_), .B(_13393_), .C(_13495_), .Y(_13394_) );
INVX1 INVX1_892 ( .gnd(gnd), .vdd(vdd), .A(_13387_), .Y(_13395_) );
NAND2X1 NAND2X1_1832 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_6_), .B(concatenador_3_nonce_7_), .Y(_13396_) );
NOR2X1 NOR2X1_2170 ( .gnd(gnd), .vdd(vdd), .A(_13396_), .B(_13384_), .Y(_13397_) );
NAND3X1 NAND3X1_699 ( .gnd(gnd), .vdd(vdd), .A(_13395_), .B(_13394_), .C(_13397_), .Y(_13398_) );
NAND2X1 NAND2X1_1833 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_10_), .B(concatenador_3_nonce_11_), .Y(_13399_) );
OAI21X1 OAI21X1_3826 ( .gnd(gnd), .vdd(vdd), .A(_13398_), .B(_13399_), .C(_13484__bF_buf2), .Y(_13400_) );
NOR2X1 NOR2X1_2171 ( .gnd(gnd), .vdd(vdd), .A(_13400_), .B(_13392_), .Y(_13377__11_) );
NOR2X1 NOR2X1_2172 ( .gnd(gnd), .vdd(vdd), .A(_13399_), .B(_13398_), .Y(_13401_) );
OAI21X1 OAI21X1_3827 ( .gnd(gnd), .vdd(vdd), .A(_13401_), .B(concatenador_3_nonce_12_), .C(_13484__bF_buf1), .Y(_13402_) );
AND2X2 AND2X2_797 ( .gnd(gnd), .vdd(vdd), .A(_13401_), .B(concatenador_3_nonce_12_), .Y(_13403_) );
NOR2X1 NOR2X1_2173 ( .gnd(gnd), .vdd(vdd), .A(_13402_), .B(_13403_), .Y(_13377__12_) );
OAI21X1 OAI21X1_3828 ( .gnd(gnd), .vdd(vdd), .A(_13403_), .B(concatenador_3_nonce_13_), .C(_13484__bF_buf0), .Y(_13404_) );
AOI21X1 AOI21X1_2295 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_13_), .B(_13403_), .C(_13404_), .Y(_13377__13_) );
OR2X2 OR2X2_88 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_0_), .B(concatenador_3_nonce_1_), .Y(_13405_) );
NAND3X1 NAND3X1_700 ( .gnd(gnd), .vdd(vdd), .A(_13507_), .B(_13388_), .C(_13405_), .Y(_13406_) );
NOR2X1 NOR2X1_2174 ( .gnd(gnd), .vdd(vdd), .A(_13501_), .B(_13406_), .Y(_13407_) );
NAND2X1 NAND2X1_1834 ( .gnd(gnd), .vdd(vdd), .A(comparador_next_bF_buf3), .B(_13407_), .Y(_13408_) );
NAND2X1 NAND2X1_1835 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_12_), .B(concatenador_3_nonce_13_), .Y(_13409_) );
NOR2X1 NOR2X1_2175 ( .gnd(gnd), .vdd(vdd), .A(_13399_), .B(_13409_), .Y(_13410_) );
INVX1 INVX1_893 ( .gnd(gnd), .vdd(vdd), .A(_13410_), .Y(_13411_) );
NOR2X1 NOR2X1_2176 ( .gnd(gnd), .vdd(vdd), .A(_13411_), .B(_13408_), .Y(_13412_) );
OAI21X1 OAI21X1_3829 ( .gnd(gnd), .vdd(vdd), .A(_13412_), .B(concatenador_3_nonce_14_), .C(_13484__bF_buf3), .Y(_13413_) );
AOI21X1 AOI21X1_2296 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_14_), .B(_13412_), .C(_13413_), .Y(_13377__14_) );
NAND3X1 NAND3X1_701 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_14_), .B(concatenador_3_nonce_15_), .C(_13410_), .Y(_13414_) );
NOR2X1 NOR2X1_2177 ( .gnd(gnd), .vdd(vdd), .A(_13414_), .B(_13408_), .Y(_13415_) );
AOI21X1 AOI21X1_2297 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_14_), .B(_13412_), .C(concatenador_3_nonce_15_), .Y(_13416_) );
NOR3X1 NOR3X1_27 ( .gnd(gnd), .vdd(vdd), .A(_13485_), .B(_13415_), .C(_13416_), .Y(_13377__15_) );
OAI21X1 OAI21X1_3830 ( .gnd(gnd), .vdd(vdd), .A(_13415_), .B(concatenador_3_nonce_16_), .C(_13484__bF_buf2), .Y(_13417_) );
AOI21X1 AOI21X1_2298 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_16_), .B(_13415_), .C(_13417_), .Y(_13377__16_) );
AND2X2 AND2X2_798 ( .gnd(gnd), .vdd(vdd), .A(_13407_), .B(comparador_next_bF_buf2), .Y(_13418_) );
NAND2X1 NAND2X1_1836 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_16_), .B(concatenador_3_nonce_17_), .Y(_13419_) );
NOR2X1 NOR2X1_2178 ( .gnd(gnd), .vdd(vdd), .A(_13419_), .B(_13414_), .Y(_13420_) );
AND2X2 AND2X2_799 ( .gnd(gnd), .vdd(vdd), .A(_13418_), .B(_13420_), .Y(_13421_) );
AOI21X1 AOI21X1_2299 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_16_), .B(_13415_), .C(concatenador_3_nonce_17_), .Y(_13422_) );
NOR3X1 NOR3X1_28 ( .gnd(gnd), .vdd(vdd), .A(_13485_), .B(_13421_), .C(_13422_), .Y(_13377__17_) );
OAI21X1 OAI21X1_3831 ( .gnd(gnd), .vdd(vdd), .A(_13421_), .B(concatenador_3_nonce_18_), .C(_13484__bF_buf1), .Y(_13423_) );
AOI21X1 AOI21X1_2300 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_18_), .B(_13421_), .C(_13423_), .Y(_13377__18_) );
NAND3X1 NAND3X1_702 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_18_), .B(_13420_), .C(_13418_), .Y(_13424_) );
NAND2X1 NAND2X1_1837 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_19_), .B(_13424_), .Y(_13425_) );
OR2X2 OR2X2_89 ( .gnd(gnd), .vdd(vdd), .A(_13424_), .B(concatenador_3_nonce_19_), .Y(_13426_) );
AOI21X1 AOI21X1_2301 ( .gnd(gnd), .vdd(vdd), .A(_13425_), .B(_13426_), .C(_13485_), .Y(_13377__19_) );
INVX1 INVX1_894 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_20_), .Y(_13427_) );
NAND3X1 NAND3X1_703 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_13_), .B(concatenador_3_nonce_14_), .C(concatenador_3_nonce_15_), .Y(_13428_) );
NOR2X1 NOR2X1_2179 ( .gnd(gnd), .vdd(vdd), .A(_13419_), .B(_13428_), .Y(_13429_) );
NAND3X1 NAND3X1_704 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_12_), .B(concatenador_3_nonce_18_), .C(concatenador_3_nonce_19_), .Y(_13430_) );
NOR2X1 NOR2X1_2180 ( .gnd(gnd), .vdd(vdd), .A(_13399_), .B(_13430_), .Y(_13431_) );
NAND2X1 NAND2X1_1838 ( .gnd(gnd), .vdd(vdd), .A(_13429_), .B(_13431_), .Y(_13432_) );
OAI21X1 OAI21X1_3832 ( .gnd(gnd), .vdd(vdd), .A(_13432_), .B(_13398_), .C(_13427_), .Y(_13433_) );
NAND2X1 NAND2X1_1839 ( .gnd(gnd), .vdd(vdd), .A(_13484__bF_buf0), .B(_13433_), .Y(_13434_) );
AND2X2 AND2X2_800 ( .gnd(gnd), .vdd(vdd), .A(_13429_), .B(_13431_), .Y(_13435_) );
NAND2X1 NAND2X1_1840 ( .gnd(gnd), .vdd(vdd), .A(_13435_), .B(_13390_), .Y(_13436_) );
NOR2X1 NOR2X1_2181 ( .gnd(gnd), .vdd(vdd), .A(_13427_), .B(_13436_), .Y(_13437_) );
NOR2X1 NOR2X1_2182 ( .gnd(gnd), .vdd(vdd), .A(_13434_), .B(_13437_), .Y(_13377__20_) );
NOR2X1 NOR2X1_2183 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_21_), .B(_13437_), .Y(_13438_) );
NAND2X1 NAND2X1_1841 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_20_), .B(concatenador_3_nonce_21_), .Y(_13439_) );
OAI21X1 OAI21X1_3833 ( .gnd(gnd), .vdd(vdd), .A(_13436_), .B(_13439_), .C(_13484__bF_buf3), .Y(_13440_) );
NOR2X1 NOR2X1_2184 ( .gnd(gnd), .vdd(vdd), .A(_13440_), .B(_13438_), .Y(_13377__21_) );
NOR3X1 NOR3X1_29 ( .gnd(gnd), .vdd(vdd), .A(_13398_), .B(_13439_), .C(_13432_), .Y(_13441_) );
OAI21X1 OAI21X1_3834 ( .gnd(gnd), .vdd(vdd), .A(_13441_), .B(concatenador_3_nonce_22_), .C(_13484__bF_buf2), .Y(_13442_) );
INVX2 INVX2_397 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_22_), .Y(_13443_) );
INVX1 INVX1_895 ( .gnd(gnd), .vdd(vdd), .A(_13439_), .Y(_13444_) );
NAND3X1 NAND3X1_705 ( .gnd(gnd), .vdd(vdd), .A(_13435_), .B(_13444_), .C(_13390_), .Y(_13445_) );
NOR2X1 NOR2X1_2185 ( .gnd(gnd), .vdd(vdd), .A(_13443_), .B(_13445_), .Y(_13446_) );
NOR2X1 NOR2X1_2186 ( .gnd(gnd), .vdd(vdd), .A(_13446_), .B(_13442_), .Y(_13377__22_) );
INVX1 INVX1_896 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_23_), .Y(_13447_) );
NOR3X1 NOR3X1_30 ( .gnd(gnd), .vdd(vdd), .A(_13443_), .B(_13447_), .C(_13445_), .Y(_13448_) );
OAI21X1 OAI21X1_3835 ( .gnd(gnd), .vdd(vdd), .A(_13446_), .B(concatenador_3_nonce_23_), .C(_13484__bF_buf1), .Y(_13449_) );
NOR2X1 NOR2X1_2187 ( .gnd(gnd), .vdd(vdd), .A(_13448_), .B(_13449_), .Y(_13377__23_) );
OAI21X1 OAI21X1_3836 ( .gnd(gnd), .vdd(vdd), .A(_13448_), .B(concatenador_3_nonce_24_), .C(_13484__bF_buf0), .Y(_13450_) );
AOI21X1 AOI21X1_2302 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_24_), .B(_13448_), .C(_13450_), .Y(_13377__24_) );
INVX1 INVX1_897 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_24_), .Y(_13451_) );
NAND3X1 NAND3X1_706 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_22_), .B(concatenador_3_nonce_23_), .C(_13441_), .Y(_13452_) );
OAI21X1 OAI21X1_3837 ( .gnd(gnd), .vdd(vdd), .A(_13452_), .B(_13451_), .C(concatenador_3_nonce_25_), .Y(_13453_) );
INVX1 INVX1_898 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_25_), .Y(_13454_) );
NAND3X1 NAND3X1_707 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_24_), .B(_13454_), .C(_13448_), .Y(_13455_) );
AOI21X1 AOI21X1_2303 ( .gnd(gnd), .vdd(vdd), .A(_13453_), .B(_13455_), .C(_13485_), .Y(_13377__25_) );
NAND3X1 NAND3X1_708 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_23_), .B(concatenador_3_nonce_24_), .C(concatenador_3_nonce_25_), .Y(_13456_) );
NOR3X1 NOR3X1_31 ( .gnd(gnd), .vdd(vdd), .A(_13443_), .B(_13456_), .C(_13445_), .Y(_13457_) );
OAI21X1 OAI21X1_3838 ( .gnd(gnd), .vdd(vdd), .A(_13457_), .B(concatenador_3_nonce_26_), .C(_13484__bF_buf3), .Y(_13458_) );
AOI21X1 AOI21X1_2304 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_26_), .B(_13457_), .C(_13458_), .Y(_13377__26_) );
INVX1 INVX1_899 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_26_), .Y(_13459_) );
INVX1 INVX1_900 ( .gnd(gnd), .vdd(vdd), .A(_13456_), .Y(_13460_) );
NAND3X1 NAND3X1_709 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_22_), .B(_13460_), .C(_13441_), .Y(_13461_) );
OAI21X1 OAI21X1_3839 ( .gnd(gnd), .vdd(vdd), .A(_13461_), .B(_13459_), .C(concatenador_3_nonce_27_), .Y(_13462_) );
INVX1 INVX1_901 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_27_), .Y(_13463_) );
NAND3X1 NAND3X1_710 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_26_), .B(_13463_), .C(_13457_), .Y(_13464_) );
AOI21X1 AOI21X1_2305 ( .gnd(gnd), .vdd(vdd), .A(_13462_), .B(_13464_), .C(_13485_), .Y(_13377__27_) );
NAND3X1 NAND3X1_711 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_22_), .B(concatenador_3_nonce_26_), .C(concatenador_3_nonce_27_), .Y(_13465_) );
NOR2X1 NOR2X1_2188 ( .gnd(gnd), .vdd(vdd), .A(_13439_), .B(_13465_), .Y(_13466_) );
NAND2X1 NAND2X1_1842 ( .gnd(gnd), .vdd(vdd), .A(_13460_), .B(_13466_), .Y(_13467_) );
NOR3X1 NOR3X1_32 ( .gnd(gnd), .vdd(vdd), .A(_13398_), .B(_13467_), .C(_13432_), .Y(_13468_) );
OAI21X1 OAI21X1_3840 ( .gnd(gnd), .vdd(vdd), .A(_13468_), .B(concatenador_3_nonce_28_), .C(_13484__bF_buf2), .Y(_13469_) );
INVX1 INVX1_902 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_28_), .Y(_13470_) );
AND2X2 AND2X2_801 ( .gnd(gnd), .vdd(vdd), .A(_13466_), .B(_13460_), .Y(_13471_) );
NAND3X1 NAND3X1_712 ( .gnd(gnd), .vdd(vdd), .A(_13435_), .B(_13471_), .C(_13390_), .Y(_13472_) );
NOR2X1 NOR2X1_2189 ( .gnd(gnd), .vdd(vdd), .A(_13470_), .B(_13472_), .Y(_13473_) );
NOR2X1 NOR2X1_2190 ( .gnd(gnd), .vdd(vdd), .A(_13473_), .B(_13469_), .Y(_13377__28_) );
INVX1 INVX1_903 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_29_), .Y(_13474_) );
NOR3X1 NOR3X1_33 ( .gnd(gnd), .vdd(vdd), .A(_13470_), .B(_13474_), .C(_13472_), .Y(_13475_) );
OAI21X1 OAI21X1_3841 ( .gnd(gnd), .vdd(vdd), .A(_13473_), .B(concatenador_3_nonce_29_), .C(_13484__bF_buf1), .Y(_13476_) );
NOR2X1 NOR2X1_2191 ( .gnd(gnd), .vdd(vdd), .A(_13475_), .B(_13476_), .Y(_13377__29_) );
OAI21X1 OAI21X1_3842 ( .gnd(gnd), .vdd(vdd), .A(_13475_), .B(concatenador_3_nonce_30_), .C(_13484__bF_buf0), .Y(_13477_) );
AOI21X1 AOI21X1_2306 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_30_), .B(_13475_), .C(_13477_), .Y(_13377__30_) );
INVX1 INVX1_904 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_30_), .Y(_13478_) );
NAND3X1 NAND3X1_713 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_28_), .B(concatenador_3_nonce_29_), .C(_13468_), .Y(_13479_) );
OAI21X1 OAI21X1_3843 ( .gnd(gnd), .vdd(vdd), .A(_13479_), .B(_13478_), .C(concatenador_3_nonce_31_), .Y(_13480_) );
INVX1 INVX1_905 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_31_), .Y(_13481_) );
NAND3X1 NAND3X1_714 ( .gnd(gnd), .vdd(vdd), .A(concatenador_3_nonce_30_), .B(_13481_), .C(_13475_), .Y(_13482_) );
AOI21X1 AOI21X1_2307 ( .gnd(gnd), .vdd(vdd), .A(_13480_), .B(_13482_), .C(_13485_), .Y(_13377__31_) );
DFFPOSX1 DFFPOSX1_1826 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_13377__0_), .Q(concatenador_3_nonce_0_) );
DFFPOSX1 DFFPOSX1_1827 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_13377__1_), .Q(concatenador_3_nonce_1_) );
DFFPOSX1 DFFPOSX1_1828 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_13377__2_), .Q(concatenador_3_nonce_2_) );
DFFPOSX1 DFFPOSX1_1829 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_13377__3_), .Q(concatenador_3_nonce_3_) );
DFFPOSX1 DFFPOSX1_1830 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_13377__4_), .Q(concatenador_3_nonce_4_) );
DFFPOSX1 DFFPOSX1_1831 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_13377__5_), .Q(concatenador_3_nonce_5_) );
DFFPOSX1 DFFPOSX1_1832 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_13377__6_), .Q(concatenador_3_nonce_6_) );
DFFPOSX1 DFFPOSX1_1833 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_13377__7_), .Q(concatenador_3_nonce_7_) );
DFFPOSX1 DFFPOSX1_1834 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_13377__8_), .Q(concatenador_3_nonce_8_) );
DFFPOSX1 DFFPOSX1_1835 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_13377__9_), .Q(concatenador_3_nonce_9_) );
DFFPOSX1 DFFPOSX1_1836 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_13377__10_), .Q(concatenador_3_nonce_10_) );
DFFPOSX1 DFFPOSX1_1837 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_13377__11_), .Q(concatenador_3_nonce_11_) );
DFFPOSX1 DFFPOSX1_1838 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_13377__12_), .Q(concatenador_3_nonce_12_) );
DFFPOSX1 DFFPOSX1_1839 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_13377__13_), .Q(concatenador_3_nonce_13_) );
DFFPOSX1 DFFPOSX1_1840 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_13377__14_), .Q(concatenador_3_nonce_14_) );
DFFPOSX1 DFFPOSX1_1841 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_13377__15_), .Q(concatenador_3_nonce_15_) );
DFFPOSX1 DFFPOSX1_1842 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_13377__16_), .Q(concatenador_3_nonce_16_) );
DFFPOSX1 DFFPOSX1_1843 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_13377__17_), .Q(concatenador_3_nonce_17_) );
DFFPOSX1 DFFPOSX1_1844 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_13377__18_), .Q(concatenador_3_nonce_18_) );
DFFPOSX1 DFFPOSX1_1845 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_13377__19_), .Q(concatenador_3_nonce_19_) );
DFFPOSX1 DFFPOSX1_1846 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_13377__20_), .Q(concatenador_3_nonce_20_) );
DFFPOSX1 DFFPOSX1_1847 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_13377__21_), .Q(concatenador_3_nonce_21_) );
DFFPOSX1 DFFPOSX1_1848 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_13377__22_), .Q(concatenador_3_nonce_22_) );
DFFPOSX1 DFFPOSX1_1849 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_13377__23_), .Q(concatenador_3_nonce_23_) );
DFFPOSX1 DFFPOSX1_1850 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_13377__24_), .Q(concatenador_3_nonce_24_) );
DFFPOSX1 DFFPOSX1_1851 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_13377__25_), .Q(concatenador_3_nonce_25_) );
DFFPOSX1 DFFPOSX1_1852 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_13377__26_), .Q(concatenador_3_nonce_26_) );
DFFPOSX1 DFFPOSX1_1853 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_13377__27_), .Q(concatenador_3_nonce_27_) );
DFFPOSX1 DFFPOSX1_1854 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_13377__28_), .Q(concatenador_3_nonce_28_) );
DFFPOSX1 DFFPOSX1_1855 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_13377__29_), .Q(concatenador_3_nonce_29_) );
DFFPOSX1 DFFPOSX1_1856 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_13377__30_), .Q(concatenador_3_nonce_30_) );
DFFPOSX1 DFFPOSX1_1857 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_13377__31_), .Q(concatenador_3_nonce_31_) );
INVX1 INVX1_906 ( .gnd(gnd), .vdd(vdd), .A(comparador_valid_bF_buf4), .Y(_13529_) );
NAND2X1 NAND2X1_1843 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf0), .B(_13529_), .Y(_13508_) );
NAND3X1 NAND3X1_715 ( .gnd(gnd), .vdd(vdd), .A(comparador_valid_bF_buf3), .B(reset_bF_buf10), .C(concatenador_nonce_0_), .Y(_13530_) );
INVX1 INVX1_907 ( .gnd(gnd), .vdd(vdd), .A(_13530_), .Y(_13509__0_) );
NAND3X1 NAND3X1_716 ( .gnd(gnd), .vdd(vdd), .A(comparador_valid_bF_buf2), .B(reset_bF_buf9), .C(concatenador_nonce_1_), .Y(_13531_) );
INVX1 INVX1_908 ( .gnd(gnd), .vdd(vdd), .A(_13531_), .Y(_13509__1_) );
NAND3X1 NAND3X1_717 ( .gnd(gnd), .vdd(vdd), .A(comparador_valid_bF_buf1), .B(reset_bF_buf8), .C(concatenador_nonce_2_), .Y(_13532_) );
INVX1 INVX1_909 ( .gnd(gnd), .vdd(vdd), .A(_13532_), .Y(_13509__2_) );
NAND3X1 NAND3X1_718 ( .gnd(gnd), .vdd(vdd), .A(comparador_valid_bF_buf0), .B(reset_bF_buf7), .C(concatenador_nonce_3_), .Y(_13533_) );
INVX1 INVX1_910 ( .gnd(gnd), .vdd(vdd), .A(_13533_), .Y(_13509__3_) );
NAND3X1 NAND3X1_719 ( .gnd(gnd), .vdd(vdd), .A(comparador_valid_bF_buf4), .B(reset_bF_buf6), .C(concatenador_nonce_4_), .Y(_13534_) );
INVX1 INVX1_911 ( .gnd(gnd), .vdd(vdd), .A(_13534_), .Y(_13509__4_) );
NAND3X1 NAND3X1_720 ( .gnd(gnd), .vdd(vdd), .A(comparador_valid_bF_buf3), .B(reset_bF_buf5), .C(concatenador_nonce_5_), .Y(_13535_) );
INVX1 INVX1_912 ( .gnd(gnd), .vdd(vdd), .A(_13535_), .Y(_13509__5_) );
NAND3X1 NAND3X1_721 ( .gnd(gnd), .vdd(vdd), .A(comparador_valid_bF_buf2), .B(reset_bF_buf4), .C(concatenador_nonce_6_), .Y(_13536_) );
INVX1 INVX1_913 ( .gnd(gnd), .vdd(vdd), .A(_13536_), .Y(_13509__6_) );
NAND3X1 NAND3X1_722 ( .gnd(gnd), .vdd(vdd), .A(comparador_valid_bF_buf1), .B(reset_bF_buf3), .C(concatenador_nonce_7_), .Y(_13537_) );
INVX1 INVX1_914 ( .gnd(gnd), .vdd(vdd), .A(_13537_), .Y(_13509__7_) );
NAND3X1 NAND3X1_723 ( .gnd(gnd), .vdd(vdd), .A(comparador_valid_bF_buf0), .B(reset_bF_buf2), .C(concatenador_nonce_8_), .Y(_13538_) );
INVX1 INVX1_915 ( .gnd(gnd), .vdd(vdd), .A(_13538_), .Y(_13509__8_) );
NAND3X1 NAND3X1_724 ( .gnd(gnd), .vdd(vdd), .A(comparador_valid_bF_buf4), .B(reset_bF_buf1), .C(concatenador_nonce_9_), .Y(_13539_) );
INVX1 INVX1_916 ( .gnd(gnd), .vdd(vdd), .A(_13539_), .Y(_13509__9_) );
NAND3X1 NAND3X1_725 ( .gnd(gnd), .vdd(vdd), .A(comparador_valid_bF_buf3), .B(reset_bF_buf0), .C(concatenador_nonce_10_), .Y(_13540_) );
INVX1 INVX1_917 ( .gnd(gnd), .vdd(vdd), .A(_13540_), .Y(_13509__10_) );
NAND3X1 NAND3X1_726 ( .gnd(gnd), .vdd(vdd), .A(comparador_valid_bF_buf2), .B(reset_bF_buf10), .C(concatenador_nonce_11_), .Y(_13541_) );
INVX1 INVX1_918 ( .gnd(gnd), .vdd(vdd), .A(_13541_), .Y(_13509__11_) );
NAND3X1 NAND3X1_727 ( .gnd(gnd), .vdd(vdd), .A(comparador_valid_bF_buf1), .B(reset_bF_buf9), .C(concatenador_nonce_12_), .Y(_13542_) );
INVX1 INVX1_919 ( .gnd(gnd), .vdd(vdd), .A(_13542_), .Y(_13509__12_) );
NAND3X1 NAND3X1_728 ( .gnd(gnd), .vdd(vdd), .A(comparador_valid_bF_buf0), .B(reset_bF_buf8), .C(concatenador_nonce_13_), .Y(_13510_) );
INVX1 INVX1_920 ( .gnd(gnd), .vdd(vdd), .A(_13510_), .Y(_13509__13_) );
NAND3X1 NAND3X1_729 ( .gnd(gnd), .vdd(vdd), .A(comparador_valid_bF_buf4), .B(reset_bF_buf7), .C(concatenador_nonce_14_), .Y(_13511_) );
INVX1 INVX1_921 ( .gnd(gnd), .vdd(vdd), .A(_13511_), .Y(_13509__14_) );
NAND3X1 NAND3X1_730 ( .gnd(gnd), .vdd(vdd), .A(comparador_valid_bF_buf3), .B(reset_bF_buf6), .C(concatenador_nonce_15_), .Y(_13512_) );
INVX1 INVX1_922 ( .gnd(gnd), .vdd(vdd), .A(_13512_), .Y(_13509__15_) );
NAND3X1 NAND3X1_731 ( .gnd(gnd), .vdd(vdd), .A(comparador_valid_bF_buf2), .B(reset_bF_buf5), .C(concatenador_nonce_16_), .Y(_13513_) );
INVX1 INVX1_923 ( .gnd(gnd), .vdd(vdd), .A(_13513_), .Y(_13509__16_) );
NAND3X1 NAND3X1_732 ( .gnd(gnd), .vdd(vdd), .A(comparador_valid_bF_buf1), .B(reset_bF_buf4), .C(concatenador_nonce_17_), .Y(_13514_) );
INVX1 INVX1_924 ( .gnd(gnd), .vdd(vdd), .A(_13514_), .Y(_13509__17_) );
NAND3X1 NAND3X1_733 ( .gnd(gnd), .vdd(vdd), .A(comparador_valid_bF_buf0), .B(reset_bF_buf3), .C(concatenador_nonce_18_), .Y(_13515_) );
INVX1 INVX1_925 ( .gnd(gnd), .vdd(vdd), .A(_13515_), .Y(_13509__18_) );
NAND3X1 NAND3X1_734 ( .gnd(gnd), .vdd(vdd), .A(comparador_valid_bF_buf4), .B(reset_bF_buf2), .C(concatenador_nonce_19_), .Y(_13516_) );
INVX1 INVX1_926 ( .gnd(gnd), .vdd(vdd), .A(_13516_), .Y(_13509__19_) );
NAND3X1 NAND3X1_735 ( .gnd(gnd), .vdd(vdd), .A(comparador_valid_bF_buf3), .B(reset_bF_buf1), .C(concatenador_nonce_20_), .Y(_13517_) );
INVX1 INVX1_927 ( .gnd(gnd), .vdd(vdd), .A(_13517_), .Y(_13509__20_) );
NAND3X1 NAND3X1_736 ( .gnd(gnd), .vdd(vdd), .A(comparador_valid_bF_buf2), .B(reset_bF_buf0), .C(concatenador_nonce_21_), .Y(_13518_) );
INVX1 INVX1_928 ( .gnd(gnd), .vdd(vdd), .A(_13518_), .Y(_13509__21_) );
NAND3X1 NAND3X1_737 ( .gnd(gnd), .vdd(vdd), .A(comparador_valid_bF_buf1), .B(reset_bF_buf10), .C(concatenador_nonce_22_), .Y(_13519_) );
INVX1 INVX1_929 ( .gnd(gnd), .vdd(vdd), .A(_13519_), .Y(_13509__22_) );
NAND3X1 NAND3X1_738 ( .gnd(gnd), .vdd(vdd), .A(comparador_valid_bF_buf0), .B(reset_bF_buf9), .C(concatenador_nonce_23_), .Y(_13520_) );
INVX1 INVX1_930 ( .gnd(gnd), .vdd(vdd), .A(_13520_), .Y(_13509__23_) );
NAND3X1 NAND3X1_739 ( .gnd(gnd), .vdd(vdd), .A(comparador_valid_bF_buf4), .B(reset_bF_buf8), .C(concatenador_nonce_24_), .Y(_13521_) );
INVX1 INVX1_931 ( .gnd(gnd), .vdd(vdd), .A(_13521_), .Y(_13509__24_) );
NAND3X1 NAND3X1_740 ( .gnd(gnd), .vdd(vdd), .A(comparador_valid_bF_buf3), .B(reset_bF_buf7), .C(concatenador_nonce_25_), .Y(_13522_) );
INVX1 INVX1_932 ( .gnd(gnd), .vdd(vdd), .A(_13522_), .Y(_13509__25_) );
NAND3X1 NAND3X1_741 ( .gnd(gnd), .vdd(vdd), .A(comparador_valid_bF_buf2), .B(reset_bF_buf6), .C(concatenador_nonce_26_), .Y(_13523_) );
INVX1 INVX1_933 ( .gnd(gnd), .vdd(vdd), .A(_13523_), .Y(_13509__26_) );
NAND3X1 NAND3X1_742 ( .gnd(gnd), .vdd(vdd), .A(comparador_valid_bF_buf1), .B(reset_bF_buf5), .C(concatenador_nonce_27_), .Y(_13524_) );
INVX1 INVX1_934 ( .gnd(gnd), .vdd(vdd), .A(_13524_), .Y(_13509__27_) );
NAND3X1 NAND3X1_743 ( .gnd(gnd), .vdd(vdd), .A(comparador_valid_bF_buf0), .B(reset_bF_buf4), .C(concatenador_nonce_28_), .Y(_13525_) );
INVX1 INVX1_935 ( .gnd(gnd), .vdd(vdd), .A(_13525_), .Y(_13509__28_) );
NAND3X1 NAND3X1_744 ( .gnd(gnd), .vdd(vdd), .A(comparador_valid_bF_buf4), .B(reset_bF_buf3), .C(concatenador_nonce_29_), .Y(_13526_) );
INVX1 INVX1_936 ( .gnd(gnd), .vdd(vdd), .A(_13526_), .Y(_13509__29_) );
NAND3X1 NAND3X1_745 ( .gnd(gnd), .vdd(vdd), .A(comparador_valid_bF_buf3), .B(reset_bF_buf2), .C(concatenador_nonce_30_), .Y(_13527_) );
INVX1 INVX1_937 ( .gnd(gnd), .vdd(vdd), .A(_13527_), .Y(_13509__30_) );
NAND3X1 NAND3X1_746 ( .gnd(gnd), .vdd(vdd), .A(comparador_valid_bF_buf2), .B(reset_bF_buf1), .C(concatenador_nonce_31_), .Y(_13528_) );
INVX1 INVX1_938 ( .gnd(gnd), .vdd(vdd), .A(_13528_), .Y(_13509__31_) );
DFFPOSX1 DFFPOSX1_1858 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_13509__0_), .Q(nonce_out_1_0_) );
DFFPOSX1 DFFPOSX1_1859 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_13509__1_), .Q(nonce_out_1_1_) );
DFFPOSX1 DFFPOSX1_1860 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_13509__2_), .Q(nonce_out_1_2_) );
DFFPOSX1 DFFPOSX1_1861 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_13509__3_), .Q(nonce_out_1_3_) );
DFFPOSX1 DFFPOSX1_1862 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_13509__4_), .Q(nonce_out_1_4_) );
DFFPOSX1 DFFPOSX1_1863 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_13509__5_), .Q(nonce_out_1_5_) );
DFFPOSX1 DFFPOSX1_1864 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_13509__6_), .Q(nonce_out_1_6_) );
DFFPOSX1 DFFPOSX1_1865 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_13509__7_), .Q(nonce_out_1_7_) );
DFFPOSX1 DFFPOSX1_1866 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_13509__8_), .Q(nonce_out_1_8_) );
DFFPOSX1 DFFPOSX1_1867 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_13509__9_), .Q(nonce_out_1_9_) );
DFFPOSX1 DFFPOSX1_1868 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_13509__10_), .Q(nonce_out_1_10_) );
DFFPOSX1 DFFPOSX1_1869 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_13509__11_), .Q(nonce_out_1_11_) );
DFFPOSX1 DFFPOSX1_1870 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_13509__12_), .Q(nonce_out_1_12_) );
DFFPOSX1 DFFPOSX1_1871 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_13509__13_), .Q(nonce_out_1_13_) );
DFFPOSX1 DFFPOSX1_1872 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_13509__14_), .Q(nonce_out_1_14_) );
DFFPOSX1 DFFPOSX1_1873 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_13509__15_), .Q(nonce_out_1_15_) );
DFFPOSX1 DFFPOSX1_1874 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_13509__16_), .Q(nonce_out_1_16_) );
DFFPOSX1 DFFPOSX1_1875 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_13509__17_), .Q(nonce_out_1_17_) );
DFFPOSX1 DFFPOSX1_1876 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_13509__18_), .Q(nonce_out_1_18_) );
DFFPOSX1 DFFPOSX1_1877 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_13509__19_), .Q(nonce_out_1_19_) );
DFFPOSX1 DFFPOSX1_1878 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_13509__20_), .Q(nonce_out_1_20_) );
DFFPOSX1 DFFPOSX1_1879 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_13509__21_), .Q(nonce_out_1_21_) );
DFFPOSX1 DFFPOSX1_1880 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_13509__22_), .Q(nonce_out_1_22_) );
DFFPOSX1 DFFPOSX1_1881 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_13509__23_), .Q(nonce_out_1_23_) );
DFFPOSX1 DFFPOSX1_1882 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_13509__24_), .Q(nonce_out_1_24_) );
DFFPOSX1 DFFPOSX1_1883 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_13509__25_), .Q(nonce_out_1_25_) );
DFFPOSX1 DFFPOSX1_1884 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_13509__26_), .Q(nonce_out_1_26_) );
DFFPOSX1 DFFPOSX1_1885 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_13509__27_), .Q(nonce_out_1_27_) );
DFFPOSX1 DFFPOSX1_1886 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_13509__28_), .Q(nonce_out_1_28_) );
DFFPOSX1 DFFPOSX1_1887 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_13509__29_), .Q(nonce_out_1_29_) );
DFFPOSX1 DFFPOSX1_1888 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_13509__30_), .Q(nonce_out_1_30_) );
DFFPOSX1 DFFPOSX1_1889 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_13509__31_), .Q(nonce_out_1_31_) );
DFFPOSX1 DFFPOSX1_1890 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_13508_), .Q(finished_1) );
INVX1 INVX1_939 ( .gnd(gnd), .vdd(vdd), .A(comparador_2_valid_bF_buf4), .Y(_13564_) );
NAND2X1 NAND2X1_1844 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf0), .B(_13564_), .Y(_13543_) );
NAND3X1 NAND3X1_747 ( .gnd(gnd), .vdd(vdd), .A(comparador_2_valid_bF_buf3), .B(reset_bF_buf10), .C(concatenador_2_nonce_0_), .Y(_13565_) );
INVX1 INVX1_940 ( .gnd(gnd), .vdd(vdd), .A(_13565_), .Y(_13544__0_) );
NAND3X1 NAND3X1_748 ( .gnd(gnd), .vdd(vdd), .A(comparador_2_valid_bF_buf2), .B(reset_bF_buf9), .C(concatenador_2_nonce_1_), .Y(_13566_) );
INVX1 INVX1_941 ( .gnd(gnd), .vdd(vdd), .A(_13566_), .Y(_13544__1_) );
NAND3X1 NAND3X1_749 ( .gnd(gnd), .vdd(vdd), .A(comparador_2_valid_bF_buf1), .B(reset_bF_buf8), .C(concatenador_2_nonce_2_), .Y(_13567_) );
INVX1 INVX1_942 ( .gnd(gnd), .vdd(vdd), .A(_13567_), .Y(_13544__2_) );
NAND3X1 NAND3X1_750 ( .gnd(gnd), .vdd(vdd), .A(comparador_2_valid_bF_buf0), .B(reset_bF_buf7), .C(concatenador_2_nonce_3_), .Y(_13568_) );
INVX1 INVX1_943 ( .gnd(gnd), .vdd(vdd), .A(_13568_), .Y(_13544__3_) );
NAND3X1 NAND3X1_751 ( .gnd(gnd), .vdd(vdd), .A(comparador_2_valid_bF_buf4), .B(reset_bF_buf6), .C(concatenador_2_nonce_4_), .Y(_13569_) );
INVX1 INVX1_944 ( .gnd(gnd), .vdd(vdd), .A(_13569_), .Y(_13544__4_) );
NAND3X1 NAND3X1_752 ( .gnd(gnd), .vdd(vdd), .A(comparador_2_valid_bF_buf3), .B(reset_bF_buf5), .C(concatenador_2_nonce_5_), .Y(_13570_) );
INVX1 INVX1_945 ( .gnd(gnd), .vdd(vdd), .A(_13570_), .Y(_13544__5_) );
NAND3X1 NAND3X1_753 ( .gnd(gnd), .vdd(vdd), .A(comparador_2_valid_bF_buf2), .B(reset_bF_buf4), .C(concatenador_2_nonce_6_), .Y(_13571_) );
INVX1 INVX1_946 ( .gnd(gnd), .vdd(vdd), .A(_13571_), .Y(_13544__6_) );
NAND3X1 NAND3X1_754 ( .gnd(gnd), .vdd(vdd), .A(comparador_2_valid_bF_buf1), .B(reset_bF_buf3), .C(concatenador_2_nonce_7_), .Y(_13572_) );
INVX1 INVX1_947 ( .gnd(gnd), .vdd(vdd), .A(_13572_), .Y(_13544__7_) );
NAND3X1 NAND3X1_755 ( .gnd(gnd), .vdd(vdd), .A(comparador_2_valid_bF_buf0), .B(reset_bF_buf2), .C(concatenador_2_nonce_8_), .Y(_13573_) );
INVX1 INVX1_948 ( .gnd(gnd), .vdd(vdd), .A(_13573_), .Y(_13544__8_) );
NAND3X1 NAND3X1_756 ( .gnd(gnd), .vdd(vdd), .A(comparador_2_valid_bF_buf4), .B(reset_bF_buf1), .C(concatenador_2_nonce_9_), .Y(_13574_) );
INVX1 INVX1_949 ( .gnd(gnd), .vdd(vdd), .A(_13574_), .Y(_13544__9_) );
NAND3X1 NAND3X1_757 ( .gnd(gnd), .vdd(vdd), .A(comparador_2_valid_bF_buf3), .B(reset_bF_buf0), .C(concatenador_2_nonce_10_), .Y(_13575_) );
INVX1 INVX1_950 ( .gnd(gnd), .vdd(vdd), .A(_13575_), .Y(_13544__10_) );
NAND3X1 NAND3X1_758 ( .gnd(gnd), .vdd(vdd), .A(comparador_2_valid_bF_buf2), .B(reset_bF_buf10), .C(concatenador_2_nonce_11_), .Y(_13576_) );
INVX1 INVX1_951 ( .gnd(gnd), .vdd(vdd), .A(_13576_), .Y(_13544__11_) );
NAND3X1 NAND3X1_759 ( .gnd(gnd), .vdd(vdd), .A(comparador_2_valid_bF_buf1), .B(reset_bF_buf9), .C(concatenador_2_nonce_12_), .Y(_13577_) );
INVX1 INVX1_952 ( .gnd(gnd), .vdd(vdd), .A(_13577_), .Y(_13544__12_) );
NAND3X1 NAND3X1_760 ( .gnd(gnd), .vdd(vdd), .A(comparador_2_valid_bF_buf0), .B(reset_bF_buf8), .C(concatenador_2_nonce_13_), .Y(_13545_) );
INVX1 INVX1_953 ( .gnd(gnd), .vdd(vdd), .A(_13545_), .Y(_13544__13_) );
NAND3X1 NAND3X1_761 ( .gnd(gnd), .vdd(vdd), .A(comparador_2_valid_bF_buf4), .B(reset_bF_buf7), .C(concatenador_2_nonce_14_), .Y(_13546_) );
INVX1 INVX1_954 ( .gnd(gnd), .vdd(vdd), .A(_13546_), .Y(_13544__14_) );
NAND3X1 NAND3X1_762 ( .gnd(gnd), .vdd(vdd), .A(comparador_2_valid_bF_buf3), .B(reset_bF_buf6), .C(concatenador_2_nonce_15_), .Y(_13547_) );
INVX1 INVX1_955 ( .gnd(gnd), .vdd(vdd), .A(_13547_), .Y(_13544__15_) );
NAND3X1 NAND3X1_763 ( .gnd(gnd), .vdd(vdd), .A(comparador_2_valid_bF_buf2), .B(reset_bF_buf5), .C(concatenador_2_nonce_16_), .Y(_13548_) );
INVX1 INVX1_956 ( .gnd(gnd), .vdd(vdd), .A(_13548_), .Y(_13544__16_) );
NAND3X1 NAND3X1_764 ( .gnd(gnd), .vdd(vdd), .A(comparador_2_valid_bF_buf1), .B(reset_bF_buf4), .C(concatenador_2_nonce_17_), .Y(_13549_) );
INVX1 INVX1_957 ( .gnd(gnd), .vdd(vdd), .A(_13549_), .Y(_13544__17_) );
NAND3X1 NAND3X1_765 ( .gnd(gnd), .vdd(vdd), .A(comparador_2_valid_bF_buf0), .B(reset_bF_buf3), .C(concatenador_2_nonce_18_), .Y(_13550_) );
INVX1 INVX1_958 ( .gnd(gnd), .vdd(vdd), .A(_13550_), .Y(_13544__18_) );
NAND3X1 NAND3X1_766 ( .gnd(gnd), .vdd(vdd), .A(comparador_2_valid_bF_buf4), .B(reset_bF_buf2), .C(concatenador_2_nonce_19_), .Y(_13551_) );
INVX1 INVX1_959 ( .gnd(gnd), .vdd(vdd), .A(_13551_), .Y(_13544__19_) );
NAND3X1 NAND3X1_767 ( .gnd(gnd), .vdd(vdd), .A(comparador_2_valid_bF_buf3), .B(reset_bF_buf1), .C(concatenador_2_nonce_20_), .Y(_13552_) );
INVX1 INVX1_960 ( .gnd(gnd), .vdd(vdd), .A(_13552_), .Y(_13544__20_) );
NAND3X1 NAND3X1_768 ( .gnd(gnd), .vdd(vdd), .A(comparador_2_valid_bF_buf2), .B(reset_bF_buf0), .C(concatenador_2_nonce_21_), .Y(_13553_) );
INVX1 INVX1_961 ( .gnd(gnd), .vdd(vdd), .A(_13553_), .Y(_13544__21_) );
NAND3X1 NAND3X1_769 ( .gnd(gnd), .vdd(vdd), .A(comparador_2_valid_bF_buf1), .B(reset_bF_buf10), .C(concatenador_2_nonce_22_), .Y(_13554_) );
INVX1 INVX1_962 ( .gnd(gnd), .vdd(vdd), .A(_13554_), .Y(_13544__22_) );
NAND3X1 NAND3X1_770 ( .gnd(gnd), .vdd(vdd), .A(comparador_2_valid_bF_buf0), .B(reset_bF_buf9), .C(concatenador_2_nonce_23_), .Y(_13555_) );
INVX1 INVX1_963 ( .gnd(gnd), .vdd(vdd), .A(_13555_), .Y(_13544__23_) );
NAND3X1 NAND3X1_771 ( .gnd(gnd), .vdd(vdd), .A(comparador_2_valid_bF_buf4), .B(reset_bF_buf8), .C(concatenador_2_nonce_24_), .Y(_13556_) );
INVX1 INVX1_964 ( .gnd(gnd), .vdd(vdd), .A(_13556_), .Y(_13544__24_) );
NAND3X1 NAND3X1_772 ( .gnd(gnd), .vdd(vdd), .A(comparador_2_valid_bF_buf3), .B(reset_bF_buf7), .C(concatenador_2_nonce_25_), .Y(_13557_) );
INVX1 INVX1_965 ( .gnd(gnd), .vdd(vdd), .A(_13557_), .Y(_13544__25_) );
NAND3X1 NAND3X1_773 ( .gnd(gnd), .vdd(vdd), .A(comparador_2_valid_bF_buf2), .B(reset_bF_buf6), .C(concatenador_2_nonce_26_), .Y(_13558_) );
INVX1 INVX1_966 ( .gnd(gnd), .vdd(vdd), .A(_13558_), .Y(_13544__26_) );
NAND3X1 NAND3X1_774 ( .gnd(gnd), .vdd(vdd), .A(comparador_2_valid_bF_buf1), .B(reset_bF_buf5), .C(concatenador_2_nonce_27_), .Y(_13559_) );
INVX1 INVX1_967 ( .gnd(gnd), .vdd(vdd), .A(_13559_), .Y(_13544__27_) );
NAND3X1 NAND3X1_775 ( .gnd(gnd), .vdd(vdd), .A(comparador_2_valid_bF_buf0), .B(reset_bF_buf4), .C(concatenador_2_nonce_28_), .Y(_13560_) );
INVX1 INVX1_968 ( .gnd(gnd), .vdd(vdd), .A(_13560_), .Y(_13544__28_) );
NAND3X1 NAND3X1_776 ( .gnd(gnd), .vdd(vdd), .A(comparador_2_valid_bF_buf4), .B(reset_bF_buf3), .C(concatenador_2_nonce_29_), .Y(_13561_) );
INVX1 INVX1_969 ( .gnd(gnd), .vdd(vdd), .A(_13561_), .Y(_13544__29_) );
NAND3X1 NAND3X1_777 ( .gnd(gnd), .vdd(vdd), .A(comparador_2_valid_bF_buf3), .B(reset_bF_buf2), .C(concatenador_2_nonce_30_), .Y(_13562_) );
INVX1 INVX1_970 ( .gnd(gnd), .vdd(vdd), .A(_13562_), .Y(_13544__30_) );
NAND3X1 NAND3X1_778 ( .gnd(gnd), .vdd(vdd), .A(comparador_2_valid_bF_buf2), .B(reset_bF_buf1), .C(concatenador_2_nonce_31_), .Y(_13563_) );
INVX1 INVX1_971 ( .gnd(gnd), .vdd(vdd), .A(_13563_), .Y(_13544__31_) );
DFFPOSX1 DFFPOSX1_1891 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_13544__0_), .Q(nonce_out_2_0_) );
DFFPOSX1 DFFPOSX1_1892 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_13544__1_), .Q(nonce_out_2_1_) );
DFFPOSX1 DFFPOSX1_1893 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_13544__2_), .Q(nonce_out_2_2_) );
DFFPOSX1 DFFPOSX1_1894 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_13544__3_), .Q(nonce_out_2_3_) );
DFFPOSX1 DFFPOSX1_1895 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_13544__4_), .Q(nonce_out_2_4_) );
DFFPOSX1 DFFPOSX1_1896 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_13544__5_), .Q(nonce_out_2_5_) );
DFFPOSX1 DFFPOSX1_1897 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf157), .D(_13544__6_), .Q(nonce_out_2_6_) );
DFFPOSX1 DFFPOSX1_1898 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf156), .D(_13544__7_), .Q(nonce_out_2_7_) );
DFFPOSX1 DFFPOSX1_1899 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf155), .D(_13544__8_), .Q(nonce_out_2_8_) );
DFFPOSX1 DFFPOSX1_1900 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf154), .D(_13544__9_), .Q(nonce_out_2_9_) );
DFFPOSX1 DFFPOSX1_1901 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf153), .D(_13544__10_), .Q(nonce_out_2_10_) );
DFFPOSX1 DFFPOSX1_1902 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf152), .D(_13544__11_), .Q(nonce_out_2_11_) );
DFFPOSX1 DFFPOSX1_1903 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf151), .D(_13544__12_), .Q(nonce_out_2_12_) );
DFFPOSX1 DFFPOSX1_1904 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf150), .D(_13544__13_), .Q(nonce_out_2_13_) );
DFFPOSX1 DFFPOSX1_1905 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf149), .D(_13544__14_), .Q(nonce_out_2_14_) );
DFFPOSX1 DFFPOSX1_1906 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf148), .D(_13544__15_), .Q(nonce_out_2_15_) );
DFFPOSX1 DFFPOSX1_1907 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf147), .D(_13544__16_), .Q(nonce_out_2_16_) );
DFFPOSX1 DFFPOSX1_1908 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf146), .D(_13544__17_), .Q(nonce_out_2_17_) );
DFFPOSX1 DFFPOSX1_1909 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf145), .D(_13544__18_), .Q(nonce_out_2_18_) );
DFFPOSX1 DFFPOSX1_1910 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf144), .D(_13544__19_), .Q(nonce_out_2_19_) );
DFFPOSX1 DFFPOSX1_1911 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf143), .D(_13544__20_), .Q(nonce_out_2_20_) );
DFFPOSX1 DFFPOSX1_1912 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf142), .D(_13544__21_), .Q(nonce_out_2_21_) );
DFFPOSX1 DFFPOSX1_1913 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf141), .D(_13544__22_), .Q(nonce_out_2_22_) );
DFFPOSX1 DFFPOSX1_1914 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf140), .D(_13544__23_), .Q(nonce_out_2_23_) );
DFFPOSX1 DFFPOSX1_1915 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf139), .D(_13544__24_), .Q(nonce_out_2_24_) );
DFFPOSX1 DFFPOSX1_1916 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf138), .D(_13544__25_), .Q(nonce_out_2_25_) );
DFFPOSX1 DFFPOSX1_1917 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf137), .D(_13544__26_), .Q(nonce_out_2_26_) );
DFFPOSX1 DFFPOSX1_1918 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf136), .D(_13544__27_), .Q(nonce_out_2_27_) );
DFFPOSX1 DFFPOSX1_1919 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf135), .D(_13544__28_), .Q(nonce_out_2_28_) );
DFFPOSX1 DFFPOSX1_1920 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf134), .D(_13544__29_), .Q(nonce_out_2_29_) );
DFFPOSX1 DFFPOSX1_1921 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf133), .D(_13544__30_), .Q(nonce_out_2_30_) );
DFFPOSX1 DFFPOSX1_1922 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf132), .D(_13544__31_), .Q(nonce_out_2_31_) );
DFFPOSX1 DFFPOSX1_1923 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf131), .D(_13543_), .Q(finished_2) );
INVX1 INVX1_972 ( .gnd(gnd), .vdd(vdd), .A(comparador_3_valid_bF_buf4), .Y(_13599_) );
NAND2X1 NAND2X1_1845 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf0), .B(_13599_), .Y(_13578_) );
NAND3X1 NAND3X1_779 ( .gnd(gnd), .vdd(vdd), .A(comparador_3_valid_bF_buf3), .B(reset_bF_buf10), .C(concatenador_3_nonce_0_), .Y(_13600_) );
INVX1 INVX1_973 ( .gnd(gnd), .vdd(vdd), .A(_13600_), .Y(_13579__0_) );
NAND3X1 NAND3X1_780 ( .gnd(gnd), .vdd(vdd), .A(comparador_3_valid_bF_buf2), .B(reset_bF_buf9), .C(concatenador_3_nonce_1_), .Y(_13601_) );
INVX1 INVX1_974 ( .gnd(gnd), .vdd(vdd), .A(_13601_), .Y(_13579__1_) );
NAND3X1 NAND3X1_781 ( .gnd(gnd), .vdd(vdd), .A(comparador_3_valid_bF_buf1), .B(reset_bF_buf8), .C(concatenador_3_nonce_2_), .Y(_13602_) );
INVX1 INVX1_975 ( .gnd(gnd), .vdd(vdd), .A(_13602_), .Y(_13579__2_) );
NAND3X1 NAND3X1_782 ( .gnd(gnd), .vdd(vdd), .A(comparador_3_valid_bF_buf0), .B(reset_bF_buf7), .C(concatenador_3_nonce_3_), .Y(_13603_) );
INVX1 INVX1_976 ( .gnd(gnd), .vdd(vdd), .A(_13603_), .Y(_13579__3_) );
NAND3X1 NAND3X1_783 ( .gnd(gnd), .vdd(vdd), .A(comparador_3_valid_bF_buf4), .B(reset_bF_buf6), .C(concatenador_3_nonce_4_), .Y(_13604_) );
INVX1 INVX1_977 ( .gnd(gnd), .vdd(vdd), .A(_13604_), .Y(_13579__4_) );
NAND3X1 NAND3X1_784 ( .gnd(gnd), .vdd(vdd), .A(comparador_3_valid_bF_buf3), .B(reset_bF_buf5), .C(concatenador_3_nonce_5_), .Y(_13605_) );
INVX1 INVX1_978 ( .gnd(gnd), .vdd(vdd), .A(_13605_), .Y(_13579__5_) );
NAND3X1 NAND3X1_785 ( .gnd(gnd), .vdd(vdd), .A(comparador_3_valid_bF_buf2), .B(reset_bF_buf4), .C(concatenador_3_nonce_6_), .Y(_13606_) );
INVX1 INVX1_979 ( .gnd(gnd), .vdd(vdd), .A(_13606_), .Y(_13579__6_) );
NAND3X1 NAND3X1_786 ( .gnd(gnd), .vdd(vdd), .A(comparador_3_valid_bF_buf1), .B(reset_bF_buf3), .C(concatenador_3_nonce_7_), .Y(_13607_) );
INVX1 INVX1_980 ( .gnd(gnd), .vdd(vdd), .A(_13607_), .Y(_13579__7_) );
NAND3X1 NAND3X1_787 ( .gnd(gnd), .vdd(vdd), .A(comparador_3_valid_bF_buf0), .B(reset_bF_buf2), .C(concatenador_3_nonce_8_), .Y(_13608_) );
INVX1 INVX1_981 ( .gnd(gnd), .vdd(vdd), .A(_13608_), .Y(_13579__8_) );
NAND3X1 NAND3X1_788 ( .gnd(gnd), .vdd(vdd), .A(comparador_3_valid_bF_buf4), .B(reset_bF_buf1), .C(concatenador_3_nonce_9_), .Y(_13609_) );
INVX1 INVX1_982 ( .gnd(gnd), .vdd(vdd), .A(_13609_), .Y(_13579__9_) );
NAND3X1 NAND3X1_789 ( .gnd(gnd), .vdd(vdd), .A(comparador_3_valid_bF_buf3), .B(reset_bF_buf0), .C(concatenador_3_nonce_10_), .Y(_13610_) );
INVX1 INVX1_983 ( .gnd(gnd), .vdd(vdd), .A(_13610_), .Y(_13579__10_) );
NAND3X1 NAND3X1_790 ( .gnd(gnd), .vdd(vdd), .A(comparador_3_valid_bF_buf2), .B(reset_bF_buf10), .C(concatenador_3_nonce_11_), .Y(_13611_) );
INVX1 INVX1_984 ( .gnd(gnd), .vdd(vdd), .A(_13611_), .Y(_13579__11_) );
NAND3X1 NAND3X1_791 ( .gnd(gnd), .vdd(vdd), .A(comparador_3_valid_bF_buf1), .B(reset_bF_buf9), .C(concatenador_3_nonce_12_), .Y(_13612_) );
INVX1 INVX1_985 ( .gnd(gnd), .vdd(vdd), .A(_13612_), .Y(_13579__12_) );
NAND3X1 NAND3X1_792 ( .gnd(gnd), .vdd(vdd), .A(comparador_3_valid_bF_buf0), .B(reset_bF_buf8), .C(concatenador_3_nonce_13_), .Y(_13580_) );
INVX1 INVX1_986 ( .gnd(gnd), .vdd(vdd), .A(_13580_), .Y(_13579__13_) );
NAND3X1 NAND3X1_793 ( .gnd(gnd), .vdd(vdd), .A(comparador_3_valid_bF_buf4), .B(reset_bF_buf7), .C(concatenador_3_nonce_14_), .Y(_13581_) );
INVX1 INVX1_987 ( .gnd(gnd), .vdd(vdd), .A(_13581_), .Y(_13579__14_) );
NAND3X1 NAND3X1_794 ( .gnd(gnd), .vdd(vdd), .A(comparador_3_valid_bF_buf3), .B(reset_bF_buf6), .C(concatenador_3_nonce_15_), .Y(_13582_) );
INVX1 INVX1_988 ( .gnd(gnd), .vdd(vdd), .A(_13582_), .Y(_13579__15_) );
NAND3X1 NAND3X1_795 ( .gnd(gnd), .vdd(vdd), .A(comparador_3_valid_bF_buf2), .B(reset_bF_buf5), .C(concatenador_3_nonce_16_), .Y(_13583_) );
INVX1 INVX1_989 ( .gnd(gnd), .vdd(vdd), .A(_13583_), .Y(_13579__16_) );
NAND3X1 NAND3X1_796 ( .gnd(gnd), .vdd(vdd), .A(comparador_3_valid_bF_buf1), .B(reset_bF_buf4), .C(concatenador_3_nonce_17_), .Y(_13584_) );
INVX1 INVX1_990 ( .gnd(gnd), .vdd(vdd), .A(_13584_), .Y(_13579__17_) );
NAND3X1 NAND3X1_797 ( .gnd(gnd), .vdd(vdd), .A(comparador_3_valid_bF_buf0), .B(reset_bF_buf3), .C(concatenador_3_nonce_18_), .Y(_13585_) );
INVX1 INVX1_991 ( .gnd(gnd), .vdd(vdd), .A(_13585_), .Y(_13579__18_) );
NAND3X1 NAND3X1_798 ( .gnd(gnd), .vdd(vdd), .A(comparador_3_valid_bF_buf4), .B(reset_bF_buf2), .C(concatenador_3_nonce_19_), .Y(_13586_) );
INVX1 INVX1_992 ( .gnd(gnd), .vdd(vdd), .A(_13586_), .Y(_13579__19_) );
NAND3X1 NAND3X1_799 ( .gnd(gnd), .vdd(vdd), .A(comparador_3_valid_bF_buf3), .B(reset_bF_buf1), .C(concatenador_3_nonce_20_), .Y(_13587_) );
INVX1 INVX1_993 ( .gnd(gnd), .vdd(vdd), .A(_13587_), .Y(_13579__20_) );
NAND3X1 NAND3X1_800 ( .gnd(gnd), .vdd(vdd), .A(comparador_3_valid_bF_buf2), .B(reset_bF_buf0), .C(concatenador_3_nonce_21_), .Y(_13588_) );
INVX1 INVX1_994 ( .gnd(gnd), .vdd(vdd), .A(_13588_), .Y(_13579__21_) );
NAND3X1 NAND3X1_801 ( .gnd(gnd), .vdd(vdd), .A(comparador_3_valid_bF_buf1), .B(reset_bF_buf10), .C(concatenador_3_nonce_22_), .Y(_13589_) );
INVX1 INVX1_995 ( .gnd(gnd), .vdd(vdd), .A(_13589_), .Y(_13579__22_) );
NAND3X1 NAND3X1_802 ( .gnd(gnd), .vdd(vdd), .A(comparador_3_valid_bF_buf0), .B(reset_bF_buf9), .C(concatenador_3_nonce_23_), .Y(_13590_) );
INVX1 INVX1_996 ( .gnd(gnd), .vdd(vdd), .A(_13590_), .Y(_13579__23_) );
NAND3X1 NAND3X1_803 ( .gnd(gnd), .vdd(vdd), .A(comparador_3_valid_bF_buf4), .B(reset_bF_buf8), .C(concatenador_3_nonce_24_), .Y(_13591_) );
INVX1 INVX1_997 ( .gnd(gnd), .vdd(vdd), .A(_13591_), .Y(_13579__24_) );
NAND3X1 NAND3X1_804 ( .gnd(gnd), .vdd(vdd), .A(comparador_3_valid_bF_buf3), .B(reset_bF_buf7), .C(concatenador_3_nonce_25_), .Y(_13592_) );
INVX1 INVX1_998 ( .gnd(gnd), .vdd(vdd), .A(_13592_), .Y(_13579__25_) );
NAND3X1 NAND3X1_805 ( .gnd(gnd), .vdd(vdd), .A(comparador_3_valid_bF_buf2), .B(reset_bF_buf6), .C(concatenador_3_nonce_26_), .Y(_13593_) );
INVX1 INVX1_999 ( .gnd(gnd), .vdd(vdd), .A(_13593_), .Y(_13579__26_) );
NAND3X1 NAND3X1_806 ( .gnd(gnd), .vdd(vdd), .A(comparador_3_valid_bF_buf1), .B(reset_bF_buf5), .C(concatenador_3_nonce_27_), .Y(_13594_) );
INVX1 INVX1_1000 ( .gnd(gnd), .vdd(vdd), .A(_13594_), .Y(_13579__27_) );
NAND3X1 NAND3X1_807 ( .gnd(gnd), .vdd(vdd), .A(comparador_3_valid_bF_buf0), .B(reset_bF_buf4), .C(concatenador_3_nonce_28_), .Y(_13595_) );
INVX1 INVX1_1001 ( .gnd(gnd), .vdd(vdd), .A(_13595_), .Y(_13579__28_) );
NAND3X1 NAND3X1_808 ( .gnd(gnd), .vdd(vdd), .A(comparador_3_valid_bF_buf4), .B(reset_bF_buf3), .C(concatenador_3_nonce_29_), .Y(_13596_) );
INVX1 INVX1_1002 ( .gnd(gnd), .vdd(vdd), .A(_13596_), .Y(_13579__29_) );
NAND3X1 NAND3X1_809 ( .gnd(gnd), .vdd(vdd), .A(comparador_3_valid_bF_buf3), .B(reset_bF_buf2), .C(concatenador_3_nonce_30_), .Y(_13597_) );
INVX1 INVX1_1003 ( .gnd(gnd), .vdd(vdd), .A(_13597_), .Y(_13579__30_) );
NAND3X1 NAND3X1_810 ( .gnd(gnd), .vdd(vdd), .A(comparador_3_valid_bF_buf2), .B(reset_bF_buf1), .C(concatenador_3_nonce_31_), .Y(_13598_) );
INVX1 INVX1_1004 ( .gnd(gnd), .vdd(vdd), .A(_13598_), .Y(_13579__31_) );
DFFPOSX1 DFFPOSX1_1924 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf130), .D(_13579__0_), .Q(nonce_out_3_0_) );
DFFPOSX1 DFFPOSX1_1925 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf129), .D(_13579__1_), .Q(nonce_out_3_1_) );
DFFPOSX1 DFFPOSX1_1926 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf128), .D(_13579__2_), .Q(nonce_out_3_2_) );
DFFPOSX1 DFFPOSX1_1927 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf127), .D(_13579__3_), .Q(nonce_out_3_3_) );
DFFPOSX1 DFFPOSX1_1928 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf126), .D(_13579__4_), .Q(nonce_out_3_4_) );
DFFPOSX1 DFFPOSX1_1929 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf125), .D(_13579__5_), .Q(nonce_out_3_5_) );
DFFPOSX1 DFFPOSX1_1930 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf124), .D(_13579__6_), .Q(nonce_out_3_6_) );
DFFPOSX1 DFFPOSX1_1931 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf123), .D(_13579__7_), .Q(nonce_out_3_7_) );
DFFPOSX1 DFFPOSX1_1932 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf122), .D(_13579__8_), .Q(nonce_out_3_8_) );
DFFPOSX1 DFFPOSX1_1933 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf121), .D(_13579__9_), .Q(nonce_out_3_9_) );
DFFPOSX1 DFFPOSX1_1934 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf120), .D(_13579__10_), .Q(nonce_out_3_10_) );
DFFPOSX1 DFFPOSX1_1935 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf119), .D(_13579__11_), .Q(nonce_out_3_11_) );
DFFPOSX1 DFFPOSX1_1936 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf118), .D(_13579__12_), .Q(nonce_out_3_12_) );
DFFPOSX1 DFFPOSX1_1937 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf117), .D(_13579__13_), .Q(nonce_out_3_13_) );
DFFPOSX1 DFFPOSX1_1938 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf116), .D(_13579__14_), .Q(nonce_out_3_14_) );
DFFPOSX1 DFFPOSX1_1939 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf115), .D(_13579__15_), .Q(nonce_out_3_15_) );
DFFPOSX1 DFFPOSX1_1940 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf114), .D(_13579__16_), .Q(nonce_out_3_16_) );
DFFPOSX1 DFFPOSX1_1941 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf113), .D(_13579__17_), .Q(nonce_out_3_17_) );
DFFPOSX1 DFFPOSX1_1942 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf112), .D(_13579__18_), .Q(nonce_out_3_18_) );
DFFPOSX1 DFFPOSX1_1943 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf111), .D(_13579__19_), .Q(nonce_out_3_19_) );
DFFPOSX1 DFFPOSX1_1944 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf110), .D(_13579__20_), .Q(nonce_out_3_20_) );
DFFPOSX1 DFFPOSX1_1945 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf109), .D(_13579__21_), .Q(nonce_out_3_21_) );
DFFPOSX1 DFFPOSX1_1946 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf108), .D(_13579__22_), .Q(nonce_out_3_22_) );
DFFPOSX1 DFFPOSX1_1947 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf107), .D(_13579__23_), .Q(nonce_out_3_23_) );
DFFPOSX1 DFFPOSX1_1948 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(_13579__24_), .Q(nonce_out_3_24_) );
DFFPOSX1 DFFPOSX1_1949 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(_13579__25_), .Q(nonce_out_3_25_) );
DFFPOSX1 DFFPOSX1_1950 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(_13579__26_), .Q(nonce_out_3_26_) );
DFFPOSX1 DFFPOSX1_1951 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(_13579__27_), .Q(nonce_out_3_27_) );
DFFPOSX1 DFFPOSX1_1952 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(_13579__28_), .Q(nonce_out_3_28_) );
DFFPOSX1 DFFPOSX1_1953 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(_13579__29_), .Q(nonce_out_3_29_) );
DFFPOSX1 DFFPOSX1_1954 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(_13579__30_), .Q(nonce_out_3_30_) );
DFFPOSX1 DFFPOSX1_1955 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(_13579__31_), .Q(nonce_out_3_31_) );
DFFPOSX1 DFFPOSX1_1956 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_13578_), .Q(finished_3) );
INVX8 INVX8_288 ( .gnd(gnd), .vdd(vdd), .A(finished_2_bF_buf4), .Y(_13615_) );
NAND3X1 NAND3X1_811 ( .gnd(gnd), .vdd(vdd), .A(finished_3_bF_buf4), .B(nonce_out_3_0_), .C(_13615__bF_buf4), .Y(_13616_) );
AOI21X1 AOI21X1_2308 ( .gnd(gnd), .vdd(vdd), .A(nonce_out_2_0_), .B(finished_2_bF_buf3), .C(finished_1_bF_buf4), .Y(_13617_) );
INVX8 INVX8_289 ( .gnd(gnd), .vdd(vdd), .A(finished_1_bF_buf3), .Y(_13618_) );
OAI21X1 OAI21X1_3844 ( .gnd(gnd), .vdd(vdd), .A(_13618__bF_buf4), .B(nonce_out_1_0_), .C(reset_bF_buf0), .Y(_13619_) );
AOI21X1 AOI21X1_2309 ( .gnd(gnd), .vdd(vdd), .A(_13617_), .B(_13616_), .C(_13619_), .Y(_13614__0_) );
NAND3X1 NAND3X1_812 ( .gnd(gnd), .vdd(vdd), .A(finished_3_bF_buf3), .B(nonce_out_3_1_), .C(_13615__bF_buf3), .Y(_13620_) );
AOI21X1 AOI21X1_2310 ( .gnd(gnd), .vdd(vdd), .A(finished_2_bF_buf2), .B(nonce_out_2_1_), .C(finished_1_bF_buf2), .Y(_13621_) );
OAI21X1 OAI21X1_3845 ( .gnd(gnd), .vdd(vdd), .A(_13618__bF_buf3), .B(nonce_out_1_1_), .C(reset_bF_buf10), .Y(_13622_) );
AOI21X1 AOI21X1_2311 ( .gnd(gnd), .vdd(vdd), .A(_13621_), .B(_13620_), .C(_13622_), .Y(_13614__1_) );
NAND3X1 NAND3X1_813 ( .gnd(gnd), .vdd(vdd), .A(finished_3_bF_buf2), .B(nonce_out_3_2_), .C(_13615__bF_buf2), .Y(_13623_) );
AOI21X1 AOI21X1_2312 ( .gnd(gnd), .vdd(vdd), .A(finished_2_bF_buf1), .B(nonce_out_2_2_), .C(finished_1_bF_buf1), .Y(_13624_) );
OAI21X1 OAI21X1_3846 ( .gnd(gnd), .vdd(vdd), .A(_13618__bF_buf2), .B(nonce_out_1_2_), .C(reset_bF_buf9), .Y(_13625_) );
AOI21X1 AOI21X1_2313 ( .gnd(gnd), .vdd(vdd), .A(_13624_), .B(_13623_), .C(_13625_), .Y(_13614__2_) );
NAND3X1 NAND3X1_814 ( .gnd(gnd), .vdd(vdd), .A(finished_3_bF_buf1), .B(nonce_out_3_3_), .C(_13615__bF_buf1), .Y(_13626_) );
AOI21X1 AOI21X1_2314 ( .gnd(gnd), .vdd(vdd), .A(finished_2_bF_buf0), .B(nonce_out_2_3_), .C(finished_1_bF_buf0), .Y(_13627_) );
OAI21X1 OAI21X1_3847 ( .gnd(gnd), .vdd(vdd), .A(_13618__bF_buf1), .B(nonce_out_1_3_), .C(reset_bF_buf8), .Y(_13628_) );
AOI21X1 AOI21X1_2315 ( .gnd(gnd), .vdd(vdd), .A(_13627_), .B(_13626_), .C(_13628_), .Y(_13614__3_) );
NAND3X1 NAND3X1_815 ( .gnd(gnd), .vdd(vdd), .A(finished_3_bF_buf0), .B(nonce_out_3_4_), .C(_13615__bF_buf0), .Y(_13629_) );
AOI21X1 AOI21X1_2316 ( .gnd(gnd), .vdd(vdd), .A(finished_2_bF_buf4), .B(nonce_out_2_4_), .C(finished_1_bF_buf4), .Y(_13630_) );
OAI21X1 OAI21X1_3848 ( .gnd(gnd), .vdd(vdd), .A(_13618__bF_buf0), .B(nonce_out_1_4_), .C(reset_bF_buf7), .Y(_13631_) );
AOI21X1 AOI21X1_2317 ( .gnd(gnd), .vdd(vdd), .A(_13630_), .B(_13629_), .C(_13631_), .Y(_13614__4_) );
NAND3X1 NAND3X1_816 ( .gnd(gnd), .vdd(vdd), .A(finished_3_bF_buf4), .B(nonce_out_3_5_), .C(_13615__bF_buf4), .Y(_13632_) );
AOI21X1 AOI21X1_2318 ( .gnd(gnd), .vdd(vdd), .A(finished_2_bF_buf3), .B(nonce_out_2_5_), .C(finished_1_bF_buf3), .Y(_13633_) );
OAI21X1 OAI21X1_3849 ( .gnd(gnd), .vdd(vdd), .A(_13618__bF_buf4), .B(nonce_out_1_5_), .C(reset_bF_buf6), .Y(_13634_) );
AOI21X1 AOI21X1_2319 ( .gnd(gnd), .vdd(vdd), .A(_13633_), .B(_13632_), .C(_13634_), .Y(_13614__5_) );
NAND3X1 NAND3X1_817 ( .gnd(gnd), .vdd(vdd), .A(finished_3_bF_buf3), .B(nonce_out_3_6_), .C(_13615__bF_buf3), .Y(_13635_) );
AOI21X1 AOI21X1_2320 ( .gnd(gnd), .vdd(vdd), .A(finished_2_bF_buf2), .B(nonce_out_2_6_), .C(finished_1_bF_buf2), .Y(_13636_) );
OAI21X1 OAI21X1_3850 ( .gnd(gnd), .vdd(vdd), .A(_13618__bF_buf3), .B(nonce_out_1_6_), .C(reset_bF_buf5), .Y(_13637_) );
AOI21X1 AOI21X1_2321 ( .gnd(gnd), .vdd(vdd), .A(_13636_), .B(_13635_), .C(_13637_), .Y(_13614__6_) );
NAND3X1 NAND3X1_818 ( .gnd(gnd), .vdd(vdd), .A(finished_3_bF_buf2), .B(nonce_out_3_7_), .C(_13615__bF_buf2), .Y(_13638_) );
AOI21X1 AOI21X1_2322 ( .gnd(gnd), .vdd(vdd), .A(finished_2_bF_buf1), .B(nonce_out_2_7_), .C(finished_1_bF_buf1), .Y(_13639_) );
OAI21X1 OAI21X1_3851 ( .gnd(gnd), .vdd(vdd), .A(_13618__bF_buf2), .B(nonce_out_1_7_), .C(reset_bF_buf4), .Y(_13640_) );
AOI21X1 AOI21X1_2323 ( .gnd(gnd), .vdd(vdd), .A(_13639_), .B(_13638_), .C(_13640_), .Y(_13614__7_) );
NAND3X1 NAND3X1_819 ( .gnd(gnd), .vdd(vdd), .A(finished_3_bF_buf1), .B(nonce_out_3_8_), .C(_13615__bF_buf1), .Y(_13641_) );
AOI21X1 AOI21X1_2324 ( .gnd(gnd), .vdd(vdd), .A(finished_2_bF_buf0), .B(nonce_out_2_8_), .C(finished_1_bF_buf0), .Y(_13642_) );
OAI21X1 OAI21X1_3852 ( .gnd(gnd), .vdd(vdd), .A(_13618__bF_buf1), .B(nonce_out_1_8_), .C(reset_bF_buf3), .Y(_13643_) );
AOI21X1 AOI21X1_2325 ( .gnd(gnd), .vdd(vdd), .A(_13642_), .B(_13641_), .C(_13643_), .Y(_13614__8_) );
NAND3X1 NAND3X1_820 ( .gnd(gnd), .vdd(vdd), .A(finished_3_bF_buf0), .B(nonce_out_3_9_), .C(_13615__bF_buf0), .Y(_13644_) );
AOI21X1 AOI21X1_2326 ( .gnd(gnd), .vdd(vdd), .A(finished_2_bF_buf4), .B(nonce_out_2_9_), .C(finished_1_bF_buf4), .Y(_13645_) );
OAI21X1 OAI21X1_3853 ( .gnd(gnd), .vdd(vdd), .A(_13618__bF_buf0), .B(nonce_out_1_9_), .C(reset_bF_buf2), .Y(_13646_) );
AOI21X1 AOI21X1_2327 ( .gnd(gnd), .vdd(vdd), .A(_13645_), .B(_13644_), .C(_13646_), .Y(_13614__9_) );
NAND3X1 NAND3X1_821 ( .gnd(gnd), .vdd(vdd), .A(finished_3_bF_buf4), .B(nonce_out_3_10_), .C(_13615__bF_buf4), .Y(_13647_) );
AOI21X1 AOI21X1_2328 ( .gnd(gnd), .vdd(vdd), .A(finished_2_bF_buf3), .B(nonce_out_2_10_), .C(finished_1_bF_buf3), .Y(_13648_) );
OAI21X1 OAI21X1_3854 ( .gnd(gnd), .vdd(vdd), .A(_13618__bF_buf4), .B(nonce_out_1_10_), .C(reset_bF_buf1), .Y(_13649_) );
AOI21X1 AOI21X1_2329 ( .gnd(gnd), .vdd(vdd), .A(_13648_), .B(_13647_), .C(_13649_), .Y(_13614__10_) );
NAND3X1 NAND3X1_822 ( .gnd(gnd), .vdd(vdd), .A(finished_3_bF_buf3), .B(nonce_out_3_11_), .C(_13615__bF_buf3), .Y(_13650_) );
AOI21X1 AOI21X1_2330 ( .gnd(gnd), .vdd(vdd), .A(finished_2_bF_buf2), .B(nonce_out_2_11_), .C(finished_1_bF_buf2), .Y(_13651_) );
OAI21X1 OAI21X1_3855 ( .gnd(gnd), .vdd(vdd), .A(_13618__bF_buf3), .B(nonce_out_1_11_), .C(reset_bF_buf0), .Y(_13652_) );
AOI21X1 AOI21X1_2331 ( .gnd(gnd), .vdd(vdd), .A(_13651_), .B(_13650_), .C(_13652_), .Y(_13614__11_) );
NAND3X1 NAND3X1_823 ( .gnd(gnd), .vdd(vdd), .A(finished_3_bF_buf2), .B(nonce_out_3_12_), .C(_13615__bF_buf2), .Y(_13653_) );
AOI21X1 AOI21X1_2332 ( .gnd(gnd), .vdd(vdd), .A(finished_2_bF_buf1), .B(nonce_out_2_12_), .C(finished_1_bF_buf1), .Y(_13654_) );
OAI21X1 OAI21X1_3856 ( .gnd(gnd), .vdd(vdd), .A(_13618__bF_buf2), .B(nonce_out_1_12_), .C(reset_bF_buf10), .Y(_13655_) );
AOI21X1 AOI21X1_2333 ( .gnd(gnd), .vdd(vdd), .A(_13654_), .B(_13653_), .C(_13655_), .Y(_13614__12_) );
NAND3X1 NAND3X1_824 ( .gnd(gnd), .vdd(vdd), .A(finished_3_bF_buf1), .B(nonce_out_3_13_), .C(_13615__bF_buf1), .Y(_13656_) );
AOI21X1 AOI21X1_2334 ( .gnd(gnd), .vdd(vdd), .A(finished_2_bF_buf0), .B(nonce_out_2_13_), .C(finished_1_bF_buf0), .Y(_13657_) );
OAI21X1 OAI21X1_3857 ( .gnd(gnd), .vdd(vdd), .A(_13618__bF_buf1), .B(nonce_out_1_13_), .C(reset_bF_buf9), .Y(_13658_) );
AOI21X1 AOI21X1_2335 ( .gnd(gnd), .vdd(vdd), .A(_13657_), .B(_13656_), .C(_13658_), .Y(_13614__13_) );
NAND3X1 NAND3X1_825 ( .gnd(gnd), .vdd(vdd), .A(finished_3_bF_buf0), .B(nonce_out_3_14_), .C(_13615__bF_buf0), .Y(_13659_) );
AOI21X1 AOI21X1_2336 ( .gnd(gnd), .vdd(vdd), .A(finished_2_bF_buf4), .B(nonce_out_2_14_), .C(finished_1_bF_buf4), .Y(_13660_) );
OAI21X1 OAI21X1_3858 ( .gnd(gnd), .vdd(vdd), .A(_13618__bF_buf0), .B(nonce_out_1_14_), .C(reset_bF_buf8), .Y(_13661_) );
AOI21X1 AOI21X1_2337 ( .gnd(gnd), .vdd(vdd), .A(_13660_), .B(_13659_), .C(_13661_), .Y(_13614__14_) );
NAND3X1 NAND3X1_826 ( .gnd(gnd), .vdd(vdd), .A(finished_3_bF_buf4), .B(nonce_out_3_15_), .C(_13615__bF_buf4), .Y(_13662_) );
AOI21X1 AOI21X1_2338 ( .gnd(gnd), .vdd(vdd), .A(finished_2_bF_buf3), .B(nonce_out_2_15_), .C(finished_1_bF_buf3), .Y(_13663_) );
OAI21X1 OAI21X1_3859 ( .gnd(gnd), .vdd(vdd), .A(_13618__bF_buf4), .B(nonce_out_1_15_), .C(reset_bF_buf7), .Y(_13664_) );
AOI21X1 AOI21X1_2339 ( .gnd(gnd), .vdd(vdd), .A(_13663_), .B(_13662_), .C(_13664_), .Y(_13614__15_) );
NAND3X1 NAND3X1_827 ( .gnd(gnd), .vdd(vdd), .A(finished_3_bF_buf3), .B(nonce_out_3_16_), .C(_13615__bF_buf3), .Y(_13665_) );
AOI21X1 AOI21X1_2340 ( .gnd(gnd), .vdd(vdd), .A(finished_2_bF_buf2), .B(nonce_out_2_16_), .C(finished_1_bF_buf2), .Y(_13666_) );
OAI21X1 OAI21X1_3860 ( .gnd(gnd), .vdd(vdd), .A(_13618__bF_buf3), .B(nonce_out_1_16_), .C(reset_bF_buf6), .Y(_13667_) );
AOI21X1 AOI21X1_2341 ( .gnd(gnd), .vdd(vdd), .A(_13666_), .B(_13665_), .C(_13667_), .Y(_13614__16_) );
NAND3X1 NAND3X1_828 ( .gnd(gnd), .vdd(vdd), .A(finished_3_bF_buf2), .B(nonce_out_3_17_), .C(_13615__bF_buf2), .Y(_13668_) );
AOI21X1 AOI21X1_2342 ( .gnd(gnd), .vdd(vdd), .A(finished_2_bF_buf1), .B(nonce_out_2_17_), .C(finished_1_bF_buf1), .Y(_13669_) );
OAI21X1 OAI21X1_3861 ( .gnd(gnd), .vdd(vdd), .A(_13618__bF_buf2), .B(nonce_out_1_17_), .C(reset_bF_buf5), .Y(_13670_) );
AOI21X1 AOI21X1_2343 ( .gnd(gnd), .vdd(vdd), .A(_13669_), .B(_13668_), .C(_13670_), .Y(_13614__17_) );
NAND3X1 NAND3X1_829 ( .gnd(gnd), .vdd(vdd), .A(finished_3_bF_buf1), .B(nonce_out_3_18_), .C(_13615__bF_buf1), .Y(_13671_) );
AOI21X1 AOI21X1_2344 ( .gnd(gnd), .vdd(vdd), .A(finished_2_bF_buf0), .B(nonce_out_2_18_), .C(finished_1_bF_buf0), .Y(_13672_) );
OAI21X1 OAI21X1_3862 ( .gnd(gnd), .vdd(vdd), .A(_13618__bF_buf1), .B(nonce_out_1_18_), .C(reset_bF_buf4), .Y(_13673_) );
AOI21X1 AOI21X1_2345 ( .gnd(gnd), .vdd(vdd), .A(_13672_), .B(_13671_), .C(_13673_), .Y(_13614__18_) );
NAND3X1 NAND3X1_830 ( .gnd(gnd), .vdd(vdd), .A(finished_3_bF_buf0), .B(nonce_out_3_19_), .C(_13615__bF_buf0), .Y(_13674_) );
AOI21X1 AOI21X1_2346 ( .gnd(gnd), .vdd(vdd), .A(finished_2_bF_buf4), .B(nonce_out_2_19_), .C(finished_1_bF_buf4), .Y(_13675_) );
OAI21X1 OAI21X1_3863 ( .gnd(gnd), .vdd(vdd), .A(_13618__bF_buf0), .B(nonce_out_1_19_), .C(reset_bF_buf3), .Y(_13676_) );
AOI21X1 AOI21X1_2347 ( .gnd(gnd), .vdd(vdd), .A(_13675_), .B(_13674_), .C(_13676_), .Y(_13614__19_) );
NAND3X1 NAND3X1_831 ( .gnd(gnd), .vdd(vdd), .A(finished_3_bF_buf4), .B(nonce_out_3_20_), .C(_13615__bF_buf4), .Y(_13677_) );
AOI21X1 AOI21X1_2348 ( .gnd(gnd), .vdd(vdd), .A(finished_2_bF_buf3), .B(nonce_out_2_20_), .C(finished_1_bF_buf3), .Y(_13678_) );
OAI21X1 OAI21X1_3864 ( .gnd(gnd), .vdd(vdd), .A(_13618__bF_buf4), .B(nonce_out_1_20_), .C(reset_bF_buf2), .Y(_13679_) );
AOI21X1 AOI21X1_2349 ( .gnd(gnd), .vdd(vdd), .A(_13678_), .B(_13677_), .C(_13679_), .Y(_13614__20_) );
NAND3X1 NAND3X1_832 ( .gnd(gnd), .vdd(vdd), .A(finished_3_bF_buf3), .B(nonce_out_3_21_), .C(_13615__bF_buf3), .Y(_13680_) );
AOI21X1 AOI21X1_2350 ( .gnd(gnd), .vdd(vdd), .A(finished_2_bF_buf2), .B(nonce_out_2_21_), .C(finished_1_bF_buf2), .Y(_13681_) );
OAI21X1 OAI21X1_3865 ( .gnd(gnd), .vdd(vdd), .A(_13618__bF_buf3), .B(nonce_out_1_21_), .C(reset_bF_buf1), .Y(_13682_) );
AOI21X1 AOI21X1_2351 ( .gnd(gnd), .vdd(vdd), .A(_13681_), .B(_13680_), .C(_13682_), .Y(_13614__21_) );
NAND3X1 NAND3X1_833 ( .gnd(gnd), .vdd(vdd), .A(finished_3_bF_buf2), .B(nonce_out_3_22_), .C(_13615__bF_buf2), .Y(_13683_) );
AOI21X1 AOI21X1_2352 ( .gnd(gnd), .vdd(vdd), .A(finished_2_bF_buf1), .B(nonce_out_2_22_), .C(finished_1_bF_buf1), .Y(_13684_) );
OAI21X1 OAI21X1_3866 ( .gnd(gnd), .vdd(vdd), .A(_13618__bF_buf2), .B(nonce_out_1_22_), .C(reset_bF_buf0), .Y(_13685_) );
AOI21X1 AOI21X1_2353 ( .gnd(gnd), .vdd(vdd), .A(_13684_), .B(_13683_), .C(_13685_), .Y(_13614__22_) );
NAND3X1 NAND3X1_834 ( .gnd(gnd), .vdd(vdd), .A(finished_3_bF_buf1), .B(nonce_out_3_23_), .C(_13615__bF_buf1), .Y(_13686_) );
AOI21X1 AOI21X1_2354 ( .gnd(gnd), .vdd(vdd), .A(finished_2_bF_buf0), .B(nonce_out_2_23_), .C(finished_1_bF_buf0), .Y(_13687_) );
OAI21X1 OAI21X1_3867 ( .gnd(gnd), .vdd(vdd), .A(_13618__bF_buf1), .B(nonce_out_1_23_), .C(reset_bF_buf10), .Y(_13688_) );
AOI21X1 AOI21X1_2355 ( .gnd(gnd), .vdd(vdd), .A(_13687_), .B(_13686_), .C(_13688_), .Y(_13614__23_) );
NAND3X1 NAND3X1_835 ( .gnd(gnd), .vdd(vdd), .A(finished_3_bF_buf0), .B(nonce_out_3_24_), .C(_13615__bF_buf0), .Y(_13689_) );
AOI21X1 AOI21X1_2356 ( .gnd(gnd), .vdd(vdd), .A(finished_2_bF_buf4), .B(nonce_out_2_24_), .C(finished_1_bF_buf4), .Y(_13690_) );
OAI21X1 OAI21X1_3868 ( .gnd(gnd), .vdd(vdd), .A(_13618__bF_buf0), .B(nonce_out_1_24_), .C(reset_bF_buf9), .Y(_13691_) );
AOI21X1 AOI21X1_2357 ( .gnd(gnd), .vdd(vdd), .A(_13690_), .B(_13689_), .C(_13691_), .Y(_13614__24_) );
NAND3X1 NAND3X1_836 ( .gnd(gnd), .vdd(vdd), .A(finished_3_bF_buf4), .B(nonce_out_3_25_), .C(_13615__bF_buf4), .Y(_13692_) );
AOI21X1 AOI21X1_2358 ( .gnd(gnd), .vdd(vdd), .A(finished_2_bF_buf3), .B(nonce_out_2_25_), .C(finished_1_bF_buf3), .Y(_13693_) );
OAI21X1 OAI21X1_3869 ( .gnd(gnd), .vdd(vdd), .A(_13618__bF_buf4), .B(nonce_out_1_25_), .C(reset_bF_buf8), .Y(_13694_) );
AOI21X1 AOI21X1_2359 ( .gnd(gnd), .vdd(vdd), .A(_13693_), .B(_13692_), .C(_13694_), .Y(_13614__25_) );
NAND3X1 NAND3X1_837 ( .gnd(gnd), .vdd(vdd), .A(finished_3_bF_buf3), .B(nonce_out_3_26_), .C(_13615__bF_buf3), .Y(_13695_) );
AOI21X1 AOI21X1_2360 ( .gnd(gnd), .vdd(vdd), .A(finished_2_bF_buf2), .B(nonce_out_2_26_), .C(finished_1_bF_buf2), .Y(_13696_) );
OAI21X1 OAI21X1_3870 ( .gnd(gnd), .vdd(vdd), .A(_13618__bF_buf3), .B(nonce_out_1_26_), .C(reset_bF_buf7), .Y(_13697_) );
AOI21X1 AOI21X1_2361 ( .gnd(gnd), .vdd(vdd), .A(_13696_), .B(_13695_), .C(_13697_), .Y(_13614__26_) );
NAND3X1 NAND3X1_838 ( .gnd(gnd), .vdd(vdd), .A(finished_3_bF_buf2), .B(nonce_out_3_27_), .C(_13615__bF_buf2), .Y(_13698_) );
AOI21X1 AOI21X1_2362 ( .gnd(gnd), .vdd(vdd), .A(finished_2_bF_buf1), .B(nonce_out_2_27_), .C(finished_1_bF_buf1), .Y(_13699_) );
OAI21X1 OAI21X1_3871 ( .gnd(gnd), .vdd(vdd), .A(_13618__bF_buf2), .B(nonce_out_1_27_), .C(reset_bF_buf6), .Y(_13700_) );
AOI21X1 AOI21X1_2363 ( .gnd(gnd), .vdd(vdd), .A(_13699_), .B(_13698_), .C(_13700_), .Y(_13614__27_) );
NAND3X1 NAND3X1_839 ( .gnd(gnd), .vdd(vdd), .A(finished_3_bF_buf1), .B(nonce_out_3_28_), .C(_13615__bF_buf1), .Y(_13701_) );
AOI21X1 AOI21X1_2364 ( .gnd(gnd), .vdd(vdd), .A(finished_2_bF_buf0), .B(nonce_out_2_28_), .C(finished_1_bF_buf0), .Y(_13702_) );
OAI21X1 OAI21X1_3872 ( .gnd(gnd), .vdd(vdd), .A(_13618__bF_buf1), .B(nonce_out_1_28_), .C(reset_bF_buf5), .Y(_13703_) );
AOI21X1 AOI21X1_2365 ( .gnd(gnd), .vdd(vdd), .A(_13702_), .B(_13701_), .C(_13703_), .Y(_13614__28_) );
NAND3X1 NAND3X1_840 ( .gnd(gnd), .vdd(vdd), .A(finished_3_bF_buf0), .B(nonce_out_3_29_), .C(_13615__bF_buf0), .Y(_13704_) );
AOI21X1 AOI21X1_2366 ( .gnd(gnd), .vdd(vdd), .A(finished_2_bF_buf4), .B(nonce_out_2_29_), .C(finished_1_bF_buf4), .Y(_13705_) );
OAI21X1 OAI21X1_3873 ( .gnd(gnd), .vdd(vdd), .A(_13618__bF_buf0), .B(nonce_out_1_29_), .C(reset_bF_buf4), .Y(_13706_) );
AOI21X1 AOI21X1_2367 ( .gnd(gnd), .vdd(vdd), .A(_13705_), .B(_13704_), .C(_13706_), .Y(_13614__29_) );
NAND3X1 NAND3X1_841 ( .gnd(gnd), .vdd(vdd), .A(finished_3_bF_buf4), .B(nonce_out_3_30_), .C(_13615__bF_buf4), .Y(_13707_) );
AOI21X1 AOI21X1_2368 ( .gnd(gnd), .vdd(vdd), .A(finished_2_bF_buf3), .B(nonce_out_2_30_), .C(finished_1_bF_buf3), .Y(_13708_) );
OAI21X1 OAI21X1_3874 ( .gnd(gnd), .vdd(vdd), .A(_13618__bF_buf4), .B(nonce_out_1_30_), .C(reset_bF_buf3), .Y(_13709_) );
AOI21X1 AOI21X1_2369 ( .gnd(gnd), .vdd(vdd), .A(_13708_), .B(_13707_), .C(_13709_), .Y(_13614__30_) );
NAND3X1 NAND3X1_842 ( .gnd(gnd), .vdd(vdd), .A(finished_3_bF_buf3), .B(nonce_out_3_31_), .C(_13615__bF_buf3), .Y(_13710_) );
AOI21X1 AOI21X1_2370 ( .gnd(gnd), .vdd(vdd), .A(finished_2_bF_buf2), .B(nonce_out_2_31_), .C(finished_1_bF_buf2), .Y(_13711_) );
OAI21X1 OAI21X1_3875 ( .gnd(gnd), .vdd(vdd), .A(_13618__bF_buf3), .B(nonce_out_1_31_), .C(reset_bF_buf2), .Y(_13712_) );
AOI21X1 AOI21X1_2371 ( .gnd(gnd), .vdd(vdd), .A(_13711_), .B(_13710_), .C(_13712_), .Y(_13614__31_) );
NOR2X1 NOR2X1_2192 ( .gnd(gnd), .vdd(vdd), .A(finished_3_bF_buf2), .B(finished_2_bF_buf1), .Y(_13713_) );
NAND3X1 NAND3X1_843 ( .gnd(gnd), .vdd(vdd), .A(_13618__bF_buf2), .B(reset_bF_buf1), .C(_13713_), .Y(_13613_) );
DFFPOSX1 DFFPOSX1_1957 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_13613_), .Q(_0_) );
DFFPOSX1 DFFPOSX1_1958 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_13614__0_), .Q(_1__0_) );
DFFPOSX1 DFFPOSX1_1959 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_13614__1_), .Q(_1__1_) );
DFFPOSX1 DFFPOSX1_1960 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_13614__2_), .Q(_1__2_) );
DFFPOSX1 DFFPOSX1_1961 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_13614__3_), .Q(_1__3_) );
DFFPOSX1 DFFPOSX1_1962 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_13614__4_), .Q(_1__4_) );
DFFPOSX1 DFFPOSX1_1963 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_13614__5_), .Q(_1__5_) );
DFFPOSX1 DFFPOSX1_1964 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_13614__6_), .Q(_1__6_) );
DFFPOSX1 DFFPOSX1_1965 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_13614__7_), .Q(_1__7_) );
DFFPOSX1 DFFPOSX1_1966 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_13614__8_), .Q(_1__8_) );
DFFPOSX1 DFFPOSX1_1967 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_13614__9_), .Q(_1__9_) );
DFFPOSX1 DFFPOSX1_1968 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_13614__10_), .Q(_1__10_) );
DFFPOSX1 DFFPOSX1_1969 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_13614__11_), .Q(_1__11_) );
DFFPOSX1 DFFPOSX1_1970 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_13614__12_), .Q(_1__12_) );
DFFPOSX1 DFFPOSX1_1971 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_13614__13_), .Q(_1__13_) );
DFFPOSX1 DFFPOSX1_1972 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_13614__14_), .Q(_1__14_) );
DFFPOSX1 DFFPOSX1_1973 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_13614__15_), .Q(_1__15_) );
DFFPOSX1 DFFPOSX1_1974 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_13614__16_), .Q(_1__16_) );
DFFPOSX1 DFFPOSX1_1975 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_13614__17_), .Q(_1__17_) );
DFFPOSX1 DFFPOSX1_1976 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_13614__18_), .Q(_1__18_) );
DFFPOSX1 DFFPOSX1_1977 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_13614__19_), .Q(_1__19_) );
DFFPOSX1 DFFPOSX1_1978 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_13614__20_), .Q(_1__20_) );
DFFPOSX1 DFFPOSX1_1979 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_13614__21_), .Q(_1__21_) );
DFFPOSX1 DFFPOSX1_1980 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_13614__22_), .Q(_1__22_) );
DFFPOSX1 DFFPOSX1_1981 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_13614__23_), .Q(_1__23_) );
DFFPOSX1 DFFPOSX1_1982 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_13614__24_), .Q(_1__24_) );
DFFPOSX1 DFFPOSX1_1983 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_13614__25_), .Q(_1__25_) );
DFFPOSX1 DFFPOSX1_1984 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_13614__26_), .Q(_1__26_) );
DFFPOSX1 DFFPOSX1_1985 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_13614__27_), .Q(_1__27_) );
DFFPOSX1 DFFPOSX1_1986 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_13614__28_), .Q(_1__28_) );
DFFPOSX1 DFFPOSX1_1987 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_13614__29_), .Q(_1__29_) );
DFFPOSX1 DFFPOSX1_1988 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_13614__30_), .Q(_1__30_) );
DFFPOSX1 DFFPOSX1_1989 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_13614__31_), .Q(_1__31_) );
endmodule
